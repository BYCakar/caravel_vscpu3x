magic
tech sky130A
magscale 1 2
timestamp 1655402775
<< metal1 >>
rect 235166 700340 235172 700392
rect 235224 700380 235230 700392
rect 305638 700380 305644 700392
rect 235224 700352 305644 700380
rect 235224 700340 235230 700352
rect 305638 700340 305644 700352
rect 305696 700340 305702 700392
rect 57882 700272 57888 700324
rect 57940 700312 57946 700324
rect 543458 700312 543464 700324
rect 57940 700284 543464 700312
rect 57940 700272 57946 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 137830 683136 137836 683188
rect 137888 683176 137894 683188
rect 580166 683176 580172 683188
rect 137888 683148 580172 683176
rect 137888 683136 137894 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 299474 640976 299480 641028
rect 299532 641016 299538 641028
rect 400674 641016 400680 641028
rect 299532 640988 400680 641016
rect 299532 640976 299538 640988
rect 400674 640976 400680 640988
rect 400732 640976 400738 641028
rect 3418 639548 3424 639600
rect 3476 639588 3482 639600
rect 317046 639588 317052 639600
rect 3476 639560 317052 639588
rect 3476 639548 3482 639560
rect 317046 639548 317052 639560
rect 317104 639548 317110 639600
rect 104894 636828 104900 636880
rect 104952 636868 104958 636880
rect 429378 636868 429384 636880
rect 104952 636840 429384 636868
rect 104952 636828 104958 636840
rect 429378 636828 429384 636840
rect 429436 636828 429442 636880
rect 169754 635468 169760 635520
rect 169812 635508 169818 635520
rect 430942 635508 430948 635520
rect 169812 635480 430948 635508
rect 169812 635468 169818 635480
rect 430942 635468 430948 635480
rect 431000 635468 431006 635520
rect 316862 634856 316868 634908
rect 316920 634896 316926 634908
rect 430574 634896 430580 634908
rect 316920 634868 430580 634896
rect 316920 634856 316926 634868
rect 430574 634856 430580 634868
rect 430632 634856 430638 634908
rect 316954 634788 316960 634840
rect 317012 634828 317018 634840
rect 430850 634828 430856 634840
rect 317012 634800 430856 634828
rect 317012 634788 317018 634800
rect 430850 634788 430856 634800
rect 430908 634788 430914 634840
rect 318794 634040 318800 634092
rect 318852 634080 318858 634092
rect 494054 634080 494060 634092
rect 318852 634052 494060 634080
rect 318852 634040 318858 634052
rect 494054 634040 494060 634052
rect 494112 634040 494118 634092
rect 298094 633632 298100 633684
rect 298152 633672 298158 633684
rect 435358 633672 435364 633684
rect 298152 633644 435364 633672
rect 298152 633632 298158 633644
rect 435358 633632 435364 633644
rect 435416 633632 435422 633684
rect 289814 633564 289820 633616
rect 289872 633604 289878 633616
rect 432598 633604 432604 633616
rect 289872 633576 432604 633604
rect 289872 633564 289878 633576
rect 432598 633564 432604 633576
rect 432656 633564 432662 633616
rect 296714 633496 296720 633548
rect 296772 633536 296778 633548
rect 494330 633536 494336 633548
rect 296772 633508 494336 633536
rect 296772 633496 296778 633508
rect 494330 633496 494336 633508
rect 494388 633496 494394 633548
rect 288434 633428 288440 633480
rect 288492 633468 288498 633480
rect 510706 633468 510712 633480
rect 288492 633440 510712 633468
rect 288492 633428 288498 633440
rect 510706 633428 510712 633440
rect 510764 633428 510770 633480
rect 316678 632952 316684 633004
rect 316736 632992 316742 633004
rect 396626 632992 396632 633004
rect 316736 632964 396632 632992
rect 316736 632952 316742 632964
rect 396626 632952 396632 632964
rect 396684 632952 396690 633004
rect 300118 632884 300124 632936
rect 300176 632924 300182 632936
rect 378594 632924 378600 632936
rect 300176 632896 378600 632924
rect 300176 632884 300182 632896
rect 378594 632884 378600 632896
rect 378652 632884 378658 632936
rect 318242 632816 318248 632868
rect 318300 632856 318306 632868
rect 428182 632856 428188 632868
rect 318300 632828 428188 632856
rect 318300 632816 318306 632828
rect 428182 632816 428188 632828
rect 428240 632816 428246 632868
rect 312538 632748 312544 632800
rect 312596 632788 312602 632800
rect 337378 632788 337384 632800
rect 312596 632760 337384 632788
rect 312596 632748 312602 632760
rect 337378 632748 337384 632760
rect 337436 632748 337442 632800
rect 319438 632680 319444 632732
rect 319496 632720 319502 632732
rect 355410 632720 355416 632732
rect 319496 632692 355416 632720
rect 319496 632680 319502 632692
rect 355410 632680 355416 632692
rect 355468 632680 355474 632732
rect 364334 632680 364340 632732
rect 364392 632720 364398 632732
rect 423674 632720 423680 632732
rect 364392 632692 423680 632720
rect 364392 632680 364398 632692
rect 423674 632680 423680 632692
rect 423732 632680 423738 632732
rect 318150 632612 318156 632664
rect 318208 632652 318214 632664
rect 359918 632652 359924 632664
rect 318208 632624 359924 632652
rect 318208 632612 318214 632624
rect 359918 632612 359924 632624
rect 359976 632612 359982 632664
rect 307018 632544 307024 632596
rect 307076 632584 307082 632596
rect 350902 632584 350908 632596
rect 307076 632556 350908 632584
rect 307076 632544 307082 632556
rect 350902 632544 350908 632556
rect 350960 632544 350966 632596
rect 313918 632476 313924 632528
rect 313976 632516 313982 632528
rect 364426 632516 364432 632528
rect 313976 632488 364432 632516
rect 313976 632476 313982 632488
rect 364426 632476 364432 632488
rect 364484 632476 364490 632528
rect 319714 632408 319720 632460
rect 319772 632448 319778 632460
rect 373442 632448 373448 632460
rect 319772 632420 373448 632448
rect 319772 632408 319778 632420
rect 373442 632408 373448 632420
rect 373500 632408 373506 632460
rect 316770 632340 316776 632392
rect 316828 632380 316834 632392
rect 383102 632380 383108 632392
rect 316828 632352 383108 632380
rect 316828 632340 316834 632352
rect 383102 632340 383108 632352
rect 383160 632340 383166 632392
rect 314010 632272 314016 632324
rect 314068 632312 314074 632324
rect 387610 632312 387616 632324
rect 314068 632284 387616 632312
rect 314068 632272 314074 632284
rect 387610 632272 387616 632284
rect 387668 632272 387674 632324
rect 315298 632204 315304 632256
rect 315356 632244 315362 632256
rect 332870 632244 332876 632256
rect 315356 632216 332876 632244
rect 315356 632204 315362 632216
rect 332870 632204 332876 632216
rect 332928 632204 332934 632256
rect 320358 632136 320364 632188
rect 320416 632176 320422 632188
rect 341886 632176 341892 632188
rect 320416 632148 341892 632176
rect 320416 632136 320422 632148
rect 341886 632136 341892 632148
rect 341944 632136 341950 632188
rect 319622 632068 319628 632120
rect 319680 632108 319686 632120
rect 323854 632108 323860 632120
rect 319680 632080 323860 632108
rect 319680 632068 319686 632080
rect 323854 632068 323860 632080
rect 323912 632068 323918 632120
rect 414658 632068 414664 632120
rect 414716 632108 414722 632120
rect 457438 632108 457444 632120
rect 414716 632080 457444 632108
rect 414716 632068 414722 632080
rect 457438 632068 457444 632080
rect 457496 632068 457502 632120
rect 284938 631320 284944 631372
rect 284996 631360 285002 631372
rect 368934 631360 368940 631372
rect 284996 631332 368940 631360
rect 284996 631320 285002 631332
rect 368934 631320 368940 631332
rect 368992 631320 368998 631372
rect 285030 631252 285036 631304
rect 285088 631292 285094 631304
rect 419166 631292 419172 631304
rect 285088 631264 419172 631292
rect 285088 631252 285094 631264
rect 419166 631252 419172 631264
rect 419224 631252 419230 631304
rect 298186 631184 298192 631236
rect 298244 631224 298250 631236
rect 432690 631224 432696 631236
rect 298244 631196 432696 631224
rect 298244 631184 298250 631196
rect 432690 631184 432696 631196
rect 432748 631184 432754 631236
rect 319806 631116 319812 631168
rect 319864 631156 319870 631168
rect 457530 631156 457536 631168
rect 319864 631128 457536 631156
rect 319864 631116 319870 631128
rect 457530 631116 457536 631128
rect 457588 631116 457594 631168
rect 291194 631048 291200 631100
rect 291252 631088 291258 631100
rect 429838 631088 429844 631100
rect 291252 631060 429844 631088
rect 291252 631048 291258 631060
rect 429838 631048 429844 631060
rect 429896 631048 429902 631100
rect 318058 630980 318064 631032
rect 318116 631020 318122 631032
rect 471146 631020 471152 631032
rect 318116 630992 471152 631020
rect 318116 630980 318122 630992
rect 471146 630980 471152 630992
rect 471204 630980 471210 631032
rect 293954 630912 293960 630964
rect 294012 630952 294018 630964
rect 510614 630952 510620 630964
rect 294012 630924 510620 630952
rect 294012 630912 294018 630924
rect 510614 630912 510620 630924
rect 510672 630912 510678 630964
rect 287054 630844 287060 630896
rect 287112 630884 287118 630896
rect 511994 630884 512000 630896
rect 287112 630856 512000 630884
rect 287112 630844 287118 630856
rect 511994 630844 512000 630856
rect 512052 630844 512058 630896
rect 319070 630776 319076 630828
rect 319128 630816 319134 630828
rect 580166 630816 580172 630828
rect 319128 630788 580172 630816
rect 319128 630776 319134 630788
rect 580166 630776 580172 630788
rect 580224 630776 580230 630828
rect 18598 630708 18604 630760
rect 18656 630748 18662 630760
rect 409874 630748 409880 630760
rect 18656 630720 409880 630748
rect 18656 630708 18662 630720
rect 409874 630708 409880 630720
rect 409932 630708 409938 630760
rect 218698 630640 218704 630692
rect 218756 630680 218762 630692
rect 414566 630680 414572 630692
rect 218756 630652 414572 630680
rect 218756 630640 218762 630652
rect 414566 630640 414572 630652
rect 414624 630640 414630 630692
rect 320358 630476 320364 630488
rect 316006 630448 320364 630476
rect 280706 629960 280712 630012
rect 280764 630000 280770 630012
rect 316006 630000 316034 630448
rect 320358 630436 320364 630448
rect 320416 630436 320422 630488
rect 280764 629972 316034 630000
rect 280764 629960 280770 629972
rect 217778 629892 217784 629944
rect 217836 629932 217842 629944
rect 319070 629932 319076 629944
rect 217836 629904 319076 629932
rect 217836 629892 217842 629904
rect 319070 629892 319076 629904
rect 319128 629892 319134 629944
rect 309778 629280 309784 629332
rect 309836 629320 309842 629332
rect 317782 629320 317788 629332
rect 309836 629292 317788 629320
rect 309836 629280 309842 629292
rect 317782 629280 317788 629292
rect 317840 629280 317846 629332
rect 100570 625744 100576 625796
rect 100628 625784 100634 625796
rect 124674 625784 124680 625796
rect 100628 625756 124680 625784
rect 100628 625744 100634 625756
rect 124674 625744 124680 625756
rect 124732 625744 124738 625796
rect 213914 625744 213920 625796
rect 213972 625784 213978 625796
rect 225414 625784 225420 625796
rect 213972 625756 225420 625784
rect 213972 625744 213978 625756
rect 225414 625744 225420 625756
rect 225472 625744 225478 625796
rect 115382 625676 115388 625728
rect 115440 625716 115446 625728
rect 124582 625716 124588 625728
rect 115440 625688 124588 625716
rect 115440 625676 115446 625688
rect 124582 625676 124588 625688
rect 124640 625676 124646 625728
rect 137738 625676 137744 625728
rect 137796 625716 137802 625728
rect 186498 625716 186504 625728
rect 137796 625688 186504 625716
rect 137796 625676 137802 625688
rect 186498 625676 186504 625688
rect 186556 625676 186562 625728
rect 206462 625676 206468 625728
rect 206520 625716 206526 625728
rect 231302 625716 231308 625728
rect 206520 625688 231308 625716
rect 206520 625676 206526 625688
rect 231302 625676 231308 625688
rect 231360 625676 231366 625728
rect 112162 625608 112168 625660
rect 112220 625648 112226 625660
rect 124490 625648 124496 625660
rect 112220 625620 124496 625648
rect 112220 625608 112226 625620
rect 124490 625608 124496 625620
rect 124548 625608 124554 625660
rect 139302 625608 139308 625660
rect 139360 625648 139366 625660
rect 162854 625648 162860 625660
rect 139360 625620 162860 625648
rect 139360 625608 139366 625620
rect 162854 625608 162860 625620
rect 162912 625608 162918 625660
rect 212534 625608 212540 625660
rect 212592 625648 212598 625660
rect 271874 625648 271880 625660
rect 212592 625620 271880 625648
rect 212592 625608 212598 625620
rect 271874 625608 271880 625620
rect 271932 625608 271938 625660
rect 83182 625540 83188 625592
rect 83240 625580 83246 625592
rect 125686 625580 125692 625592
rect 83240 625552 125692 625580
rect 83240 625540 83246 625552
rect 125686 625540 125692 625552
rect 125744 625540 125750 625592
rect 135162 625540 135168 625592
rect 135220 625580 135226 625592
rect 160278 625580 160284 625592
rect 135220 625552 160284 625580
rect 135220 625540 135226 625552
rect 160278 625540 160284 625552
rect 160336 625540 160342 625592
rect 217870 625540 217876 625592
rect 217928 625580 217934 625592
rect 242894 625580 242900 625592
rect 217928 625552 242900 625580
rect 217928 625540 217934 625552
rect 242894 625540 242900 625552
rect 242952 625540 242958 625592
rect 109586 625472 109592 625524
rect 109644 625512 109650 625524
rect 122834 625512 122840 625524
rect 109644 625484 122840 625512
rect 109644 625472 109650 625484
rect 122834 625472 122840 625484
rect 122892 625472 122898 625524
rect 136358 625472 136364 625524
rect 136416 625512 136422 625524
rect 166166 625512 166172 625524
rect 136416 625484 166172 625512
rect 136416 625472 136422 625484
rect 166166 625472 166172 625484
rect 166224 625472 166230 625524
rect 218882 625472 218888 625524
rect 218940 625512 218946 625524
rect 251910 625512 251916 625524
rect 218940 625484 251916 625512
rect 218940 625472 218946 625484
rect 251910 625472 251916 625484
rect 251968 625472 251974 625524
rect 106366 625404 106372 625456
rect 106424 625444 106430 625456
rect 120902 625444 120908 625456
rect 106424 625416 120908 625444
rect 106424 625404 106430 625416
rect 120902 625404 120908 625416
rect 120960 625404 120966 625456
rect 139118 625404 139124 625456
rect 139176 625444 139182 625456
rect 174446 625444 174452 625456
rect 139176 625416 174452 625444
rect 139176 625404 139182 625416
rect 174446 625404 174452 625416
rect 174504 625404 174510 625456
rect 218790 625404 218796 625456
rect 218848 625444 218854 625456
rect 263594 625444 263600 625456
rect 218848 625416 263600 625444
rect 218848 625404 218854 625416
rect 263594 625404 263600 625416
rect 263652 625404 263658 625456
rect 103790 625336 103796 625388
rect 103848 625376 103854 625388
rect 122282 625376 122288 625388
rect 103848 625348 122288 625376
rect 103848 625336 103854 625348
rect 122282 625336 122288 625348
rect 122340 625336 122346 625388
rect 134886 625336 134892 625388
rect 134944 625376 134950 625388
rect 180334 625376 180340 625388
rect 134944 625348 180340 625376
rect 134944 625336 134950 625348
rect 180334 625336 180340 625348
rect 180392 625336 180398 625388
rect 189994 625336 190000 625388
rect 190052 625376 190058 625388
rect 204438 625376 204444 625388
rect 190052 625348 204444 625376
rect 190052 625336 190058 625348
rect 204438 625336 204444 625348
rect 204496 625336 204502 625388
rect 209774 625336 209780 625388
rect 209832 625376 209838 625388
rect 260190 625376 260196 625388
rect 209832 625348 260196 625376
rect 209832 625336 209838 625348
rect 260190 625336 260196 625348
rect 260248 625336 260254 625388
rect 54846 625268 54852 625320
rect 54904 625308 54910 625320
rect 88978 625308 88984 625320
rect 54904 625280 88984 625308
rect 54904 625268 54910 625280
rect 88978 625268 88984 625280
rect 89036 625268 89042 625320
rect 124214 625268 124220 625320
rect 124272 625308 124278 625320
rect 171870 625308 171876 625320
rect 124272 625280 171876 625308
rect 124272 625268 124278 625280
rect 171870 625268 171876 625280
rect 171928 625268 171934 625320
rect 214006 625268 214012 625320
rect 214064 625308 214070 625320
rect 269206 625308 269212 625320
rect 214064 625280 269212 625308
rect 214064 625268 214070 625280
rect 269206 625268 269212 625280
rect 269264 625268 269270 625320
rect 55122 625200 55128 625252
rect 55180 625240 55186 625252
rect 92198 625240 92204 625252
rect 55180 625212 92204 625240
rect 55180 625200 55186 625212
rect 92198 625200 92204 625212
rect 92256 625200 92262 625252
rect 94774 625200 94780 625252
rect 94832 625240 94838 625252
rect 121638 625240 121644 625252
rect 94832 625212 121644 625240
rect 94832 625200 94838 625212
rect 121638 625200 121644 625212
rect 121696 625200 121702 625252
rect 135254 625200 135260 625252
rect 135312 625240 135318 625252
rect 183646 625240 183652 625252
rect 135312 625212 183652 625240
rect 135312 625200 135318 625212
rect 183646 625200 183652 625212
rect 183704 625200 183710 625252
rect 192570 625200 192576 625252
rect 192628 625240 192634 625252
rect 201678 625240 201684 625252
rect 192628 625212 201684 625240
rect 192628 625200 192634 625212
rect 201678 625200 201684 625212
rect 201736 625200 201742 625252
rect 219342 625200 219348 625252
rect 219400 625240 219406 625252
rect 275094 625240 275100 625252
rect 219400 625212 275100 625240
rect 219400 625200 219406 625212
rect 275094 625200 275100 625212
rect 275152 625200 275158 625252
rect 56502 625132 56508 625184
rect 56560 625172 56566 625184
rect 77386 625172 77392 625184
rect 56560 625144 77392 625172
rect 56560 625132 56566 625144
rect 77386 625132 77392 625144
rect 77444 625132 77450 625184
rect 133874 625132 133880 625184
rect 133932 625172 133938 625184
rect 133932 625144 139808 625172
rect 133932 625132 133938 625144
rect 139780 625104 139808 625144
rect 139854 625132 139860 625184
rect 139912 625172 139918 625184
rect 157518 625172 157524 625184
rect 139912 625144 157524 625172
rect 139912 625132 139918 625144
rect 157518 625132 157524 625144
rect 157576 625132 157582 625184
rect 195698 625132 195704 625184
rect 195756 625172 195762 625184
rect 200850 625172 200856 625184
rect 195756 625144 200856 625172
rect 195756 625132 195762 625144
rect 200850 625132 200856 625144
rect 200908 625132 200914 625184
rect 289078 625132 289084 625184
rect 289136 625172 289142 625184
rect 317598 625172 317604 625184
rect 289136 625144 317604 625172
rect 289136 625132 289142 625144
rect 317598 625132 317604 625144
rect 317656 625132 317662 625184
rect 140130 625104 140136 625116
rect 139780 625076 140136 625104
rect 140130 625064 140136 625076
rect 140188 625064 140194 625116
rect 215294 624044 215300 624096
rect 215352 624084 215358 624096
rect 234614 624084 234620 624096
rect 215352 624056 234620 624084
rect 215352 624044 215358 624056
rect 234614 624044 234620 624056
rect 234672 624044 234678 624096
rect 219618 623976 219624 624028
rect 219676 624016 219682 624028
rect 246022 624016 246028 624028
rect 219676 623988 246028 624016
rect 219676 623976 219682 623988
rect 246022 623976 246028 623988
rect 246080 623976 246086 624028
rect 59354 623908 59360 623960
rect 59412 623948 59418 623960
rect 97994 623948 98000 623960
rect 59412 623920 98000 623948
rect 59412 623908 59418 623920
rect 97994 623908 98000 623920
rect 98052 623908 98058 623960
rect 210418 623908 210424 623960
rect 210476 623948 210482 623960
rect 237558 623948 237564 623960
rect 210476 623920 237564 623948
rect 210476 623908 210482 623920
rect 237558 623908 237564 623920
rect 237616 623908 237622 623960
rect 57790 623840 57796 623892
rect 57848 623880 57854 623892
rect 80606 623880 80612 623892
rect 57848 623852 80612 623880
rect 57848 623840 57854 623852
rect 80606 623840 80612 623852
rect 80664 623840 80670 623892
rect 86402 623840 86408 623892
rect 86460 623880 86466 623892
rect 124306 623880 124312 623892
rect 86460 623852 124312 623880
rect 86460 623840 86466 623852
rect 124306 623840 124312 623852
rect 124364 623840 124370 623892
rect 133138 623840 133144 623892
rect 133196 623880 133202 623892
rect 151262 623880 151268 623892
rect 133196 623852 151268 623880
rect 133196 623840 133202 623852
rect 151262 623840 151268 623852
rect 151320 623840 151326 623892
rect 206278 623840 206284 623892
rect 206336 623880 206342 623892
rect 254486 623880 254492 623892
rect 206336 623852 254492 623880
rect 206336 623840 206342 623852
rect 254486 623840 254492 623852
rect 254544 623840 254550 623892
rect 69014 623772 69020 623824
rect 69072 623812 69078 623824
rect 124398 623812 124404 623824
rect 69072 623784 124404 623812
rect 69072 623772 69078 623784
rect 124398 623772 124404 623784
rect 124456 623772 124462 623824
rect 136634 623772 136640 623824
rect 136692 623812 136698 623824
rect 168742 623812 168748 623824
rect 136692 623784 168748 623812
rect 136692 623772 136698 623784
rect 168742 623772 168748 623784
rect 168800 623772 168806 623824
rect 204254 623772 204260 623824
rect 204312 623812 204318 623824
rect 277670 623812 277676 623824
rect 204312 623784 277676 623812
rect 204312 623772 204318 623784
rect 277670 623772 277676 623784
rect 277728 623772 277734 623824
rect 217962 622820 217968 622872
rect 218020 622860 218026 622872
rect 228726 622860 228732 622872
rect 218020 622832 228732 622860
rect 218020 622820 218026 622832
rect 228726 622820 228732 622832
rect 228784 622820 228790 622872
rect 135070 622752 135076 622804
rect 135128 622792 135134 622804
rect 145558 622792 145564 622804
rect 135128 622764 145564 622792
rect 135128 622752 135134 622764
rect 145558 622752 145564 622764
rect 145616 622752 145622 622804
rect 214558 622752 214564 622804
rect 214616 622792 214622 622804
rect 257614 622792 257620 622804
rect 214616 622764 257620 622792
rect 214616 622752 214622 622764
rect 257614 622752 257620 622764
rect 257672 622752 257678 622804
rect 126238 622684 126244 622736
rect 126296 622724 126302 622736
rect 177850 622724 177856 622736
rect 126296 622696 177856 622724
rect 126296 622684 126302 622696
rect 177850 622684 177856 622696
rect 177908 622684 177914 622736
rect 204346 622684 204352 622736
rect 204404 622724 204410 622736
rect 222838 622724 222844 622736
rect 204404 622696 222844 622724
rect 204404 622684 204410 622696
rect 222838 622684 222844 622696
rect 222896 622684 222902 622736
rect 55030 622616 55036 622668
rect 55088 622656 55094 622668
rect 62942 622656 62948 622668
rect 55088 622628 62948 622656
rect 55088 622616 55094 622628
rect 62942 622616 62948 622628
rect 63000 622616 63006 622668
rect 136450 622616 136456 622668
rect 136508 622656 136514 622668
rect 149146 622656 149152 622668
rect 136508 622628 149152 622656
rect 136508 622616 136514 622628
rect 149146 622616 149152 622628
rect 149204 622616 149210 622668
rect 208394 622616 208400 622668
rect 208452 622656 208458 622668
rect 240318 622656 240324 622668
rect 208452 622628 240324 622656
rect 208452 622616 208458 622628
rect 240318 622616 240324 622628
rect 240376 622616 240382 622668
rect 54938 622548 54944 622600
rect 54996 622588 55002 622600
rect 65518 622588 65524 622600
rect 54996 622560 65524 622588
rect 54996 622548 55002 622560
rect 65518 622548 65524 622560
rect 65576 622548 65582 622600
rect 136542 622548 136548 622600
rect 136600 622588 136606 622600
rect 154574 622588 154580 622600
rect 136600 622560 154580 622588
rect 136600 622548 136606 622560
rect 154574 622548 154580 622560
rect 154632 622548 154638 622600
rect 206370 622548 206376 622600
rect 206428 622588 206434 622600
rect 248690 622588 248696 622600
rect 206428 622560 248696 622588
rect 206428 622548 206434 622560
rect 248690 622548 248696 622560
rect 248748 622548 248754 622600
rect 56318 622480 56324 622532
rect 56376 622520 56382 622532
rect 71222 622520 71228 622532
rect 56376 622492 71228 622520
rect 56376 622480 56382 622492
rect 71222 622480 71228 622492
rect 71280 622480 71286 622532
rect 134978 622480 134984 622532
rect 135036 622520 135042 622532
rect 142982 622520 142988 622532
rect 135036 622492 142988 622520
rect 135036 622480 135042 622492
rect 142982 622480 142988 622492
rect 143040 622480 143046 622532
rect 211798 622480 211804 622532
rect 211856 622520 211862 622532
rect 266262 622520 266268 622532
rect 211856 622492 266268 622520
rect 211856 622480 211862 622492
rect 266262 622480 266268 622492
rect 266320 622480 266326 622532
rect 280706 622480 280712 622532
rect 280764 622480 280770 622532
rect 56410 622412 56416 622464
rect 56468 622452 56474 622464
rect 74626 622452 74632 622464
rect 56468 622424 74632 622452
rect 56468 622412 56474 622424
rect 74626 622412 74632 622424
rect 74684 622412 74690 622464
rect 137922 622412 137928 622464
rect 137980 622452 137986 622464
rect 218698 622452 218704 622464
rect 137980 622424 218704 622452
rect 137980 622412 137986 622424
rect 218698 622412 218704 622424
rect 218756 622412 218762 622464
rect 118234 622344 118240 622396
rect 118292 622384 118298 622396
rect 121546 622384 121552 622396
rect 118292 622356 121552 622384
rect 118292 622344 118298 622356
rect 121546 622344 121552 622356
rect 121604 622344 121610 622396
rect 198274 622344 198280 622396
rect 198332 622384 198338 622396
rect 202230 622384 202236 622396
rect 198332 622356 202236 622384
rect 198332 622344 198338 622356
rect 202230 622344 202236 622356
rect 202288 622344 202294 622396
rect 217318 622344 217324 622396
rect 217376 622384 217382 622396
rect 219710 622384 219716 622396
rect 217376 622356 219716 622384
rect 217376 622344 217382 622356
rect 219710 622344 219716 622356
rect 219768 622344 219774 622396
rect 280724 622328 280752 622480
rect 280706 622276 280712 622328
rect 280764 622276 280770 622328
rect 432598 621732 432604 621784
rect 432656 621772 432662 621784
rect 483198 621772 483204 621784
rect 432656 621744 483204 621772
rect 432656 621732 432662 621744
rect 483198 621732 483204 621744
rect 483256 621732 483262 621784
rect 432690 621664 432696 621716
rect 432748 621704 432754 621716
rect 501230 621704 501236 621716
rect 432748 621676 501236 621704
rect 432748 621664 432754 621676
rect 501230 621664 501236 621676
rect 501288 621664 501294 621716
rect 465166 620984 465172 621036
rect 465224 621024 465230 621036
rect 515398 621024 515404 621036
rect 465224 620996 515404 621024
rect 465224 620984 465230 620996
rect 515398 620984 515404 620996
rect 515456 620984 515462 621036
rect 429838 620916 429844 620968
rect 429896 620956 429902 620968
rect 456794 620956 456800 620968
rect 429896 620928 456800 620956
rect 429896 620916 429902 620928
rect 456794 620916 456800 620928
rect 456852 620916 456858 620968
rect 213178 619624 213184 619676
rect 213236 619664 213242 619676
rect 216674 619664 216680 619676
rect 213236 619636 216680 619664
rect 213236 619624 213242 619636
rect 216674 619624 216680 619636
rect 216732 619624 216738 619676
rect 311158 619624 311164 619676
rect 311216 619664 311222 619676
rect 317966 619664 317972 619676
rect 311216 619636 317972 619664
rect 311216 619624 311222 619636
rect 317966 619624 317972 619636
rect 318024 619624 318030 619676
rect 208486 616836 208492 616888
rect 208544 616876 208550 616888
rect 216674 616876 216680 616888
rect 208544 616848 216680 616876
rect 208544 616836 208550 616848
rect 216674 616836 216680 616848
rect 216732 616836 216738 616888
rect 286318 615476 286324 615528
rect 286376 615516 286382 615528
rect 317966 615516 317972 615528
rect 286376 615488 317972 615516
rect 286376 615476 286382 615488
rect 317966 615476 317972 615488
rect 318024 615476 318030 615528
rect 287698 609968 287704 610020
rect 287756 610008 287762 610020
rect 317874 610008 317880 610020
rect 287756 609980 317880 610008
rect 287756 609968 287762 609980
rect 317874 609968 317880 609980
rect 317932 609968 317938 610020
rect 435358 608540 435364 608592
rect 435416 608580 435422 608592
rect 456794 608580 456800 608592
rect 435416 608552 456800 608580
rect 435416 608540 435422 608552
rect 456794 608540 456800 608552
rect 456852 608540 456858 608592
rect 132494 607180 132500 607232
rect 132552 607220 132558 607232
rect 136726 607220 136732 607232
rect 132552 607192 136732 607220
rect 132552 607180 132558 607192
rect 136726 607180 136732 607192
rect 136784 607180 136790 607232
rect 204898 607180 204904 607232
rect 204956 607220 204962 607232
rect 216674 607220 216680 607232
rect 204956 607192 216680 607220
rect 204956 607180 204962 607192
rect 216674 607180 216680 607192
rect 216732 607180 216738 607232
rect 304258 605820 304264 605872
rect 304316 605860 304322 605872
rect 317966 605860 317972 605872
rect 304316 605832 317972 605860
rect 304316 605820 304322 605832
rect 317966 605820 317972 605832
rect 318024 605820 318030 605872
rect 294598 600312 294604 600364
rect 294656 600352 294662 600364
rect 317598 600352 317604 600364
rect 294656 600324 317604 600352
rect 294656 600312 294662 600324
rect 317598 600312 317604 600324
rect 317656 600312 317662 600364
rect 200942 598000 200948 598052
rect 201000 598040 201006 598052
rect 203058 598040 203064 598052
rect 201000 598012 203064 598040
rect 201000 598000 201006 598012
rect 203058 598000 203064 598012
rect 203116 598000 203122 598052
rect 287790 596164 287796 596216
rect 287848 596204 287854 596216
rect 317598 596204 317604 596216
rect 287848 596176 317604 596204
rect 287848 596164 287854 596176
rect 317598 596164 317604 596176
rect 317656 596164 317662 596216
rect 207014 593376 207020 593428
rect 207072 593416 207078 593428
rect 216674 593416 216680 593428
rect 207072 593388 216680 593416
rect 207072 593376 207078 593388
rect 216674 593376 216680 593388
rect 216732 593376 216738 593428
rect 302234 589908 302240 589960
rect 302292 589948 302298 589960
rect 319806 589948 319812 589960
rect 302292 589920 319812 589948
rect 302292 589908 302298 589920
rect 319806 589908 319812 589920
rect 319864 589908 319870 589960
rect 124122 589364 124128 589416
rect 124180 589404 124186 589416
rect 134610 589404 134616 589416
rect 124180 589376 134616 589404
rect 124180 589364 124186 589376
rect 134610 589364 134616 589376
rect 134668 589364 134674 589416
rect 134518 589296 134524 589348
rect 134576 589336 134582 589348
rect 136726 589336 136732 589348
rect 134576 589308 136732 589336
rect 134576 589296 134582 589308
rect 136726 589296 136732 589308
rect 136784 589296 136790 589348
rect 203242 589296 203248 589348
rect 203300 589336 203306 589348
rect 204530 589336 204536 589348
rect 203300 589308 204536 589336
rect 203300 589296 203306 589308
rect 204530 589296 204536 589308
rect 204588 589296 204594 589348
rect 210510 589296 210516 589348
rect 210568 589336 210574 589348
rect 216674 589336 216680 589348
rect 210568 589308 216680 589336
rect 210568 589296 210574 589308
rect 216674 589296 216680 589308
rect 216732 589296 216738 589348
rect 283650 589296 283656 589348
rect 283708 589336 283714 589348
rect 302234 589336 302240 589348
rect 283708 589308 302240 589336
rect 283708 589296 283714 589308
rect 302234 589296 302240 589308
rect 302292 589296 302298 589348
rect 211154 586848 211160 586900
rect 211212 586888 211218 586900
rect 216674 586888 216680 586900
rect 211212 586860 216680 586888
rect 211212 586848 211218 586860
rect 216674 586848 216680 586860
rect 216732 586848 216738 586900
rect 293218 586508 293224 586560
rect 293276 586548 293282 586560
rect 317414 586548 317420 586560
rect 293276 586520 317420 586548
rect 293276 586508 293282 586520
rect 317414 586508 317420 586520
rect 317472 586508 317478 586560
rect 515398 585760 515404 585812
rect 515456 585800 515462 585812
rect 580166 585800 580172 585812
rect 515456 585772 580172 585800
rect 515456 585760 515462 585772
rect 580166 585760 580172 585772
rect 580224 585760 580230 585812
rect 57514 583720 57520 583772
rect 57572 583760 57578 583772
rect 58618 583760 58624 583772
rect 57572 583732 58624 583760
rect 57572 583720 57578 583732
rect 58618 583720 58624 583732
rect 58676 583720 58682 583772
rect 304350 582360 304356 582412
rect 304408 582400 304414 582412
rect 317966 582400 317972 582412
rect 304408 582372 317972 582400
rect 304408 582360 304414 582372
rect 317966 582360 317972 582372
rect 318024 582360 318030 582412
rect 217686 581680 217692 581732
rect 217744 581720 217750 581732
rect 218698 581720 218704 581732
rect 217744 581692 218704 581720
rect 217744 581680 217750 581692
rect 218698 581680 218704 581692
rect 218756 581680 218762 581732
rect 125594 576852 125600 576904
rect 125652 576892 125658 576904
rect 136726 576892 136732 576904
rect 125652 576864 136732 576892
rect 125652 576852 125658 576864
rect 136726 576852 136732 576864
rect 136784 576852 136790 576904
rect 300210 576852 300216 576904
rect 300268 576892 300274 576904
rect 317874 576892 317880 576904
rect 300268 576864 317880 576892
rect 300268 576852 300274 576864
rect 317874 576852 317880 576864
rect 317932 576852 317938 576904
rect 206554 574064 206560 574116
rect 206612 574104 206618 574116
rect 216674 574104 216680 574116
rect 206612 574076 216680 574104
rect 206612 574064 206618 574076
rect 216674 574064 216680 574076
rect 216732 574064 216738 574116
rect 513282 572704 513288 572756
rect 513340 572744 513346 572756
rect 560938 572744 560944 572756
rect 513340 572716 560944 572744
rect 513340 572704 513346 572716
rect 560938 572704 560944 572716
rect 560996 572704 561002 572756
rect 57330 572296 57336 572348
rect 57388 572336 57394 572348
rect 58710 572336 58716 572348
rect 57388 572308 58716 572336
rect 57388 572296 57394 572308
rect 58710 572296 58716 572308
rect 58768 572296 58774 572348
rect 210602 571344 210608 571396
rect 210660 571384 210666 571396
rect 216674 571384 216680 571396
rect 210660 571356 216680 571384
rect 210660 571344 210666 571356
rect 216674 571344 216680 571356
rect 216732 571344 216738 571396
rect 289170 571344 289176 571396
rect 289228 571384 289234 571396
rect 317966 571384 317972 571396
rect 289228 571356 317972 571384
rect 289228 571344 289234 571356
rect 317966 571344 317972 571356
rect 318024 571344 318030 571396
rect 209038 562300 209044 562352
rect 209096 562340 209102 562352
rect 217410 562340 217416 562352
rect 209096 562312 217416 562340
rect 209096 562300 209102 562312
rect 217410 562300 217416 562312
rect 217468 562300 217474 562352
rect 57882 561144 57888 561196
rect 57940 561184 57946 561196
rect 137278 561184 137284 561196
rect 57940 561156 137284 561184
rect 57940 561144 57946 561156
rect 137278 561144 137284 561156
rect 137336 561144 137342 561196
rect 3418 561076 3424 561128
rect 3476 561116 3482 561128
rect 304350 561116 304356 561128
rect 3476 561088 304356 561116
rect 3476 561076 3482 561088
rect 304350 561076 304356 561088
rect 304408 561076 304414 561128
rect 201034 560464 201040 560516
rect 201092 560504 201098 560516
rect 202874 560504 202880 560516
rect 201092 560476 202880 560504
rect 201092 560464 201098 560476
rect 202874 560464 202880 560476
rect 202932 560464 202938 560516
rect 217686 560260 217692 560312
rect 217744 560300 217750 560312
rect 220170 560300 220176 560312
rect 217744 560272 220176 560300
rect 217744 560260 217750 560272
rect 220170 560260 220176 560272
rect 220228 560260 220234 560312
rect 57146 560192 57152 560244
rect 57204 560232 57210 560244
rect 62114 560232 62120 560244
rect 57204 560204 62120 560232
rect 57204 560192 57210 560204
rect 62114 560192 62120 560204
rect 62172 560192 62178 560244
rect 137646 560192 137652 560244
rect 137704 560232 137710 560244
rect 140774 560232 140780 560244
rect 137704 560204 140780 560232
rect 137704 560192 137710 560204
rect 140774 560192 140780 560204
rect 140832 560192 140838 560244
rect 204530 560232 204536 560244
rect 142126 560204 204536 560232
rect 106274 560124 106280 560176
rect 106332 560164 106338 560176
rect 124582 560164 124588 560176
rect 106332 560136 124588 560164
rect 106332 560124 106338 560136
rect 124582 560124 124588 560136
rect 124640 560124 124646 560176
rect 134610 560124 134616 560176
rect 134668 560164 134674 560176
rect 142126 560164 142154 560204
rect 204530 560192 204536 560204
rect 204588 560232 204594 560244
rect 302234 560232 302240 560244
rect 204588 560204 302240 560232
rect 204588 560192 204594 560204
rect 302234 560192 302240 560204
rect 302292 560192 302298 560244
rect 134668 560136 142154 560164
rect 134668 560124 134674 560136
rect 98086 560056 98092 560108
rect 98144 560096 98150 560108
rect 122834 560096 122840 560108
rect 98144 560068 122840 560096
rect 98144 560056 98150 560068
rect 122834 560056 122840 560068
rect 122892 560056 122898 560108
rect 96798 559988 96804 560040
rect 96856 560028 96862 560040
rect 124490 560028 124496 560040
rect 96856 560000 124496 560028
rect 96856 559988 96862 560000
rect 124490 559988 124496 560000
rect 124548 559988 124554 560040
rect 164326 559988 164332 560040
rect 164384 560028 164390 560040
rect 200850 560028 200856 560040
rect 164384 560000 200856 560028
rect 164384 559988 164390 560000
rect 200850 559988 200856 560000
rect 200908 559988 200914 560040
rect 93854 559920 93860 559972
rect 93912 559960 93918 559972
rect 124674 559960 124680 559972
rect 93912 559932 124680 559960
rect 93912 559920 93918 559932
rect 124674 559920 124680 559932
rect 124732 559920 124738 559972
rect 182358 559920 182364 559972
rect 182416 559960 182422 559972
rect 218882 559960 218888 559972
rect 182416 559932 218888 559960
rect 182416 559920 182422 559932
rect 218882 559920 218888 559932
rect 218940 559920 218946 559972
rect 260834 559920 260840 559972
rect 260892 559960 260898 559972
rect 316954 559960 316960 559972
rect 260892 559932 316960 559960
rect 260892 559920 260898 559932
rect 316954 559920 316960 559932
rect 317012 559920 317018 559972
rect 57054 559852 57060 559904
rect 57112 559892 57118 559904
rect 67726 559892 67732 559904
rect 57112 559864 67732 559892
rect 57112 559852 57118 559864
rect 67726 559852 67732 559864
rect 67784 559852 67790 559904
rect 86954 559852 86960 559904
rect 87012 559892 87018 559904
rect 120902 559892 120908 559904
rect 87012 559864 120908 559892
rect 87012 559852 87018 559864
rect 120902 559852 120908 559864
rect 120960 559852 120966 559904
rect 137738 559852 137744 559904
rect 137796 559892 137802 559904
rect 145098 559892 145104 559904
rect 137796 559864 145104 559892
rect 137796 559852 137802 559864
rect 145098 559852 145104 559864
rect 145156 559852 145162 559904
rect 157978 559852 157984 559904
rect 158036 559892 158042 559904
rect 203334 559892 203340 559904
rect 158036 559864 203340 559892
rect 158036 559852 158042 559864
rect 203334 559852 203340 559864
rect 203392 559852 203398 559904
rect 258074 559852 258080 559904
rect 258132 559892 258138 559904
rect 316862 559892 316868 559904
rect 258132 559864 316868 559892
rect 258132 559852 258138 559864
rect 316862 559852 316868 559864
rect 316920 559852 316926 559904
rect 59078 559784 59084 559836
rect 59136 559824 59142 559836
rect 82906 559824 82912 559836
rect 59136 559796 82912 559824
rect 59136 559784 59142 559796
rect 82906 559784 82912 559796
rect 82964 559784 82970 559836
rect 87046 559784 87052 559836
rect 87104 559824 87110 559836
rect 121546 559824 121552 559836
rect 87104 559796 121552 559824
rect 87104 559784 87110 559796
rect 121546 559784 121552 559796
rect 121604 559784 121610 559836
rect 139026 559784 139032 559836
rect 139084 559824 139090 559836
rect 150618 559824 150624 559836
rect 139084 559796 150624 559824
rect 139084 559784 139090 559796
rect 150618 559784 150624 559796
rect 150676 559784 150682 559836
rect 154574 559784 154580 559836
rect 154632 559824 154638 559836
rect 201678 559824 201684 559836
rect 154632 559796 201684 559824
rect 154632 559784 154638 559796
rect 201678 559784 201684 559796
rect 201736 559784 201742 559836
rect 216122 559784 216128 559836
rect 216180 559824 216186 559836
rect 282914 559824 282920 559836
rect 216180 559796 282920 559824
rect 216180 559784 216186 559796
rect 282914 559784 282920 559796
rect 282972 559784 282978 559836
rect 54846 559716 54852 559768
rect 54904 559756 54910 559768
rect 78674 559756 78680 559768
rect 54904 559728 78680 559756
rect 54904 559716 54910 559728
rect 78674 559716 78680 559728
rect 78732 559716 78738 559768
rect 85574 559716 85580 559768
rect 85632 559756 85638 559768
rect 121730 559756 121736 559768
rect 85632 559728 121736 559756
rect 85632 559716 85638 559728
rect 121730 559716 121736 559728
rect 121788 559716 121794 559768
rect 134886 559716 134892 559768
rect 134944 559756 134950 559768
rect 151814 559756 151820 559768
rect 134944 559728 151820 559756
rect 134944 559716 134950 559728
rect 151814 559716 151820 559728
rect 151872 559716 151878 559768
rect 156046 559716 156052 559768
rect 156104 559756 156110 559768
rect 204438 559756 204444 559768
rect 156104 559728 204444 559756
rect 156104 559716 156110 559728
rect 204438 559716 204444 559728
rect 204496 559716 204502 559768
rect 247034 559716 247040 559768
rect 247092 559756 247098 559768
rect 319714 559756 319720 559768
rect 247092 559728 319720 559756
rect 247092 559716 247098 559728
rect 319714 559716 319720 559728
rect 319772 559716 319778 559768
rect 67634 559648 67640 559700
rect 67692 559688 67698 559700
rect 121914 559688 121920 559700
rect 67692 559660 121920 559688
rect 67692 559648 67698 559660
rect 121914 559648 121920 559660
rect 121972 559648 121978 559700
rect 136358 559648 136364 559700
rect 136416 559688 136422 559700
rect 161658 559688 161664 559700
rect 136416 559660 161664 559688
rect 136416 559648 136422 559660
rect 161658 559648 161664 559660
rect 161716 559648 161722 559700
rect 179690 559648 179696 559700
rect 179748 559688 179754 559700
rect 281534 559688 281540 559700
rect 179748 559660 281540 559688
rect 179748 559648 179754 559660
rect 281534 559648 281540 559660
rect 281592 559648 281598 559700
rect 63494 559580 63500 559632
rect 63552 559620 63558 559632
rect 122926 559620 122932 559632
rect 63552 559592 122932 559620
rect 63552 559580 63558 559592
rect 122926 559580 122932 559592
rect 122984 559580 122990 559632
rect 138842 559580 138848 559632
rect 138900 559620 138906 559632
rect 165614 559620 165620 559632
rect 138900 559592 165620 559620
rect 138900 559580 138906 559592
rect 165614 559580 165620 559592
rect 165672 559580 165678 559632
rect 180794 559580 180800 559632
rect 180852 559620 180858 559632
rect 283190 559620 283196 559632
rect 180852 559592 283196 559620
rect 180852 559580 180858 559592
rect 283190 559580 283196 559592
rect 283248 559580 283254 559632
rect 3418 559512 3424 559564
rect 3476 559552 3482 559564
rect 286318 559552 286324 559564
rect 3476 559524 286324 559552
rect 3476 559512 3482 559524
rect 286318 559512 286324 559524
rect 286376 559512 286382 559564
rect 217870 559308 217876 559360
rect 217928 559348 217934 559360
rect 222194 559348 222200 559360
rect 217928 559320 222200 559348
rect 217928 559308 217934 559320
rect 222194 559308 222200 559320
rect 222252 559308 222258 559360
rect 219342 559036 219348 559088
rect 219400 559076 219406 559088
rect 223574 559076 223580 559088
rect 219400 559048 223580 559076
rect 219400 559036 219406 559048
rect 223574 559036 223580 559048
rect 223632 559036 223638 559088
rect 139118 558900 139124 558952
rect 139176 558940 139182 558952
rect 142154 558940 142160 558952
rect 139176 558912 142160 558940
rect 139176 558900 139182 558912
rect 142154 558900 142160 558912
rect 142212 558900 142218 558952
rect 57422 558832 57428 558884
rect 57480 558872 57486 558884
rect 60734 558872 60740 558884
rect 57480 558844 60740 558872
rect 57480 558832 57486 558844
rect 60734 558832 60740 558844
rect 60792 558832 60798 558884
rect 100754 558764 100760 558816
rect 100812 558804 100818 558816
rect 102870 558804 102876 558816
rect 100812 558776 102876 558804
rect 100812 558764 100818 558776
rect 102870 558764 102876 558776
rect 102928 558764 102934 558816
rect 116578 558764 116584 558816
rect 116636 558804 116642 558816
rect 120166 558804 120172 558816
rect 116636 558776 120172 558804
rect 116636 558764 116642 558776
rect 120166 558764 120172 558776
rect 120224 558764 120230 558816
rect 161566 558764 161572 558816
rect 161624 558804 161630 558816
rect 168466 558804 168472 558816
rect 161624 558776 168472 558804
rect 161624 558764 161630 558776
rect 168466 558764 168472 558776
rect 168524 558764 168530 558816
rect 173894 558764 173900 558816
rect 173952 558804 173958 558816
rect 179598 558804 179604 558816
rect 173952 558776 179604 558804
rect 173952 558764 173958 558776
rect 179598 558764 179604 558776
rect 179656 558764 179662 558816
rect 225138 558764 225144 558816
rect 225196 558804 225202 558816
rect 227990 558804 227996 558816
rect 225196 558776 227996 558804
rect 225196 558764 225202 558776
rect 227990 558764 227996 558776
rect 228048 558764 228054 558816
rect 260098 558764 260104 558816
rect 260156 558804 260162 558816
rect 262766 558804 262772 558816
rect 260156 558776 262772 558804
rect 260156 558764 260162 558776
rect 262766 558764 262772 558776
rect 262824 558764 262830 558816
rect 278038 558764 278044 558816
rect 278096 558804 278102 558816
rect 280246 558804 280252 558816
rect 278096 558776 280252 558804
rect 278096 558764 278102 558776
rect 280246 558764 280252 558776
rect 280304 558764 280310 558816
rect 60274 558696 60280 558748
rect 60332 558736 60338 558748
rect 62758 558736 62764 558748
rect 60332 558708 62764 558736
rect 60332 558696 60338 558708
rect 62758 558696 62764 558708
rect 62816 558696 62822 558748
rect 119338 558696 119344 558748
rect 119396 558736 119402 558748
rect 120718 558736 120724 558748
rect 119396 558708 120724 558736
rect 119396 558696 119402 558708
rect 120718 558696 120724 558708
rect 120776 558696 120782 558748
rect 147674 558628 147680 558680
rect 147732 558668 147738 558680
rect 162302 558668 162308 558680
rect 147732 558640 162308 558668
rect 147732 558628 147738 558640
rect 162302 558628 162308 558640
rect 162360 558628 162366 558680
rect 151354 558560 151360 558612
rect 151412 558600 151418 558612
rect 164878 558600 164884 558612
rect 151412 558572 164884 558600
rect 151412 558560 151418 558572
rect 164878 558560 164884 558572
rect 164936 558560 164942 558612
rect 231946 558560 231952 558612
rect 232004 558600 232010 558612
rect 259638 558600 259644 558612
rect 232004 558572 259644 558600
rect 232004 558560 232010 558572
rect 259638 558560 259644 558572
rect 259696 558560 259702 558612
rect 142890 558492 142896 558544
rect 142948 558532 142954 558544
rect 160738 558532 160744 558544
rect 142948 558504 160744 558532
rect 142948 558492 142954 558504
rect 160738 558492 160744 558504
rect 160796 558492 160802 558544
rect 222286 558492 222292 558544
rect 222344 558532 222350 558544
rect 253934 558532 253940 558544
rect 222344 558504 253940 558532
rect 222344 558492 222350 558504
rect 253934 558492 253940 558504
rect 253992 558492 253998 558544
rect 68738 558424 68744 558476
rect 68796 558464 68802 558476
rect 71038 558464 71044 558476
rect 68796 558436 71044 558464
rect 68796 558424 68802 558436
rect 71038 558424 71044 558436
rect 71096 558424 71102 558476
rect 82722 558424 82728 558476
rect 82780 558464 82786 558476
rect 88978 558464 88984 558476
rect 82780 558436 88984 558464
rect 82780 558424 82786 558436
rect 88978 558424 88984 558436
rect 89036 558424 89042 558476
rect 140314 558424 140320 558476
rect 140372 558464 140378 558476
rect 159358 558464 159364 558476
rect 140372 558436 159364 558464
rect 140372 558424 140378 558436
rect 159358 558424 159364 558436
rect 159416 558424 159422 558476
rect 188338 558424 188344 558476
rect 188396 558464 188402 558476
rect 200206 558464 200212 558476
rect 188396 558436 200212 558464
rect 188396 558424 188402 558436
rect 200206 558424 200212 558436
rect 200264 558424 200270 558476
rect 212626 558424 212632 558476
rect 212684 558464 212690 558476
rect 251174 558464 251180 558476
rect 212684 558436 251180 558464
rect 212684 558424 212690 558436
rect 251174 558424 251180 558436
rect 251232 558424 251238 558476
rect 77018 558356 77024 558408
rect 77076 558396 77082 558408
rect 85666 558396 85672 558408
rect 77076 558368 85672 558396
rect 77076 558356 77082 558368
rect 85666 558356 85672 558368
rect 85724 558356 85730 558408
rect 94498 558356 94504 558408
rect 94556 558396 94562 558408
rect 104158 558396 104164 558408
rect 94556 558368 104164 558396
rect 94556 558356 94562 558368
rect 104158 558356 104164 558368
rect 104216 558356 104222 558408
rect 112438 558356 112444 558408
rect 112496 558396 112502 558408
rect 117406 558396 117412 558408
rect 112496 558368 117412 558396
rect 112496 558356 112502 558368
rect 117406 558356 117412 558368
rect 117464 558356 117470 558408
rect 129734 558356 129740 558408
rect 129792 558396 129798 558408
rect 153838 558396 153844 558408
rect 129792 558368 153844 558396
rect 129792 558356 129798 558368
rect 153838 558356 153844 558368
rect 153896 558356 153902 558408
rect 154666 558356 154672 558408
rect 154724 558396 154730 558408
rect 171318 558396 171324 558408
rect 154724 558368 171324 558396
rect 154724 558356 154730 558368
rect 171318 558356 171324 558368
rect 171376 558356 171382 558408
rect 187878 558356 187884 558408
rect 187936 558396 187942 558408
rect 233878 558396 233884 558408
rect 187936 558368 233884 558396
rect 187936 558356 187942 558368
rect 233878 558356 233884 558368
rect 233936 558356 233942 558408
rect 62850 558288 62856 558340
rect 62908 558328 62914 558340
rect 80698 558328 80704 558340
rect 62908 558300 80704 558328
rect 62908 558288 62914 558300
rect 80698 558288 80704 558300
rect 80756 558288 80762 558340
rect 86034 558288 86040 558340
rect 86092 558328 86098 558340
rect 108298 558328 108304 558340
rect 86092 558300 108304 558328
rect 86092 558288 86098 558300
rect 108298 558288 108304 558300
rect 108356 558288 108362 558340
rect 111886 558288 111892 558340
rect 111944 558328 111950 558340
rect 123110 558328 123116 558340
rect 111944 558300 123116 558328
rect 111944 558288 111950 558300
rect 123110 558288 123116 558300
rect 123168 558288 123174 558340
rect 133966 558288 133972 558340
rect 134024 558328 134030 558340
rect 197446 558328 197452 558340
rect 134024 558300 197452 558328
rect 134024 558288 134030 558300
rect 197446 558288 197452 558300
rect 197504 558288 197510 558340
rect 227714 558288 227720 558340
rect 227772 558328 227778 558340
rect 245654 558328 245660 558340
rect 227772 558300 245660 558328
rect 227772 558288 227778 558300
rect 245654 558288 245660 558300
rect 245712 558288 245718 558340
rect 249794 558288 249800 558340
rect 249852 558328 249858 558340
rect 294598 558328 294604 558340
rect 249852 558300 294604 558328
rect 249852 558288 249858 558300
rect 294598 558288 294604 558300
rect 294656 558288 294662 558340
rect 71314 558220 71320 558272
rect 71372 558260 71378 558272
rect 93946 558260 93952 558272
rect 71372 558232 93952 558260
rect 71372 558220 71378 558232
rect 93946 558220 93952 558232
rect 94004 558220 94010 558272
rect 100202 558220 100208 558272
rect 100260 558260 100266 558272
rect 115198 558260 115204 558272
rect 100260 558232 115204 558260
rect 100260 558220 100266 558232
rect 115198 558220 115204 558232
rect 115256 558220 115262 558272
rect 118694 558220 118700 558272
rect 118752 558260 118758 558272
rect 144914 558260 144920 558272
rect 118752 558232 144920 558260
rect 118752 558220 118758 558232
rect 144914 558220 144920 558232
rect 144972 558220 144978 558272
rect 158714 558220 158720 558272
rect 158772 558260 158778 558272
rect 182910 558260 182916 558272
rect 158772 558232 182916 558260
rect 158772 558220 158778 558232
rect 182910 558220 182916 558232
rect 182968 558220 182974 558272
rect 190454 558220 190460 558272
rect 190512 558260 190518 558272
rect 257062 558260 257068 558272
rect 190512 558232 257068 558260
rect 190512 558220 190518 558232
rect 257062 558220 257068 558232
rect 257120 558220 257126 558272
rect 273254 558220 273260 558272
rect 273312 558260 273318 558272
rect 318242 558260 318248 558272
rect 273312 558232 318248 558260
rect 273312 558220 273318 558232
rect 318242 558220 318248 558232
rect 318300 558220 318306 558272
rect 58894 558152 58900 558204
rect 58952 558192 58958 558204
rect 74534 558192 74540 558204
rect 58952 558164 74540 558192
rect 58952 558152 58958 558164
rect 74534 558152 74540 558164
rect 74592 558152 74598 558204
rect 79870 558152 79876 558204
rect 79928 558192 79934 558204
rect 114554 558192 114560 558204
rect 79928 558164 114560 558192
rect 79928 558152 79934 558164
rect 114554 558152 114560 558164
rect 114612 558152 114618 558204
rect 132586 558152 132592 558204
rect 132644 558192 132650 558204
rect 177022 558192 177028 558204
rect 132644 558164 177028 558192
rect 132644 558152 132650 558164
rect 177022 558152 177028 558164
rect 177080 558152 177086 558204
rect 177298 558152 177304 558204
rect 177356 558192 177362 558204
rect 188614 558192 188620 558204
rect 177356 558164 188620 558192
rect 177356 558152 177362 558164
rect 188614 558152 188620 558164
rect 188672 558152 188678 558204
rect 191834 558152 191840 558204
rect 191892 558192 191898 558204
rect 276934 558192 276940 558204
rect 191892 558164 276940 558192
rect 191892 558152 191898 558164
rect 276934 558152 276940 558164
rect 276992 558152 276998 558204
rect 71774 557880 71780 557932
rect 71832 557920 71838 557932
rect 73798 557920 73804 557932
rect 71832 557892 73804 557920
rect 71832 557880 71838 557892
rect 73798 557880 73804 557892
rect 73856 557880 73862 557932
rect 184198 557880 184204 557932
rect 184256 557920 184262 557932
rect 185486 557920 185492 557932
rect 184256 557892 185492 557920
rect 184256 557880 184262 557892
rect 185486 557880 185492 557892
rect 185544 557880 185550 557932
rect 264238 557880 264244 557932
rect 264296 557920 264302 557932
rect 265342 557920 265348 557932
rect 264296 557892 265348 557920
rect 264296 557880 264302 557892
rect 265342 557880 265348 557892
rect 265400 557880 265406 557932
rect 262858 557608 262864 557660
rect 262916 557648 262922 557660
rect 268654 557648 268660 557660
rect 262916 557620 268660 557648
rect 262916 557608 262922 557620
rect 268654 557608 268660 557620
rect 268712 557608 268718 557660
rect 64138 557540 64144 557592
rect 64196 557580 64202 557592
rect 65058 557580 65064 557592
rect 64196 557552 65064 557580
rect 64196 557540 64202 557552
rect 65058 557540 65064 557552
rect 65116 557540 65122 557592
rect 222930 557540 222936 557592
rect 222988 557580 222994 557592
rect 224402 557580 224408 557592
rect 222988 557552 224408 557580
rect 222988 557540 222994 557552
rect 224402 557540 224408 557552
rect 224460 557540 224466 557592
rect 267734 557540 267740 557592
rect 267792 557580 267798 557592
rect 317414 557580 317420 557592
rect 267792 557552 317420 557580
rect 267792 557540 267798 557552
rect 317414 557540 317420 557552
rect 317472 557540 317478 557592
rect 219250 557472 219256 557524
rect 219308 557512 219314 557524
rect 223666 557512 223672 557524
rect 219308 557484 223672 557512
rect 219308 557472 219314 557484
rect 223666 557472 223672 557484
rect 223724 557472 223730 557524
rect 178034 557064 178040 557116
rect 178092 557104 178098 557116
rect 206554 557104 206560 557116
rect 178092 557076 206560 557104
rect 178092 557064 178098 557076
rect 206554 557064 206560 557076
rect 206612 557064 206618 557116
rect 269482 557064 269488 557116
rect 269540 557104 269546 557116
rect 300210 557104 300216 557116
rect 269540 557076 300216 557104
rect 269540 557064 269546 557076
rect 300210 557064 300216 557076
rect 300268 557064 300274 557116
rect 57330 556996 57336 557048
rect 57388 557036 57394 557048
rect 81710 557036 81716 557048
rect 57388 557008 81716 557036
rect 57388 556996 57394 557008
rect 81710 556996 81716 557008
rect 81768 556996 81774 557048
rect 122834 556996 122840 557048
rect 122892 557036 122898 557048
rect 202138 557036 202144 557048
rect 122892 557008 202144 557036
rect 122892 556996 122898 557008
rect 202138 556996 202144 557008
rect 202196 556996 202202 557048
rect 229278 556996 229284 557048
rect 229336 557036 229342 557048
rect 281258 557036 281264 557048
rect 229336 557008 281264 557036
rect 229336 556996 229342 557008
rect 281258 556996 281264 557008
rect 281316 556996 281322 557048
rect 78858 556928 78864 556980
rect 78916 556968 78922 556980
rect 121454 556968 121460 556980
rect 78916 556940 121460 556968
rect 78916 556928 78922 556940
rect 121454 556928 121460 556940
rect 121512 556928 121518 556980
rect 143534 556928 143540 556980
rect 143592 556968 143598 556980
rect 156414 556968 156420 556980
rect 143592 556940 156420 556968
rect 143592 556928 143598 556940
rect 156414 556928 156420 556940
rect 156472 556928 156478 556980
rect 159818 556928 159824 556980
rect 159876 556968 159882 556980
rect 173434 556968 173440 556980
rect 159876 556940 173440 556968
rect 159876 556928 159882 556940
rect 173434 556928 173440 556940
rect 173492 556928 173498 556980
rect 194594 556928 194600 556980
rect 194652 556968 194658 556980
rect 283650 556968 283656 556980
rect 194652 556940 283656 556968
rect 194652 556928 194658 556940
rect 283650 556928 283656 556940
rect 283708 556928 283714 556980
rect 63770 556860 63776 556912
rect 63828 556900 63834 556912
rect 123570 556900 123576 556912
rect 63828 556872 123576 556900
rect 63828 556860 63834 556872
rect 123570 556860 123576 556872
rect 123628 556860 123634 556912
rect 138934 556860 138940 556912
rect 138992 556900 138998 556912
rect 160094 556900 160100 556912
rect 138992 556872 160100 556900
rect 138992 556860 138998 556872
rect 160094 556860 160100 556872
rect 160152 556860 160158 556912
rect 179506 556860 179512 556912
rect 179564 556900 179570 556912
rect 281902 556900 281908 556912
rect 179564 556872 281908 556900
rect 179564 556860 179570 556872
rect 281902 556860 281908 556872
rect 281960 556860 281966 556912
rect 4798 556792 4804 556844
rect 4856 556832 4862 556844
rect 318334 556832 318340 556844
rect 4856 556804 318340 556832
rect 4856 556792 4862 556804
rect 318334 556792 318340 556804
rect 318392 556792 318398 556844
rect 219526 556724 219532 556776
rect 219584 556764 219590 556776
rect 219894 556764 219900 556776
rect 219584 556736 219900 556764
rect 219584 556724 219590 556736
rect 219894 556724 219900 556736
rect 219952 556724 219958 556776
rect 193214 555704 193220 555756
rect 193272 555744 193278 555756
rect 218790 555744 218796 555756
rect 193272 555716 218796 555744
rect 193272 555704 193278 555716
rect 218790 555704 218796 555716
rect 218848 555704 218854 555756
rect 266538 555704 266544 555756
rect 266596 555744 266602 555756
rect 307018 555744 307024 555756
rect 266596 555716 307024 555744
rect 266596 555704 266602 555716
rect 307018 555704 307024 555716
rect 307076 555704 307082 555756
rect 168374 555636 168380 555688
rect 168432 555676 168438 555688
rect 200666 555676 200672 555688
rect 168432 555648 200672 555676
rect 168432 555636 168438 555648
rect 200666 555636 200672 555648
rect 200724 555636 200730 555688
rect 240778 555636 240784 555688
rect 240836 555676 240842 555688
rect 283466 555676 283472 555688
rect 240836 555648 283472 555676
rect 240836 555636 240842 555648
rect 283466 555636 283472 555648
rect 283524 555636 283530 555688
rect 59262 555568 59268 555620
rect 59320 555608 59326 555620
rect 92566 555608 92572 555620
rect 59320 555580 92572 555608
rect 59320 555568 59326 555580
rect 92566 555568 92572 555580
rect 92624 555568 92630 555620
rect 100386 555568 100392 555620
rect 100444 555608 100450 555620
rect 123478 555608 123484 555620
rect 100444 555580 123484 555608
rect 100444 555568 100450 555580
rect 123478 555568 123484 555580
rect 123536 555568 123542 555620
rect 137830 555568 137836 555620
rect 137888 555608 137894 555620
rect 149054 555608 149060 555620
rect 137888 555580 149060 555608
rect 137888 555568 137894 555580
rect 149054 555568 149060 555580
rect 149112 555568 149118 555620
rect 157886 555568 157892 555620
rect 157944 555608 157950 555620
rect 203242 555608 203248 555620
rect 157944 555580 203248 555608
rect 157944 555568 157950 555580
rect 203242 555568 203248 555580
rect 203300 555568 203306 555620
rect 245102 555568 245108 555620
rect 245160 555608 245166 555620
rect 318150 555608 318156 555620
rect 245160 555580 318156 555608
rect 245160 555568 245166 555580
rect 318150 555568 318156 555580
rect 318208 555568 318214 555620
rect 64874 555500 64880 555552
rect 64932 555540 64938 555552
rect 122190 555540 122196 555552
rect 64932 555512 122196 555540
rect 64932 555500 64938 555512
rect 122190 555500 122196 555512
rect 122248 555500 122254 555552
rect 138566 555500 138572 555552
rect 138624 555540 138630 555552
rect 169110 555540 169116 555552
rect 138624 555512 169116 555540
rect 138624 555500 138630 555512
rect 169110 555500 169116 555512
rect 169168 555500 169174 555552
rect 181346 555500 181352 555552
rect 181404 555540 181410 555552
rect 281718 555540 281724 555552
rect 181404 555512 281724 555540
rect 181404 555500 181410 555512
rect 281718 555500 281724 555512
rect 281776 555500 281782 555552
rect 3510 555432 3516 555484
rect 3568 555472 3574 555484
rect 319714 555472 319720 555484
rect 3568 555444 319720 555472
rect 3568 555432 3574 555444
rect 319714 555432 319720 555444
rect 319772 555432 319778 555484
rect 129826 554208 129832 554260
rect 129884 554248 129890 554260
rect 202966 554248 202972 554260
rect 129884 554220 202972 554248
rect 129884 554208 129890 554220
rect 202966 554208 202972 554220
rect 203024 554208 203030 554260
rect 246482 554208 246488 554260
rect 246540 554248 246546 554260
rect 287698 554248 287704 554260
rect 246540 554220 287704 554248
rect 246540 554208 246546 554220
rect 287698 554208 287704 554220
rect 287756 554208 287762 554260
rect 73246 554140 73252 554192
rect 73304 554180 73310 554192
rect 108574 554180 108580 554192
rect 73304 554152 108580 554180
rect 73304 554140 73310 554152
rect 108574 554140 108580 554152
rect 108632 554140 108638 554192
rect 122926 554140 122932 554192
rect 122984 554180 122990 554192
rect 201862 554180 201868 554192
rect 122984 554152 201868 554180
rect 122984 554140 122990 554152
rect 201862 554140 201868 554152
rect 201920 554140 201926 554192
rect 263686 554140 263692 554192
rect 263744 554180 263750 554192
rect 315298 554180 315304 554192
rect 263744 554152 315304 554180
rect 263744 554140 263750 554152
rect 315298 554140 315304 554152
rect 315356 554140 315362 554192
rect 58526 554072 58532 554124
rect 58584 554112 58590 554124
rect 110414 554112 110420 554124
rect 58584 554084 110420 554112
rect 58584 554072 58590 554084
rect 110414 554072 110420 554084
rect 110472 554072 110478 554124
rect 195974 554072 195980 554124
rect 196032 554112 196038 554124
rect 283374 554112 283380 554124
rect 196032 554084 283380 554112
rect 196032 554072 196038 554084
rect 283374 554072 283380 554084
rect 283432 554072 283438 554124
rect 66714 554004 66720 554056
rect 66772 554044 66778 554056
rect 121178 554044 121184 554056
rect 66772 554016 121184 554044
rect 66772 554004 66778 554016
rect 121178 554004 121184 554016
rect 121236 554004 121242 554056
rect 182266 554004 182272 554056
rect 182324 554044 182330 554056
rect 281994 554044 282000 554056
rect 182324 554016 282000 554044
rect 182324 554004 182330 554016
rect 281994 554004 282000 554016
rect 282052 554004 282058 554056
rect 3510 553392 3516 553444
rect 3568 553432 3574 553444
rect 317966 553432 317972 553444
rect 3568 553404 317972 553432
rect 3568 553392 3574 553404
rect 317966 553392 317972 553404
rect 318024 553392 318030 553444
rect 226426 552916 226432 552968
rect 226484 552956 226490 552968
rect 280798 552956 280804 552968
rect 226484 552928 280804 552956
rect 226484 552916 226490 552928
rect 280798 552916 280804 552928
rect 280856 552916 280862 552968
rect 59446 552848 59452 552900
rect 59504 552888 59510 552900
rect 75914 552888 75920 552900
rect 59504 552860 75920 552888
rect 59504 552848 59510 552860
rect 75914 552848 75920 552860
rect 75972 552848 75978 552900
rect 88610 552848 88616 552900
rect 88668 552888 88674 552900
rect 103514 552888 103520 552900
rect 88668 552860 103520 552888
rect 88668 552848 88674 552860
rect 103514 552848 103520 552860
rect 103572 552848 103578 552900
rect 106918 552848 106924 552900
rect 106976 552888 106982 552900
rect 123386 552888 123392 552900
rect 106976 552860 123392 552888
rect 106976 552848 106982 552860
rect 123386 552848 123392 552860
rect 123444 552848 123450 552900
rect 128998 552848 129004 552900
rect 129056 552888 129062 552900
rect 203150 552888 203156 552900
rect 129056 552860 203156 552888
rect 129056 552848 129062 552860
rect 203150 552848 203156 552860
rect 203208 552848 203214 552900
rect 256694 552848 256700 552900
rect 256752 552888 256758 552900
rect 316770 552888 316776 552900
rect 256752 552860 316776 552888
rect 256752 552848 256758 552860
rect 316770 552848 316776 552860
rect 316828 552848 316834 552900
rect 75270 552780 75276 552832
rect 75328 552820 75334 552832
rect 96982 552820 96988 552832
rect 75328 552792 96988 552820
rect 75328 552780 75334 552792
rect 96982 552780 96988 552792
rect 97040 552780 97046 552832
rect 121454 552780 121460 552832
rect 121512 552820 121518 552832
rect 201126 552820 201132 552832
rect 121512 552792 201132 552820
rect 121512 552780 121518 552792
rect 201126 552780 201132 552792
rect 201184 552780 201190 552832
rect 250806 552780 250812 552832
rect 250864 552820 250870 552832
rect 319622 552820 319628 552832
rect 250864 552792 319628 552820
rect 250864 552780 250870 552792
rect 319622 552780 319628 552792
rect 319680 552780 319686 552832
rect 57698 552712 57704 552764
rect 57756 552752 57762 552764
rect 77386 552752 77392 552764
rect 57756 552724 77392 552752
rect 57756 552712 57762 552724
rect 77386 552712 77392 552724
rect 77444 552712 77450 552764
rect 80054 552712 80060 552764
rect 80112 552752 80118 552764
rect 120810 552752 120816 552764
rect 80112 552724 120816 552752
rect 80112 552712 80118 552724
rect 120810 552712 120816 552724
rect 120868 552712 120874 552764
rect 138474 552712 138480 552764
rect 138532 552752 138538 552764
rect 160646 552752 160652 552764
rect 138532 552724 160652 552752
rect 138532 552712 138538 552724
rect 160646 552712 160652 552724
rect 160704 552712 160710 552764
rect 196342 552712 196348 552764
rect 196400 552752 196406 552764
rect 283282 552752 283288 552764
rect 196400 552724 283288 552752
rect 196400 552712 196406 552724
rect 283282 552712 283288 552724
rect 283340 552712 283346 552764
rect 69014 552644 69020 552696
rect 69072 552684 69078 552696
rect 114646 552684 114652 552696
rect 69072 552656 114652 552684
rect 69072 552644 69078 552656
rect 114646 552644 114652 552656
rect 114704 552644 114710 552696
rect 138658 552644 138664 552696
rect 138716 552684 138722 552696
rect 174906 552684 174912 552696
rect 138716 552656 174912 552684
rect 138716 552644 138722 552656
rect 174906 552644 174912 552656
rect 174964 552644 174970 552696
rect 179138 552644 179144 552696
rect 179196 552684 179202 552696
rect 271230 552684 271236 552696
rect 179196 552656 271236 552684
rect 179196 552644 179202 552656
rect 271230 552644 271236 552656
rect 271288 552644 271294 552696
rect 192110 551624 192116 551676
rect 192168 551664 192174 551676
rect 217318 551664 217324 551676
rect 192168 551636 217324 551664
rect 192168 551624 192174 551636
rect 217318 551624 217324 551636
rect 217376 551624 217382 551676
rect 281534 551624 281540 551676
rect 281592 551664 281598 551676
rect 293218 551664 293224 551676
rect 281592 551636 293224 551664
rect 281592 551624 281598 551636
rect 293218 551624 293224 551636
rect 293276 551624 293282 551676
rect 176654 551556 176660 551608
rect 176712 551596 176718 551608
rect 210510 551596 210516 551608
rect 176712 551568 210516 551596
rect 176712 551556 176718 551568
rect 210510 551556 210516 551568
rect 210568 551556 210574 551608
rect 260006 551556 260012 551608
rect 260064 551596 260070 551608
rect 289170 551596 289176 551608
rect 260064 551568 289176 551596
rect 260064 551556 260070 551568
rect 289170 551556 289176 551568
rect 289228 551556 289234 551608
rect 80974 551488 80980 551540
rect 81032 551528 81038 551540
rect 122098 551528 122104 551540
rect 81032 551500 122104 551528
rect 81032 551488 81038 551500
rect 122098 551488 122104 551500
rect 122156 551488 122162 551540
rect 144086 551488 144092 551540
rect 144144 551528 144150 551540
rect 201770 551528 201776 551540
rect 144144 551500 201776 551528
rect 144144 551488 144150 551500
rect 201770 551488 201776 551500
rect 201828 551488 201834 551540
rect 253658 551488 253664 551540
rect 253716 551528 253722 551540
rect 316678 551528 316684 551540
rect 253716 551500 316684 551528
rect 253716 551488 253722 551500
rect 316678 551488 316684 551500
rect 316736 551488 316742 551540
rect 57514 551420 57520 551472
rect 57572 551460 57578 551472
rect 89806 551460 89812 551472
rect 57572 551432 89812 551460
rect 57572 551420 57578 551432
rect 89806 551420 89812 551432
rect 89864 551420 89870 551472
rect 93946 551420 93952 551472
rect 94004 551460 94010 551472
rect 114646 551460 114652 551472
rect 94004 551432 114652 551460
rect 94004 551420 94010 551432
rect 114646 551420 114652 551432
rect 114704 551420 114710 551472
rect 121546 551420 121552 551472
rect 121604 551460 121610 551472
rect 201586 551460 201592 551472
rect 121604 551432 201592 551460
rect 121604 551420 121610 551432
rect 201586 551420 201592 551432
rect 201644 551420 201650 551472
rect 211614 551420 211620 551472
rect 211672 551460 211678 551472
rect 280982 551460 280988 551472
rect 211672 551432 280988 551460
rect 211672 551420 211678 551432
rect 280982 551420 280988 551432
rect 281040 551420 281046 551472
rect 282914 551420 282920 551472
rect 282972 551460 282978 551472
rect 304258 551460 304264 551472
rect 282972 551432 304264 551460
rect 282972 551420 282978 551432
rect 304258 551420 304264 551432
rect 304316 551420 304322 551472
rect 58986 551352 58992 551404
rect 59044 551392 59050 551404
rect 102502 551392 102508 551404
rect 59044 551364 102508 551392
rect 59044 551352 59050 551364
rect 102502 551352 102508 551364
rect 102560 551352 102566 551404
rect 200666 551352 200672 551404
rect 200724 551392 200730 551404
rect 281810 551392 281816 551404
rect 200724 551364 281816 551392
rect 200724 551352 200730 551364
rect 281810 551352 281816 551364
rect 281868 551352 281874 551404
rect 65978 551284 65984 551336
rect 66036 551324 66042 551336
rect 123202 551324 123208 551336
rect 66036 551296 123208 551324
rect 66036 551284 66042 551296
rect 123202 551284 123208 551296
rect 123260 551284 123266 551336
rect 139394 551284 139400 551336
rect 139452 551324 139458 551336
rect 159082 551324 159088 551336
rect 139452 551296 159088 551324
rect 139452 551284 139458 551296
rect 159082 551284 159088 551296
rect 159140 551284 159146 551336
rect 186314 551284 186320 551336
rect 186372 551324 186378 551336
rect 283558 551324 283564 551336
rect 186372 551296 283564 551324
rect 186372 551284 186378 551296
rect 283558 551284 283564 551296
rect 283616 551284 283622 551336
rect 176746 550128 176752 550180
rect 176804 550168 176810 550180
rect 225046 550168 225052 550180
rect 176804 550140 225052 550168
rect 176804 550128 176810 550140
rect 225046 550128 225052 550140
rect 225104 550128 225110 550180
rect 228634 550128 228640 550180
rect 228692 550168 228698 550180
rect 280890 550168 280896 550180
rect 228692 550140 280896 550168
rect 228692 550128 228698 550140
rect 280890 550128 280896 550140
rect 280948 550128 280954 550180
rect 80698 550060 80704 550112
rect 80756 550100 80762 550112
rect 109678 550100 109684 550112
rect 80756 550072 109684 550100
rect 80756 550060 80762 550072
rect 109678 550060 109684 550072
rect 109736 550060 109742 550112
rect 142614 550060 142620 550112
rect 142672 550100 142678 550112
rect 202322 550100 202328 550112
rect 142672 550072 202328 550100
rect 142672 550060 142678 550072
rect 202322 550060 202328 550072
rect 202380 550060 202386 550112
rect 251542 550060 251548 550112
rect 251600 550100 251606 550112
rect 313918 550100 313924 550112
rect 251600 550072 313924 550100
rect 251600 550060 251606 550072
rect 313918 550060 313924 550072
rect 313976 550060 313982 550112
rect 59538 549992 59544 550044
rect 59596 550032 59602 550044
rect 101030 550032 101036 550044
rect 59596 550004 101036 550032
rect 59596 549992 59602 550004
rect 101030 549992 101036 550004
rect 101088 549992 101094 550044
rect 120258 549992 120264 550044
rect 120316 550032 120322 550044
rect 190546 550032 190552 550044
rect 120316 550004 190552 550032
rect 120316 549992 120322 550004
rect 190546 549992 190552 550004
rect 190604 549992 190610 550044
rect 193490 549992 193496 550044
rect 193548 550032 193554 550044
rect 213178 550032 213184 550044
rect 193548 550004 213184 550032
rect 193548 549992 193554 550004
rect 213178 549992 213184 550004
rect 213236 549992 213242 550044
rect 242894 549992 242900 550044
rect 242952 550032 242958 550044
rect 314010 550032 314016 550044
rect 242952 550004 314016 550032
rect 242952 549992 242958 550004
rect 314010 549992 314016 550004
rect 314068 549992 314074 550044
rect 69106 549924 69112 549976
rect 69164 549964 69170 549976
rect 120994 549964 121000 549976
rect 69164 549936 121000 549964
rect 69164 549924 69170 549936
rect 120994 549924 121000 549936
rect 121052 549924 121058 549976
rect 138750 549924 138756 549976
rect 138808 549964 138814 549976
rect 153378 549964 153384 549976
rect 138808 549936 153384 549964
rect 138808 549924 138814 549936
rect 153378 549924 153384 549936
rect 153436 549924 153442 549976
rect 189074 549924 189080 549976
rect 189132 549964 189138 549976
rect 262858 549964 262864 549976
rect 189132 549936 262864 549964
rect 189132 549924 189138 549936
rect 262858 549924 262864 549936
rect 262916 549924 262922 549976
rect 271598 549924 271604 549976
rect 271656 549964 271662 549976
rect 289078 549964 289084 549976
rect 271656 549936 289084 549964
rect 271656 549924 271662 549936
rect 289078 549924 289084 549936
rect 289136 549924 289142 549976
rect 70946 549856 70952 549908
rect 71004 549896 71010 549908
rect 121822 549896 121828 549908
rect 71004 549868 121828 549896
rect 71004 549856 71010 549868
rect 121822 549856 121828 549868
rect 121880 549856 121886 549908
rect 147766 549856 147772 549908
rect 147824 549896 147830 549908
rect 167086 549896 167092 549908
rect 147824 549868 167092 549896
rect 147824 549856 147830 549868
rect 167086 549856 167092 549868
rect 167144 549856 167150 549908
rect 187050 549856 187056 549908
rect 187108 549896 187114 549908
rect 283098 549896 283104 549908
rect 187108 549868 283104 549896
rect 187108 549856 187114 549868
rect 283098 549856 283104 549868
rect 283156 549856 283162 549908
rect 40034 549176 40040 549228
rect 40092 549216 40098 549228
rect 317966 549216 317972 549228
rect 40092 549188 317972 549216
rect 40092 549176 40098 549188
rect 317966 549176 317972 549188
rect 318024 549176 318030 549228
rect 199194 548700 199200 548752
rect 199252 548740 199258 548752
rect 215938 548740 215944 548752
rect 199252 548712 215944 548740
rect 199252 548700 199258 548712
rect 215938 548700 215944 548712
rect 215996 548700 216002 548752
rect 88426 548632 88432 548684
rect 88484 548672 88490 548684
rect 104894 548672 104900 548684
rect 88484 548644 104900 548672
rect 88484 548632 88490 548644
rect 104894 548632 104900 548644
rect 104952 548632 104958 548684
rect 189902 548632 189908 548684
rect 189960 548672 189966 548684
rect 206462 548672 206468 548684
rect 189960 548644 206468 548672
rect 189960 548632 189966 548644
rect 206462 548632 206468 548644
rect 206520 548632 206526 548684
rect 76742 548564 76748 548616
rect 76800 548604 76806 548616
rect 112438 548604 112444 548616
rect 76800 548576 112444 548604
rect 76800 548564 76806 548576
rect 112438 548564 112444 548576
rect 112496 548564 112502 548616
rect 205634 548564 205640 548616
rect 205692 548604 205698 548616
rect 264238 548604 264244 548616
rect 205692 548576 264244 548604
rect 205692 548564 205698 548576
rect 264238 548564 264244 548576
rect 264296 548564 264302 548616
rect 59170 548496 59176 548548
rect 59228 548536 59234 548548
rect 108206 548536 108212 548548
rect 59228 548508 108212 548536
rect 59228 548496 59234 548508
rect 108206 548496 108212 548508
rect 108264 548496 108270 548548
rect 136910 548496 136916 548548
rect 136968 548536 136974 548548
rect 201494 548536 201500 548548
rect 136968 548508 201500 548536
rect 136968 548496 136974 548508
rect 201494 548496 201500 548508
rect 201552 548496 201558 548548
rect 210142 548496 210148 548548
rect 210200 548536 210206 548548
rect 281166 548536 281172 548548
rect 210200 548508 281172 548536
rect 210200 548496 210206 548508
rect 281166 548496 281172 548508
rect 281224 548496 281230 548548
rect 57606 547340 57612 547392
rect 57664 547380 57670 547392
rect 91738 547380 91744 547392
rect 57664 547352 91744 547380
rect 57664 547340 57670 547352
rect 91738 547340 91744 547352
rect 91796 547340 91802 547392
rect 140498 547340 140504 547392
rect 140556 547380 140562 547392
rect 188338 547380 188344 547392
rect 140556 547352 188344 547380
rect 140556 547340 140562 547352
rect 188338 547340 188344 547352
rect 188396 547340 188402 547392
rect 190638 547340 190644 547392
rect 190696 547380 190702 547392
rect 204898 547380 204904 547392
rect 190696 547352 204904 547380
rect 190696 547340 190702 547352
rect 204898 547340 204904 547352
rect 204956 547340 204962 547392
rect 211062 547340 211068 547392
rect 211120 547380 211126 547392
rect 235994 547380 236000 547392
rect 211120 547352 236000 547380
rect 211120 547340 211126 547352
rect 235994 547340 236000 547352
rect 236052 547340 236058 547392
rect 259546 547340 259552 547392
rect 259604 547380 259610 547392
rect 309778 547380 309784 547392
rect 259604 547352 309784 547380
rect 259604 547340 259610 547352
rect 309778 547340 309784 547352
rect 309836 547340 309842 547392
rect 84562 547272 84568 547324
rect 84620 547312 84626 547324
rect 122006 547312 122012 547324
rect 84620 547284 122012 547312
rect 84620 547272 84626 547284
rect 122006 547272 122012 547284
rect 122064 547272 122070 547324
rect 124674 547272 124680 547324
rect 124732 547312 124738 547324
rect 201218 547312 201224 547324
rect 124732 547284 201224 547312
rect 124732 547272 124738 547284
rect 201218 547272 201224 547284
rect 201276 547272 201282 547324
rect 235074 547272 235080 547324
rect 235132 547312 235138 547324
rect 319530 547312 319536 547324
rect 235132 547284 319536 547312
rect 235132 547272 235138 547284
rect 319530 547272 319536 547284
rect 319588 547272 319594 547324
rect 62758 547204 62764 547256
rect 62816 547244 62822 547256
rect 105354 547244 105360 547256
rect 62816 547216 105360 547244
rect 62816 547204 62822 547216
rect 105354 547204 105360 547216
rect 105412 547204 105418 547256
rect 185578 547204 185584 547256
rect 185636 547244 185642 547256
rect 274634 547244 274640 547256
rect 185636 547216 274640 547244
rect 185636 547204 185642 547216
rect 274634 547204 274640 547216
rect 274692 547204 274698 547256
rect 63126 547136 63132 547188
rect 63184 547176 63190 547188
rect 110506 547176 110512 547188
rect 63184 547148 110512 547176
rect 63184 547136 63190 547148
rect 110506 547136 110512 547148
rect 110564 547136 110570 547188
rect 122650 547136 122656 547188
rect 122708 547176 122714 547188
rect 137462 547176 137468 547188
rect 122708 547148 137468 547176
rect 122708 547136 122714 547148
rect 137462 547136 137468 547148
rect 137520 547136 137526 547188
rect 147674 547136 147680 547188
rect 147732 547176 147738 547188
rect 184198 547176 184204 547188
rect 147732 547148 184204 547176
rect 147732 547136 147738 547148
rect 184198 547136 184204 547148
rect 184256 547136 184262 547188
rect 187786 547136 187792 547188
rect 187844 547176 187850 547188
rect 283006 547176 283012 547188
rect 187844 547148 283012 547176
rect 187844 547136 187850 547148
rect 283006 547136 283012 547148
rect 283064 547136 283070 547188
rect 273254 547068 273260 547120
rect 273312 547108 273318 547120
rect 274450 547108 274456 547120
rect 273312 547080 274456 547108
rect 273312 547068 273318 547080
rect 274450 547068 274456 547080
rect 274508 547068 274514 547120
rect 139854 546456 139860 546508
rect 139912 546496 139918 546508
rect 141878 546496 141884 546508
rect 139912 546468 141884 546496
rect 139912 546456 139918 546468
rect 141878 546456 141884 546468
rect 141936 546456 141942 546508
rect 184934 545980 184940 546032
rect 184992 546020 184998 546032
rect 216030 546020 216036 546032
rect 184992 545992 216036 546020
rect 184992 545980 184998 545992
rect 216030 545980 216036 545992
rect 216088 545980 216094 546032
rect 138290 545912 138296 545964
rect 138348 545952 138354 545964
rect 200758 545952 200764 545964
rect 138348 545924 200764 545952
rect 138348 545912 138354 545924
rect 200758 545912 200764 545924
rect 200816 545912 200822 545964
rect 206370 545912 206376 545964
rect 206428 545952 206434 545964
rect 241514 545952 241520 545964
rect 206428 545924 241520 545952
rect 206428 545912 206434 545924
rect 241514 545912 241520 545924
rect 241572 545912 241578 545964
rect 267274 545912 267280 545964
rect 267332 545952 267338 545964
rect 300118 545952 300124 545964
rect 267332 545924 300124 545952
rect 267332 545912 267338 545924
rect 300118 545912 300124 545924
rect 300176 545912 300182 545964
rect 82446 545844 82452 545896
rect 82504 545884 82510 545896
rect 116578 545884 116584 545896
rect 82504 545856 116584 545884
rect 82504 545844 82510 545856
rect 116578 545844 116584 545856
rect 116636 545844 116642 545896
rect 139026 545844 139032 545896
rect 139084 545884 139090 545896
rect 202046 545884 202052 545896
rect 139084 545856 202052 545884
rect 139084 545844 139090 545856
rect 202046 545844 202052 545856
rect 202104 545844 202110 545896
rect 217870 545844 217876 545896
rect 217928 545884 217934 545896
rect 260098 545884 260104 545896
rect 217928 545856 260104 545884
rect 217928 545844 217934 545856
rect 260098 545844 260104 545856
rect 260156 545844 260162 545896
rect 275186 545844 275192 545896
rect 275244 545884 275250 545896
rect 312538 545884 312544 545896
rect 275244 545856 312544 545884
rect 275244 545844 275250 545856
rect 312538 545844 312544 545856
rect 312596 545844 312602 545896
rect 57238 545776 57244 545828
rect 57296 545816 57302 545828
rect 103238 545816 103244 545828
rect 57296 545788 103244 545816
rect 57296 545776 57302 545788
rect 103238 545776 103244 545788
rect 103296 545776 103302 545828
rect 198550 545776 198556 545828
rect 198608 545816 198614 545828
rect 278038 545816 278044 545828
rect 198608 545788 278044 545816
rect 198608 545776 198614 545788
rect 278038 545776 278044 545788
rect 278096 545776 278102 545828
rect 71682 545708 71688 545760
rect 71740 545748 71746 545760
rect 123018 545748 123024 545760
rect 71740 545720 123024 545748
rect 71740 545708 71746 545720
rect 123018 545708 123024 545720
rect 123076 545708 123082 545760
rect 127618 545708 127624 545760
rect 127676 545748 127682 545760
rect 194686 545748 194692 545760
rect 127676 545720 194692 545748
rect 127676 545708 127682 545720
rect 194686 545708 194692 545720
rect 194744 545708 194750 545760
rect 197814 545708 197820 545760
rect 197872 545748 197878 545760
rect 210602 545748 210608 545760
rect 197872 545720 210608 545748
rect 197872 545708 197878 545720
rect 210602 545708 210608 545720
rect 210660 545708 210666 545760
rect 234338 545708 234344 545760
rect 234396 545748 234402 545760
rect 319438 545748 319444 545760
rect 234396 545720 319444 545748
rect 234396 545708 234402 545720
rect 319438 545708 319444 545720
rect 319496 545708 319502 545760
rect 289538 545096 289544 545148
rect 289596 545136 289602 545148
rect 313918 545136 313924 545148
rect 289596 545108 313924 545136
rect 289596 545096 289602 545108
rect 313918 545096 313924 545108
rect 313976 545096 313982 545148
rect 154574 544756 154580 544808
rect 154632 544796 154638 544808
rect 155494 544796 155500 544808
rect 154632 544768 155500 544796
rect 154632 544756 154638 544768
rect 155494 544756 155500 544768
rect 155552 544756 155558 544808
rect 171318 544552 171324 544604
rect 171376 544592 171382 544604
rect 203426 544592 203432 544604
rect 171376 544564 203432 544592
rect 171376 544552 171382 544564
rect 203426 544552 203432 544564
rect 203484 544552 203490 544604
rect 161382 544484 161388 544536
rect 161440 544524 161446 544536
rect 203058 544524 203064 544536
rect 161440 544496 203064 544524
rect 161440 544484 161446 544496
rect 203058 544484 203064 544496
rect 203116 544484 203122 544536
rect 219158 544484 219164 544536
rect 219216 544524 219222 544536
rect 227162 544524 227168 544536
rect 219216 544496 227168 544524
rect 219216 544484 219222 544496
rect 227162 544484 227168 544496
rect 227220 544484 227226 544536
rect 270126 544484 270132 544536
rect 270184 544524 270190 544536
rect 287790 544524 287796 544536
rect 270184 544496 287796 544524
rect 270184 544484 270190 544496
rect 287790 544484 287796 544496
rect 287848 544484 287854 544536
rect 94590 544416 94596 544468
rect 94648 544456 94654 544468
rect 123294 544456 123300 544468
rect 94648 544428 123300 544456
rect 94648 544416 94654 544428
rect 123294 544416 123300 544428
rect 123352 544416 123358 544468
rect 137922 544416 137928 544468
rect 137980 544456 137986 544468
rect 149790 544456 149796 544468
rect 137980 544428 149796 544456
rect 137980 544416 137986 544428
rect 149790 544416 149796 544428
rect 149848 544416 149854 544468
rect 152642 544416 152648 544468
rect 152700 544456 152706 544468
rect 201954 544456 201960 544468
rect 152700 544428 201960 544456
rect 152700 544416 152706 544428
rect 201954 544416 201960 544428
rect 202012 544416 202018 544468
rect 220722 544416 220728 544468
rect 220780 544456 220786 544468
rect 247126 544456 247132 544468
rect 220780 544428 247132 544456
rect 220780 544416 220786 544428
rect 247126 544416 247132 544428
rect 247184 544416 247190 544468
rect 279510 544416 279516 544468
rect 279568 544456 279574 544468
rect 311158 544456 311164 544468
rect 279568 544428 311164 544456
rect 279568 544416 279574 544428
rect 311158 544416 311164 544428
rect 311216 544416 311222 544468
rect 71038 544348 71044 544400
rect 71096 544388 71102 544400
rect 108942 544388 108948 544400
rect 71096 544360 108948 544388
rect 71096 544348 71102 544360
rect 108942 544348 108948 544360
rect 109000 544348 109006 544400
rect 131206 544348 131212 544400
rect 131264 544388 131270 544400
rect 177298 544388 177304 544400
rect 131264 544360 177304 544388
rect 131264 544348 131270 544360
rect 177298 544348 177304 544360
rect 177356 544348 177362 544400
rect 184198 544348 184204 544400
rect 184256 544388 184262 544400
rect 281626 544388 281632 544400
rect 184256 544360 281632 544388
rect 184256 544348 184262 544360
rect 281626 544348 281632 544360
rect 281684 544348 281690 544400
rect 290918 544144 290924 544196
rect 290976 544184 290982 544196
rect 290976 544156 296714 544184
rect 290976 544144 290982 544156
rect 287422 544076 287428 544128
rect 287480 544116 287486 544128
rect 287480 544088 295472 544116
rect 287480 544076 287486 544088
rect 69106 544008 69112 544060
rect 69164 544048 69170 544060
rect 70302 544048 70308 544060
rect 69164 544020 70308 544048
rect 69164 544008 69170 544020
rect 70302 544008 70308 544020
rect 70360 544008 70366 544060
rect 104158 544008 104164 544060
rect 104216 544008 104222 544060
rect 113266 544008 113272 544060
rect 113324 544048 113330 544060
rect 121086 544048 121092 544060
rect 113324 544020 121092 544048
rect 113324 544008 113330 544020
rect 121086 544008 121092 544020
rect 121144 544008 121150 544060
rect 121546 544008 121552 544060
rect 121604 544048 121610 544060
rect 122558 544048 122564 544060
rect 121604 544020 122564 544048
rect 121604 544008 121610 544020
rect 122558 544008 122564 544020
rect 122616 544008 122622 544060
rect 63494 543872 63500 543924
rect 63552 543912 63558 543924
rect 64506 543912 64512 543924
rect 63552 543884 64512 543912
rect 63552 543872 63558 543884
rect 64506 543872 64512 543884
rect 64564 543872 64570 543924
rect 78674 543872 78680 543924
rect 78732 543912 78738 543924
rect 79594 543912 79600 543924
rect 78732 543884 79600 543912
rect 78732 543872 78738 543884
rect 79594 543872 79600 543884
rect 79652 543872 79658 543924
rect 88426 543872 88432 543924
rect 88484 543912 88490 543924
rect 89622 543912 89628 543924
rect 88484 543884 89628 543912
rect 88484 543872 88490 543884
rect 89622 543872 89628 543884
rect 89680 543872 89686 543924
rect 89806 543872 89812 543924
rect 89864 543912 89870 543924
rect 91002 543912 91008 543924
rect 89864 543884 91008 543912
rect 89864 543872 89870 543884
rect 91002 543872 91008 543884
rect 91060 543872 91066 543924
rect 100754 543872 100760 543924
rect 100812 543912 100818 543924
rect 101766 543912 101772 543924
rect 100812 543884 101772 543912
rect 100812 543872 100818 543884
rect 101766 543872 101772 543884
rect 101824 543872 101830 543924
rect 61654 543668 61660 543720
rect 61712 543708 61718 543720
rect 64138 543708 64144 543720
rect 61712 543680 64144 543708
rect 61712 543668 61718 543680
rect 64138 543668 64144 543680
rect 64196 543668 64202 543720
rect 88978 543668 88984 543720
rect 89036 543708 89042 543720
rect 90358 543708 90364 543720
rect 89036 543680 90364 543708
rect 89036 543668 89042 543680
rect 90358 543668 90364 543680
rect 90416 543668 90422 543720
rect 104176 543708 104204 544008
rect 291194 543940 291200 543992
rect 291252 543980 291258 543992
rect 292390 543980 292396 543992
rect 291252 543952 292396 543980
rect 291252 543940 291258 543952
rect 292390 543940 292396 543952
rect 292448 543940 292454 543992
rect 293954 543940 293960 543992
rect 294012 543980 294018 543992
rect 295242 543980 295248 543992
rect 294012 543952 295248 543980
rect 294012 543940 294018 543952
rect 295242 543940 295248 543952
rect 295300 543940 295306 543992
rect 295444 543980 295472 544088
rect 296686 544048 296714 544156
rect 314010 544048 314016 544060
rect 296686 544020 314016 544048
rect 314010 544008 314016 544020
rect 314068 544008 314074 544060
rect 314378 543980 314384 543992
rect 295444 543952 314384 543980
rect 314378 543940 314384 543952
rect 314436 543940 314442 543992
rect 106274 543872 106280 543924
rect 106332 543912 106338 543924
rect 107562 543912 107568 543924
rect 106332 543884 107568 543912
rect 106332 543872 106338 543884
rect 107562 543872 107568 543884
rect 107620 543872 107626 543924
rect 114554 543872 114560 543924
rect 114612 543912 114618 543924
rect 115382 543912 115388 543924
rect 114612 543884 115388 543912
rect 114612 543872 114618 543884
rect 115382 543872 115388 543884
rect 115440 543872 115446 543924
rect 124214 543872 124220 543924
rect 124272 543912 124278 543924
rect 125410 543912 125416 543924
rect 124272 543884 125416 543912
rect 124272 543872 124278 543884
rect 125410 543872 125416 543884
rect 125468 543872 125474 543924
rect 125594 543872 125600 543924
rect 125652 543912 125658 543924
rect 126882 543912 126888 543924
rect 125652 543884 126888 543912
rect 125652 543872 125658 543884
rect 126882 543872 126888 543884
rect 126940 543872 126946 543924
rect 129734 543872 129740 543924
rect 129792 543912 129798 543924
rect 130470 543912 130476 543924
rect 129792 543884 130476 543912
rect 129792 543872 129798 543884
rect 130470 543872 130476 543884
rect 130528 543872 130534 543924
rect 136634 543872 136640 543924
rect 136692 543912 136698 543924
rect 137646 543912 137652 543924
rect 136692 543884 137652 543912
rect 136692 543872 136698 543884
rect 137646 543872 137652 543884
rect 137704 543872 137710 543924
rect 142154 543872 142160 543924
rect 142212 543912 142218 543924
rect 143350 543912 143356 543924
rect 142212 543884 143356 543912
rect 142212 543872 142218 543884
rect 143350 543872 143356 543884
rect 143408 543872 143414 543924
rect 143534 543872 143540 543924
rect 143592 543912 143598 543924
rect 144730 543912 144736 543924
rect 143592 543884 144736 543912
rect 143592 543872 143598 543884
rect 144730 543872 144736 543884
rect 144788 543872 144794 543924
rect 158714 543872 158720 543924
rect 158772 543912 158778 543924
rect 159818 543912 159824 543924
rect 158772 543884 159824 543912
rect 158772 543872 158778 543884
rect 159818 543872 159824 543884
rect 159876 543872 159882 543924
rect 161566 543872 161572 543924
rect 161624 543912 161630 543924
rect 162670 543912 162676 543924
rect 161624 543884 162676 543912
rect 161624 543872 161630 543884
rect 162670 543872 162676 543884
rect 162728 543872 162734 543924
rect 164326 543872 164332 543924
rect 164384 543912 164390 543924
rect 165522 543912 165528 543924
rect 164384 543884 165528 543912
rect 164384 543872 164390 543884
rect 165522 543872 165528 543884
rect 165580 543872 165586 543924
rect 179506 543872 179512 543924
rect 179564 543912 179570 543924
rect 180610 543912 180616 543924
rect 179564 543884 180616 543912
rect 179564 543872 179570 543884
rect 180610 543872 180616 543884
rect 180668 543872 180674 543924
rect 180794 543872 180800 543924
rect 180852 543912 180858 543924
rect 181990 543912 181996 543924
rect 180852 543884 181996 543912
rect 180852 543872 180858 543884
rect 181990 543872 181996 543884
rect 182048 543872 182054 543924
rect 191834 543872 191840 543924
rect 191892 543912 191898 543924
rect 192754 543912 192760 543924
rect 191892 543884 192760 543912
rect 191892 543872 191898 543884
rect 192754 543872 192760 543884
rect 192812 543872 192818 543924
rect 193214 543872 193220 543924
rect 193272 543912 193278 543924
rect 194226 543912 194232 543924
rect 193272 543884 194232 543912
rect 193272 543872 193278 543884
rect 194226 543872 194232 543884
rect 194284 543872 194290 543924
rect 195974 543872 195980 543924
rect 196032 543912 196038 543924
rect 197078 543912 197084 543924
rect 196032 543884 197084 543912
rect 196032 543872 196038 543884
rect 197078 543872 197084 543884
rect 197136 543872 197142 543924
rect 208394 543872 208400 543924
rect 208452 543912 208458 543924
rect 209222 543912 209228 543924
rect 208452 543884 209228 543912
rect 208452 543872 208458 543884
rect 209222 543872 209228 543884
rect 209280 543872 209286 543924
rect 212534 543872 212540 543924
rect 212592 543912 212598 543924
rect 213546 543912 213552 543924
rect 212592 543884 213552 543912
rect 212592 543872 212598 543884
rect 213546 543872 213552 543884
rect 213604 543872 213610 543924
rect 213914 543872 213920 543924
rect 213972 543912 213978 543924
rect 215018 543912 215024 543924
rect 213972 543884 215024 543912
rect 213972 543872 213978 543884
rect 215018 543872 215024 543884
rect 215076 543872 215082 543924
rect 222194 543872 222200 543924
rect 222252 543912 222258 543924
rect 222838 543912 222844 543924
rect 222252 543884 222844 543912
rect 222252 543872 222258 543884
rect 222838 543872 222844 543884
rect 222896 543872 222902 543924
rect 256694 543872 256700 543924
rect 256752 543912 256758 543924
rect 257982 543912 257988 543924
rect 256752 543884 257988 543912
rect 256752 543872 256758 543884
rect 257982 543872 257988 543884
rect 258040 543872 258046 543924
rect 285214 543872 285220 543924
rect 285272 543912 285278 543924
rect 314102 543912 314108 543924
rect 285272 543884 314108 543912
rect 285272 543872 285278 543884
rect 314102 543872 314108 543884
rect 314160 543872 314166 543924
rect 137554 543804 137560 543856
rect 137612 543844 137618 543856
rect 139762 543844 139768 543856
rect 137612 543816 139768 543844
rect 137612 543804 137618 543816
rect 139762 543804 139768 543816
rect 139820 543804 139826 543856
rect 252278 543804 252284 543856
rect 252336 543844 252342 543856
rect 317966 543844 317972 543856
rect 252336 543816 317972 543844
rect 252336 543804 252342 543816
rect 317966 543804 317972 543816
rect 318024 543804 318030 543856
rect 237926 543736 237932 543788
rect 237984 543776 237990 543788
rect 316678 543776 316684 543788
rect 237984 543748 316684 543776
rect 237984 543736 237990 543748
rect 316678 543736 316684 543748
rect 316736 543736 316742 543788
rect 106090 543708 106096 543720
rect 104176 543680 106096 543708
rect 106090 543668 106096 543680
rect 106148 543668 106154 543720
rect 108298 543668 108304 543720
rect 108356 543708 108362 543720
rect 111794 543708 111800 543720
rect 108356 543680 111800 543708
rect 108356 543668 108362 543680
rect 111794 543668 111800 543680
rect 111852 543668 111858 543720
rect 115198 543668 115204 543720
rect 115256 543708 115262 543720
rect 116118 543708 116124 543720
rect 115256 543680 116124 543708
rect 115256 543668 115262 543680
rect 116118 543668 116124 543680
rect 116176 543668 116182 543720
rect 135438 543668 135444 543720
rect 135496 543708 135502 543720
rect 137370 543708 137376 543720
rect 135496 543680 137376 543708
rect 135496 543668 135502 543680
rect 137370 543668 137376 543680
rect 137428 543668 137434 543720
rect 146202 543668 146208 543720
rect 146260 543708 146266 543720
rect 146260 543680 200114 543708
rect 146260 543668 146266 543680
rect 55122 543600 55128 543652
rect 55180 543640 55186 543652
rect 67358 543640 67364 543652
rect 55180 543612 67364 543640
rect 55180 543600 55186 543612
rect 67358 543600 67364 543612
rect 67416 543600 67422 543652
rect 91094 543600 91100 543652
rect 91152 543640 91158 543652
rect 96798 543640 96804 543652
rect 91152 543612 96804 543640
rect 91152 543600 91158 543612
rect 96798 543600 96804 543612
rect 96856 543600 96862 543652
rect 134978 543600 134984 543652
rect 135036 543640 135042 543652
rect 146938 543640 146944 543652
rect 135036 543612 146944 543640
rect 135036 543600 135042 543612
rect 146938 543600 146944 543612
rect 146996 543600 147002 543652
rect 159358 543600 159364 543652
rect 159416 543640 159422 543652
rect 163406 543640 163412 543652
rect 159416 543612 163412 543640
rect 159416 543600 159422 543612
rect 163406 543600 163412 543612
rect 163464 543600 163470 543652
rect 165706 543600 165712 543652
rect 165764 543640 165770 543652
rect 169846 543640 169852 543652
rect 165764 543612 169852 543640
rect 165764 543600 165770 543612
rect 169846 543600 169852 543612
rect 169904 543600 169910 543652
rect 200086 543640 200114 543680
rect 201402 543668 201408 543720
rect 201460 543708 201466 543720
rect 206278 543708 206284 543720
rect 201460 543680 206284 543708
rect 201460 543668 201466 543680
rect 206278 543668 206284 543680
rect 206336 543668 206342 543720
rect 207106 543668 207112 543720
rect 207164 543708 207170 543720
rect 209038 543708 209044 543720
rect 207164 543680 209044 543708
rect 207164 543668 207170 543680
rect 209038 543668 209044 543680
rect 209096 543668 209102 543720
rect 217226 543668 217232 543720
rect 217284 543708 217290 543720
rect 218606 543708 218612 543720
rect 217284 543680 218612 543708
rect 217284 543668 217290 543680
rect 218606 543668 218612 543680
rect 218664 543668 218670 543720
rect 219526 543668 219532 543720
rect 219584 543708 219590 543720
rect 221458 543708 221464 543720
rect 219584 543680 221464 543708
rect 219584 543668 219590 543680
rect 221458 543668 221464 543680
rect 221516 543668 221522 543720
rect 224402 543668 224408 543720
rect 224460 543708 224466 543720
rect 225782 543708 225788 543720
rect 224460 543680 225788 543708
rect 224460 543668 224466 543680
rect 225782 543668 225788 543680
rect 225840 543668 225846 543720
rect 202230 543640 202236 543652
rect 200086 543612 202236 543640
rect 202230 543600 202236 543612
rect 202288 543600 202294 543652
rect 203518 543600 203524 543652
rect 203576 543640 203582 543652
rect 211798 543640 211804 543652
rect 203576 543612 211804 543640
rect 203576 543600 203582 543612
rect 211798 543600 211804 543612
rect 211856 543600 211862 543652
rect 217594 543600 217600 543652
rect 217652 543640 217658 543652
rect 219250 543640 219256 543652
rect 217652 543612 219256 543640
rect 217652 543600 217658 543612
rect 219250 543600 219256 543612
rect 219308 543600 219314 543652
rect 55030 543532 55036 543584
rect 55088 543572 55094 543584
rect 88886 543572 88892 543584
rect 55088 543544 88892 543572
rect 55088 543532 55094 543544
rect 88886 543532 88892 543544
rect 88944 543532 88950 543584
rect 96062 543532 96068 543584
rect 96120 543572 96126 543584
rect 106918 543572 106924 543584
rect 96120 543544 106924 543572
rect 96120 543532 96126 543544
rect 106918 543532 106924 543544
rect 106976 543532 106982 543584
rect 118234 543532 118240 543584
rect 118292 543572 118298 543584
rect 126238 543572 126244 543584
rect 118292 543544 126244 543572
rect 118292 543532 118298 543544
rect 126238 543532 126244 543544
rect 126296 543532 126302 543584
rect 131850 543532 131856 543584
rect 131908 543572 131914 543584
rect 133138 543572 133144 543584
rect 131908 543544 133144 543572
rect 131908 543532 131914 543544
rect 133138 543532 133144 543544
rect 133196 543532 133202 543584
rect 135162 543532 135168 543584
rect 135220 543572 135226 543584
rect 151262 543572 151268 543584
rect 135220 543544 151268 543572
rect 135220 543532 135226 543544
rect 151262 543532 151268 543544
rect 151320 543532 151326 543584
rect 164878 543532 164884 543584
rect 164936 543572 164942 543584
rect 172698 543572 172704 543584
rect 164936 543544 172704 543572
rect 164936 543532 164942 543544
rect 172698 543532 172704 543544
rect 172756 543532 172762 543584
rect 57790 543464 57796 543516
rect 57848 543504 57854 543516
rect 93210 543504 93216 543516
rect 57848 543476 93216 543504
rect 57848 543464 57854 543476
rect 93210 543464 93216 543476
rect 93268 543464 93274 543516
rect 110414 543464 110420 543516
rect 110472 543504 110478 543516
rect 119338 543504 119344 543516
rect 110472 543476 119344 543504
rect 110472 543464 110478 543476
rect 119338 543464 119344 543476
rect 119396 543464 119402 543516
rect 120442 543464 120448 543516
rect 120500 543504 120506 543516
rect 122650 543504 122656 543516
rect 120500 543476 122656 543504
rect 120500 543464 120506 543476
rect 122650 543464 122656 543476
rect 122708 543464 122714 543516
rect 136542 543464 136548 543516
rect 136600 543504 136606 543516
rect 157702 543504 157708 543516
rect 136600 543476 157708 543504
rect 136600 543464 136606 543476
rect 157702 543464 157708 543476
rect 157760 543464 157766 543516
rect 237190 543464 237196 543516
rect 237248 543504 237254 543516
rect 284294 543504 284300 543516
rect 237248 543476 284300 543504
rect 237248 543464 237254 543476
rect 284294 543464 284300 543476
rect 284352 543464 284358 543516
rect 58710 543396 58716 543448
rect 58768 543436 58774 543448
rect 95326 543436 95332 543448
rect 58768 543408 95332 543436
rect 58768 543396 58774 543408
rect 95326 543396 95332 543408
rect 95384 543396 95390 543448
rect 114002 543396 114008 543448
rect 114060 543436 114066 543448
rect 124398 543436 124404 543448
rect 114060 543408 124404 543436
rect 114060 543396 114066 543408
rect 124398 543396 124404 543408
rect 124456 543396 124462 543448
rect 135070 543396 135076 543448
rect 135128 543436 135134 543448
rect 156966 543436 156972 543448
rect 135128 543408 156972 543436
rect 135128 543396 135134 543408
rect 156966 543396 156972 543408
rect 157024 543396 157030 543448
rect 164142 543396 164148 543448
rect 164200 543436 164206 543448
rect 173986 543436 173992 543448
rect 164200 543408 173992 543436
rect 164200 543396 164206 543408
rect 173986 543396 173992 543408
rect 174044 543396 174050 543448
rect 277302 543396 277308 543448
rect 277360 543436 277366 543448
rect 303062 543436 303068 543448
rect 277360 543408 303068 543436
rect 277360 543396 277366 543408
rect 303062 543396 303068 543408
rect 303120 543396 303126 543448
rect 56502 543328 56508 543380
rect 56560 543368 56566 543380
rect 83918 543368 83924 543380
rect 56560 543340 83924 543368
rect 56560 543328 56566 543340
rect 83918 543328 83924 543340
rect 83976 543328 83982 543380
rect 85298 543328 85304 543380
rect 85356 543368 85362 543380
rect 121914 543368 121920 543380
rect 85356 543340 121920 543368
rect 85356 543328 85362 543340
rect 121914 543328 121920 543340
rect 121972 543328 121978 543380
rect 139302 543328 139308 543380
rect 139360 543368 139366 543380
rect 164878 543368 164884 543380
rect 139360 543340 164884 543368
rect 139360 543328 139366 543340
rect 164878 543328 164884 543340
rect 164936 543328 164942 543380
rect 199930 543328 199936 543380
rect 199988 543368 199994 543380
rect 210418 543368 210424 543380
rect 199988 543340 210424 543368
rect 199988 543328 199994 543340
rect 210418 543328 210424 543340
rect 210476 543328 210482 543380
rect 252922 543328 252928 543380
rect 252980 543368 252986 543380
rect 301774 543368 301780 543380
rect 252980 543340 301780 543368
rect 252980 543328 252986 543340
rect 301774 543328 301780 543340
rect 301832 543328 301838 543380
rect 56410 543260 56416 543312
rect 56468 543300 56474 543312
rect 99650 543300 99656 543312
rect 56468 543272 99656 543300
rect 56468 543260 56474 543272
rect 99650 543260 99656 543272
rect 99708 543260 99714 543312
rect 106826 543260 106832 543312
rect 106884 543300 106890 543312
rect 125686 543300 125692 543312
rect 106884 543272 125692 543300
rect 106884 543260 106890 543272
rect 125686 543260 125692 543272
rect 125744 543260 125750 543312
rect 139210 543260 139216 543312
rect 139268 543300 139274 543312
rect 175550 543300 175556 543312
rect 139268 543272 175556 543300
rect 139268 543260 139274 543272
rect 175550 543260 175556 543272
rect 175608 543260 175614 543312
rect 195606 543260 195612 543312
rect 195664 543300 195670 543312
rect 206462 543300 206468 543312
rect 195664 543272 206468 543300
rect 195664 543260 195670 543272
rect 206462 543260 206468 543272
rect 206520 543260 206526 543312
rect 242250 543260 242256 543312
rect 242308 543300 242314 543312
rect 301590 543300 301596 543312
rect 242308 543272 301596 543300
rect 242308 543260 242314 543272
rect 301590 543260 301596 543272
rect 301648 543260 301654 543312
rect 54938 543192 54944 543244
rect 54996 543232 55002 543244
rect 98914 543232 98920 543244
rect 54996 543204 98920 543232
rect 54996 543192 55002 543204
rect 98914 543192 98920 543204
rect 98972 543192 98978 543244
rect 103974 543192 103980 543244
rect 104032 543232 104038 543244
rect 104032 543204 118096 543232
rect 104032 543192 104038 543204
rect 56318 543124 56324 543176
rect 56376 543164 56382 543176
rect 73798 543164 73804 543176
rect 56376 543136 73804 543164
rect 56376 543124 56382 543136
rect 73798 543124 73804 543136
rect 73856 543124 73862 543176
rect 78122 543124 78128 543176
rect 78180 543164 78186 543176
rect 78180 543136 117728 543164
rect 78180 543124 78186 543136
rect 58802 543056 58808 543108
rect 58860 543096 58866 543108
rect 116854 543096 116860 543108
rect 58860 543068 116860 543096
rect 58860 543056 58866 543068
rect 116854 543056 116860 543068
rect 116912 543056 116918 543108
rect 58618 542988 58624 543040
rect 58676 543028 58682 543040
rect 117590 543028 117596 543040
rect 58676 543000 117596 543028
rect 58676 542988 58682 543000
rect 117590 542988 117596 543000
rect 117648 542988 117654 543040
rect 117700 542960 117728 543136
rect 118068 543028 118096 543204
rect 128262 543192 128268 543244
rect 128320 543232 128326 543244
rect 157978 543232 157984 543244
rect 128320 543204 157984 543232
rect 128320 543192 128326 543204
rect 157978 543192 157984 543204
rect 158036 543192 158042 543244
rect 160738 543192 160744 543244
rect 160796 543232 160802 543244
rect 167730 543232 167736 543244
rect 160796 543204 167736 543232
rect 160796 543192 160802 543204
rect 167730 543192 167736 543204
rect 167788 543192 167794 543244
rect 170582 543192 170588 543244
rect 170640 543232 170646 543244
rect 201034 543232 201040 543244
rect 170640 543204 201040 543232
rect 170640 543192 170646 543204
rect 201034 543192 201040 543204
rect 201092 543192 201098 543244
rect 202138 543192 202144 543244
rect 202196 543232 202202 543244
rect 216122 543232 216128 543244
rect 202196 543204 216128 543232
rect 202196 543192 202202 543204
rect 216122 543192 216128 543204
rect 216180 543192 216186 543244
rect 217962 543192 217968 543244
rect 218020 543232 218026 543244
rect 230014 543232 230020 543244
rect 218020 543204 230020 543232
rect 218020 543192 218026 543204
rect 230014 543192 230020 543204
rect 230072 543192 230078 543244
rect 231486 543192 231492 543244
rect 231544 543232 231550 543244
rect 238754 543232 238760 543244
rect 231544 543204 238760 543232
rect 231544 543192 231550 543204
rect 238754 543192 238760 543204
rect 238812 543192 238818 543244
rect 278038 543192 278044 543244
rect 278096 543232 278102 543244
rect 319622 543232 319628 543244
rect 278096 543204 319628 543232
rect 278096 543192 278102 543204
rect 319622 543192 319628 543204
rect 319680 543192 319686 543244
rect 136450 543124 136456 543176
rect 136508 543164 136514 543176
rect 171962 543164 171968 543176
rect 136508 543136 171968 543164
rect 136508 543124 136514 543136
rect 171962 543124 171968 543136
rect 172020 543124 172026 543176
rect 176286 543124 176292 543176
rect 176344 543164 176350 543176
rect 214558 543164 214564 543176
rect 176344 543136 214564 543164
rect 176344 543124 176350 543136
rect 214558 543124 214564 543136
rect 214616 543124 214622 543176
rect 220078 543124 220084 543176
rect 220136 543164 220142 543176
rect 232866 543164 232872 543176
rect 220136 543136 232872 543164
rect 220136 543124 220142 543136
rect 232866 543124 232872 543136
rect 232924 543124 232930 543176
rect 238662 543124 238668 543176
rect 238720 543164 238726 543176
rect 319438 543164 319444 543176
rect 238720 543136 319444 543164
rect 238720 543124 238726 543136
rect 319438 543124 319444 543136
rect 319496 543124 319502 543176
rect 118970 543056 118976 543108
rect 119028 543096 119034 543108
rect 134518 543096 134524 543108
rect 119028 543068 134524 543096
rect 119028 543056 119034 543068
rect 134518 543056 134524 543068
rect 134576 543056 134582 543108
rect 202782 543056 202788 543108
rect 202840 543096 202846 543108
rect 211062 543096 211068 543108
rect 202840 543068 211068 543096
rect 202840 543056 202846 543068
rect 211062 543056 211068 543068
rect 211120 543056 211126 543108
rect 216398 543056 216404 543108
rect 216456 543096 216462 543108
rect 240778 543096 240784 543108
rect 216456 543068 240784 543096
rect 216456 543056 216462 543068
rect 240778 543056 240784 543068
rect 240836 543056 240842 543108
rect 245838 543056 245844 543108
rect 245896 543096 245902 543108
rect 281074 543096 281080 543108
rect 245896 543068 281080 543096
rect 245896 543056 245902 543068
rect 281074 543056 281080 543068
rect 281132 543056 281138 543108
rect 124306 543028 124312 543040
rect 118068 543000 124312 543028
rect 124306 542988 124312 543000
rect 124364 542988 124370 543040
rect 126146 542988 126152 543040
rect 126204 543028 126210 543040
rect 200942 543028 200948 543040
rect 126204 543000 200948 543028
rect 126204 542988 126210 543000
rect 200942 542988 200948 543000
rect 201000 542988 201006 543040
rect 218698 542988 218704 543040
rect 218756 543028 218762 543040
rect 233602 543028 233608 543040
rect 218756 543000 233608 543028
rect 218756 542988 218762 543000
rect 233602 542988 233608 543000
rect 233660 542988 233666 543040
rect 284938 543028 284944 543040
rect 240796 543000 284944 543028
rect 240796 542972 240824 543000
rect 284938 542988 284944 543000
rect 284996 542988 285002 543040
rect 299566 542988 299572 543040
rect 299624 543028 299630 543040
rect 318058 543028 318064 543040
rect 299624 543000 318064 543028
rect 299624 542988 299630 543000
rect 318058 542988 318064 543000
rect 318116 542988 318122 543040
rect 122190 542960 122196 542972
rect 117700 542932 122196 542960
rect 122190 542920 122196 542932
rect 122248 542920 122254 542972
rect 240778 542920 240784 542972
rect 240836 542920 240842 542972
rect 275922 542920 275928 542972
rect 275980 542960 275986 542972
rect 301958 542960 301964 542972
rect 275980 542932 301964 542960
rect 275980 542920 275986 542932
rect 301958 542920 301964 542932
rect 302016 542920 302022 542972
rect 270862 542852 270868 542904
rect 270920 542892 270926 542904
rect 300578 542892 300584 542904
rect 270920 542864 300584 542892
rect 270920 542852 270926 542864
rect 300578 542852 300584 542864
rect 300636 542852 300642 542904
rect 273714 542784 273720 542836
rect 273772 542824 273778 542836
rect 304258 542824 304264 542836
rect 273772 542796 304264 542824
rect 273772 542784 273778 542796
rect 304258 542784 304264 542796
rect 304316 542784 304322 542836
rect 276566 542716 276572 542768
rect 276624 542756 276630 542768
rect 318150 542756 318156 542768
rect 276624 542728 318156 542756
rect 276624 542716 276630 542728
rect 318150 542716 318156 542728
rect 318208 542716 318214 542768
rect 257246 542648 257252 542700
rect 257304 542688 257310 542700
rect 300394 542688 300400 542700
rect 257304 542660 300400 542688
rect 257304 542648 257310 542660
rect 300394 542648 300400 542660
rect 300452 542648 300458 542700
rect 283098 542580 283104 542632
rect 283156 542620 283162 542632
rect 300118 542620 300124 542632
rect 283156 542592 300124 542620
rect 283156 542580 283162 542592
rect 300118 542580 300124 542592
rect 300176 542580 300182 542632
rect 284478 542512 284484 542564
rect 284536 542552 284542 542564
rect 301682 542552 301688 542564
rect 284536 542524 301688 542552
rect 284536 542512 284542 542524
rect 301682 542512 301688 542524
rect 301740 542512 301746 542564
rect 280154 542444 280160 542496
rect 280212 542484 280218 542496
rect 301866 542484 301872 542496
rect 280212 542456 301872 542484
rect 280212 542444 280218 542456
rect 301866 542444 301872 542456
rect 301924 542444 301930 542496
rect 154114 542376 154120 542428
rect 154172 542416 154178 542428
rect 161382 542416 161388 542428
rect 154172 542388 161388 542416
rect 154172 542376 154178 542388
rect 161382 542376 161388 542388
rect 161440 542376 161446 542428
rect 296714 542376 296720 542428
rect 296772 542416 296778 542428
rect 302878 542416 302884 542428
rect 296772 542388 302884 542416
rect 296772 542376 296778 542388
rect 302878 542376 302884 542388
rect 302936 542376 302942 542428
rect 292546 541980 302234 542008
rect 235810 541832 235816 541884
rect 235868 541872 235874 541884
rect 292546 541872 292574 541980
rect 302050 541872 302056 541884
rect 235868 541844 292574 541872
rect 297376 541844 302056 541872
rect 235868 541832 235874 541844
rect 268746 541764 268752 541816
rect 268804 541804 268810 541816
rect 297376 541804 297404 541844
rect 302050 541832 302056 541844
rect 302108 541832 302114 541884
rect 302206 541872 302234 541980
rect 319530 541872 319536 541884
rect 302206 541844 319536 541872
rect 319530 541832 319536 541844
rect 319588 541832 319594 541884
rect 268804 541776 297404 541804
rect 268804 541764 268810 541776
rect 298094 541764 298100 541816
rect 298152 541804 298158 541816
rect 298830 541804 298836 541816
rect 298152 541776 298836 541804
rect 298152 541764 298158 541776
rect 298830 541764 298836 541776
rect 298888 541764 298894 541816
rect 281626 541696 281632 541748
rect 281684 541736 281690 541748
rect 316862 541736 316868 541748
rect 281684 541708 316868 541736
rect 281684 541696 281690 541708
rect 316862 541696 316868 541708
rect 316920 541696 316926 541748
rect 265894 541628 265900 541680
rect 265952 541668 265958 541680
rect 300302 541668 300308 541680
rect 265952 541640 300308 541668
rect 265952 541628 265958 541640
rect 300302 541628 300308 541640
rect 300360 541628 300366 541680
rect 260834 541560 260840 541612
rect 260892 541600 260898 541612
rect 317138 541600 317144 541612
rect 260892 541572 317144 541600
rect 260892 541560 260898 541572
rect 317138 541560 317144 541572
rect 317196 541560 317202 541612
rect 243630 541492 243636 541544
rect 243688 541532 243694 541544
rect 300670 541532 300676 541544
rect 243688 541504 300676 541532
rect 243688 541492 243694 541504
rect 300670 541492 300676 541504
rect 300728 541492 300734 541544
rect 244366 541424 244372 541476
rect 244424 541464 244430 541476
rect 302970 541464 302976 541476
rect 244424 541436 302976 541464
rect 244424 541424 244430 541436
rect 302970 541424 302976 541436
rect 303028 541424 303034 541476
rect 255866 541356 255872 541408
rect 255924 541396 255930 541408
rect 317966 541396 317972 541408
rect 255924 541368 317972 541396
rect 255924 541356 255930 541368
rect 317966 541356 317972 541368
rect 318024 541356 318030 541408
rect 240042 541288 240048 541340
rect 240100 541328 240106 541340
rect 303154 541328 303160 541340
rect 240100 541300 303160 541328
rect 240100 541288 240106 541300
rect 303154 541288 303160 541300
rect 303212 541288 303218 541340
rect 254394 541220 254400 541272
rect 254452 541260 254458 541272
rect 319806 541260 319812 541272
rect 254452 541232 319812 541260
rect 254452 541220 254458 541232
rect 319806 541220 319812 541232
rect 319864 541220 319870 541272
rect 236454 541152 236460 541204
rect 236512 541192 236518 541204
rect 304350 541192 304356 541204
rect 236512 541164 304356 541192
rect 236512 541152 236518 541164
rect 304350 541152 304356 541164
rect 304408 541152 304414 541204
rect 319622 541152 319628 541204
rect 319680 541192 319686 541204
rect 319680 541164 319852 541192
rect 319680 541152 319686 541164
rect 319824 541136 319852 541164
rect 249426 541084 249432 541136
rect 249484 541124 249490 541136
rect 318334 541124 318340 541136
rect 249484 541096 318340 541124
rect 249484 541084 249490 541096
rect 318334 541084 318340 541096
rect 318392 541084 318398 541136
rect 319806 541084 319812 541136
rect 319864 541084 319870 541136
rect 247218 541016 247224 541068
rect 247276 541056 247282 541068
rect 319622 541056 319628 541068
rect 247276 541028 319628 541056
rect 247276 541016 247282 541028
rect 319622 541016 319628 541028
rect 319680 541016 319686 541068
rect 272334 540948 272340 541000
rect 272392 540988 272398 541000
rect 300486 540988 300492 541000
rect 272392 540960 300492 540988
rect 272392 540948 272398 540960
rect 300486 540948 300492 540960
rect 300544 540948 300550 541000
rect 295978 540744 295984 540796
rect 296036 540784 296042 540796
rect 296036 540756 306374 540784
rect 296036 540744 296042 540756
rect 306346 540648 306374 540756
rect 317230 540648 317236 540660
rect 306346 540620 317236 540648
rect 317230 540608 317236 540620
rect 317288 540608 317294 540660
rect 293770 540540 293776 540592
rect 293828 540580 293834 540592
rect 314286 540580 314292 540592
rect 293828 540552 314292 540580
rect 293828 540540 293834 540552
rect 314286 540540 314292 540552
rect 314344 540540 314350 540592
rect 293126 540472 293132 540524
rect 293184 540512 293190 540524
rect 314470 540512 314476 540524
rect 293184 540484 314476 540512
rect 293184 540472 293190 540484
rect 314470 540472 314476 540484
rect 314528 540472 314534 540524
rect 278774 540404 278780 540456
rect 278832 540444 278838 540456
rect 300854 540444 300860 540456
rect 278832 540416 300860 540444
rect 278832 540404 278838 540416
rect 300854 540404 300860 540416
rect 300912 540404 300918 540456
rect 265158 540336 265164 540388
rect 265216 540376 265222 540388
rect 318794 540376 318800 540388
rect 265216 540348 318800 540376
rect 265216 540336 265222 540348
rect 318794 540336 318800 540348
rect 318852 540336 318858 540388
rect 263042 540268 263048 540320
rect 263100 540308 263106 540320
rect 307018 540308 307024 540320
rect 263100 540280 307024 540308
rect 263100 540268 263106 540280
rect 307018 540268 307024 540280
rect 307076 540268 307082 540320
rect 273070 540200 273076 540252
rect 273128 540240 273134 540252
rect 319346 540240 319352 540252
rect 273128 540212 319352 540240
rect 273128 540200 273134 540212
rect 319346 540200 319352 540212
rect 319404 540200 319410 540252
rect 262306 540132 262312 540184
rect 262364 540172 262370 540184
rect 318426 540172 318432 540184
rect 262364 540144 318432 540172
rect 262364 540132 262370 540144
rect 318426 540132 318432 540144
rect 318484 540132 318490 540184
rect 3602 540064 3608 540116
rect 3660 540104 3666 540116
rect 312538 540104 312544 540116
rect 3660 540076 312544 540104
rect 3660 540064 3666 540076
rect 312538 540064 312544 540076
rect 312596 540064 312602 540116
rect 300854 539520 300860 539572
rect 300912 539560 300918 539572
rect 318058 539560 318064 539572
rect 300912 539532 318064 539560
rect 300912 539520 300918 539532
rect 318058 539520 318064 539532
rect 318116 539520 318122 539572
rect 304350 535372 304356 535424
rect 304408 535412 304414 535424
rect 317598 535412 317604 535424
rect 304408 535384 317604 535412
rect 304408 535372 304414 535384
rect 317598 535372 317604 535384
rect 317656 535372 317662 535424
rect 302326 532176 302332 532228
rect 302384 532216 302390 532228
rect 304350 532216 304356 532228
rect 302384 532188 304356 532216
rect 302384 532176 302390 532188
rect 304350 532176 304356 532188
rect 304408 532176 304414 532228
rect 300670 529864 300676 529916
rect 300728 529904 300734 529916
rect 317598 529904 317604 529916
rect 300728 529876 317604 529904
rect 300728 529864 300734 529876
rect 317598 529864 317604 529876
rect 317656 529864 317662 529916
rect 303154 525716 303160 525768
rect 303212 525756 303218 525768
rect 317690 525756 317696 525768
rect 303212 525728 317696 525756
rect 303212 525716 303218 525728
rect 317690 525716 317696 525728
rect 317748 525716 317754 525768
rect 431218 525240 431224 525292
rect 431276 525280 431282 525292
rect 431402 525280 431408 525292
rect 431276 525252 431408 525280
rect 431276 525240 431282 525252
rect 431402 525240 431408 525252
rect 431460 525240 431466 525292
rect 430942 525104 430948 525156
rect 431000 525144 431006 525156
rect 431218 525144 431224 525156
rect 431000 525116 431224 525144
rect 431000 525104 431006 525116
rect 431218 525104 431224 525116
rect 431276 525104 431282 525156
rect 430666 524968 430672 525020
rect 430724 525008 430730 525020
rect 430942 525008 430948 525020
rect 430724 524980 430948 525008
rect 430724 524968 430730 524980
rect 430942 524968 430948 524980
rect 431000 524968 431006 525020
rect 319346 524696 319352 524748
rect 319404 524696 319410 524748
rect 319364 524544 319392 524696
rect 319346 524492 319352 524544
rect 319404 524492 319410 524544
rect 319438 524424 319444 524476
rect 319496 524464 319502 524476
rect 319806 524464 319812 524476
rect 319496 524436 319812 524464
rect 319496 524424 319502 524436
rect 319806 524424 319812 524436
rect 319864 524424 319870 524476
rect 319162 523676 319168 523728
rect 319220 523716 319226 523728
rect 319622 523716 319628 523728
rect 319220 523688 319628 523716
rect 319220 523676 319226 523688
rect 319622 523676 319628 523688
rect 319680 523676 319686 523728
rect 318794 520684 318800 520736
rect 318852 520724 318858 520736
rect 319898 520724 319904 520736
rect 318852 520696 319904 520724
rect 318852 520684 318858 520696
rect 319898 520684 319904 520696
rect 319956 520684 319962 520736
rect 314378 520208 314384 520260
rect 314436 520248 314442 520260
rect 476114 520248 476120 520260
rect 314436 520220 476120 520248
rect 314436 520208 314442 520220
rect 476114 520208 476120 520220
rect 476172 520208 476178 520260
rect 317230 520140 317236 520192
rect 317288 520180 317294 520192
rect 457438 520180 457444 520192
rect 317288 520152 457444 520180
rect 317288 520140 317294 520152
rect 457438 520140 457444 520152
rect 457496 520140 457502 520192
rect 300578 520072 300584 520124
rect 300636 520112 300642 520124
rect 430850 520112 430856 520124
rect 300636 520084 430856 520112
rect 300636 520072 300642 520084
rect 430850 520072 430856 520084
rect 430908 520072 430914 520124
rect 300394 520004 300400 520056
rect 300452 520044 300458 520056
rect 431310 520044 431316 520056
rect 300452 520016 431316 520044
rect 300452 520004 300458 520016
rect 431310 520004 431316 520016
rect 431368 520004 431374 520056
rect 301866 519936 301872 519988
rect 301924 519976 301930 519988
rect 430666 519976 430672 519988
rect 301924 519948 430672 519976
rect 301924 519936 301930 519948
rect 430666 519936 430672 519948
rect 430724 519936 430730 519988
rect 303062 519868 303068 519920
rect 303120 519908 303126 519920
rect 431218 519908 431224 519920
rect 303120 519880 431224 519908
rect 303120 519868 303126 519880
rect 431218 519868 431224 519880
rect 431276 519868 431282 519920
rect 319254 519800 319260 519852
rect 319312 519840 319318 519852
rect 430942 519840 430948 519852
rect 319312 519812 430948 519840
rect 319312 519800 319318 519812
rect 430942 519800 430948 519812
rect 431000 519800 431006 519852
rect 319438 519732 319444 519784
rect 319496 519772 319502 519784
rect 431402 519772 431408 519784
rect 319496 519744 431408 519772
rect 319496 519732 319502 519744
rect 431402 519732 431408 519744
rect 431460 519732 431466 519784
rect 301958 519188 301964 519240
rect 302016 519228 302022 519240
rect 351270 519228 351276 519240
rect 302016 519200 351276 519228
rect 302016 519188 302022 519200
rect 351270 519188 351276 519200
rect 351328 519188 351334 519240
rect 305638 519120 305644 519172
rect 305696 519160 305702 519172
rect 369302 519160 369308 519172
rect 305696 519132 369308 519160
rect 305696 519120 305702 519132
rect 369302 519120 369308 519132
rect 369360 519120 369366 519172
rect 304258 519052 304264 519104
rect 304316 519092 304322 519104
rect 396902 519092 396908 519104
rect 304316 519064 396908 519092
rect 304316 519052 304322 519064
rect 396902 519052 396908 519064
rect 396960 519052 396966 519104
rect 318150 518984 318156 519036
rect 318208 519024 318214 519036
rect 414934 519024 414940 519036
rect 318208 518996 414940 519024
rect 318208 518984 318214 518996
rect 414934 518984 414940 518996
rect 414992 518984 414998 519036
rect 324866 518916 324872 518968
rect 324924 518956 324930 518968
rect 429194 518956 429200 518968
rect 324924 518928 429200 518956
rect 324924 518916 324930 518928
rect 429194 518916 429200 518928
rect 429252 518916 429258 518968
rect 319806 518848 319812 518900
rect 319864 518888 319870 518900
rect 346670 518888 346676 518900
rect 319864 518860 346676 518888
rect 319864 518848 319870 518860
rect 346670 518848 346676 518860
rect 346728 518848 346734 518900
rect 319530 518780 319536 518832
rect 319588 518820 319594 518832
rect 333238 518820 333244 518832
rect 319588 518792 333244 518820
rect 319588 518780 319594 518792
rect 333238 518780 333244 518792
rect 333296 518780 333302 518832
rect 318426 518712 318432 518764
rect 318484 518752 318490 518764
rect 328730 518752 328736 518764
rect 318484 518724 328736 518752
rect 318484 518712 318490 518724
rect 328730 518712 328736 518724
rect 328788 518712 328794 518764
rect 318334 518644 318340 518696
rect 318392 518684 318398 518696
rect 423950 518684 423956 518696
rect 318392 518656 423956 518684
rect 318392 518644 318398 518656
rect 423950 518644 423956 518656
rect 424008 518644 424014 518696
rect 307018 518576 307024 518628
rect 307076 518616 307082 518628
rect 401594 518616 401600 518628
rect 307076 518588 401600 518616
rect 307076 518576 307082 518588
rect 401594 518576 401600 518588
rect 401652 518576 401658 518628
rect 318058 518508 318064 518560
rect 318116 518548 318122 518560
rect 406010 518548 406016 518560
rect 318116 518520 406016 518548
rect 318116 518508 318122 518520
rect 406010 518508 406016 518520
rect 406068 518508 406074 518560
rect 302050 518440 302056 518492
rect 302108 518480 302114 518492
rect 387886 518480 387892 518492
rect 302108 518452 387892 518480
rect 302108 518440 302114 518452
rect 387886 518440 387892 518452
rect 387944 518440 387950 518492
rect 300302 518372 300308 518424
rect 300360 518412 300366 518424
rect 383654 518412 383660 518424
rect 300360 518384 383660 518412
rect 300360 518372 300366 518384
rect 383654 518372 383660 518384
rect 383712 518372 383718 518424
rect 319346 518304 319352 518356
rect 319404 518344 319410 518356
rect 364702 518344 364708 518356
rect 319404 518316 364708 518344
rect 319404 518304 319410 518316
rect 364702 518304 364708 518316
rect 364760 518304 364766 518356
rect 319162 518236 319168 518288
rect 319220 518276 319226 518288
rect 360286 518276 360292 518288
rect 319220 518248 360292 518276
rect 319220 518236 319226 518248
rect 360286 518236 360292 518248
rect 360344 518236 360350 518288
rect 317138 518168 317144 518220
rect 317196 518208 317202 518220
rect 342254 518208 342260 518220
rect 317196 518180 342260 518208
rect 317196 518168 317202 518180
rect 342254 518168 342260 518180
rect 342312 518168 342318 518220
rect 301774 518100 301780 518152
rect 301832 518140 301838 518152
rect 431126 518140 431132 518152
rect 301832 518112 431132 518140
rect 301832 518100 301838 518112
rect 431126 518100 431132 518112
rect 431184 518100 431190 518152
rect 302970 518032 302976 518084
rect 303028 518072 303034 518084
rect 419534 518072 419540 518084
rect 303028 518044 419540 518072
rect 303028 518032 303034 518044
rect 419534 518032 419540 518044
rect 419592 518032 419598 518084
rect 300486 517964 300492 518016
rect 300544 518004 300550 518016
rect 410518 518004 410524 518016
rect 300544 517976 410524 518004
rect 300544 517964 300550 517976
rect 410518 517964 410524 517976
rect 410576 517964 410582 518016
rect 314470 517420 314476 517472
rect 314528 517460 314534 517472
rect 512270 517460 512276 517472
rect 314528 517432 512276 517460
rect 314528 517420 314534 517432
rect 512270 517420 512276 517432
rect 512328 517420 512334 517472
rect 317046 517352 317052 517404
rect 317104 517392 317110 517404
rect 495434 517392 495440 517404
rect 317104 517364 495440 517392
rect 317104 517352 317110 517364
rect 495434 517352 495440 517364
rect 495492 517352 495498 517404
rect 302878 517284 302884 517336
rect 302936 517324 302942 517336
rect 459554 517324 459560 517336
rect 302936 517296 459560 517324
rect 302936 517284 302942 517296
rect 459554 517284 459560 517296
rect 459612 517284 459618 517336
rect 314194 517216 314200 517268
rect 314252 517256 314258 517268
rect 457714 517256 457720 517268
rect 314252 517228 457720 517256
rect 314252 517216 314258 517228
rect 457714 517216 457720 517228
rect 457772 517216 457778 517268
rect 300118 517148 300124 517200
rect 300176 517188 300182 517200
rect 430574 517188 430580 517200
rect 300176 517160 430580 517188
rect 300176 517148 300182 517160
rect 430574 517148 430580 517160
rect 430632 517148 430638 517200
rect 301590 517080 301596 517132
rect 301648 517120 301654 517132
rect 431034 517120 431040 517132
rect 301648 517092 431040 517120
rect 301648 517080 301654 517092
rect 431034 517080 431040 517092
rect 431092 517080 431098 517132
rect 301682 517012 301688 517064
rect 301740 517052 301746 517064
rect 430758 517052 430764 517064
rect 301740 517024 430764 517052
rect 301740 517012 301746 517024
rect 430758 517012 430764 517024
rect 430816 517012 430822 517064
rect 302602 516128 302608 516180
rect 302660 516168 302666 516180
rect 519538 516168 519544 516180
rect 302660 516140 519544 516168
rect 302660 516128 302666 516140
rect 519538 516128 519544 516140
rect 519596 516128 519602 516180
rect 301498 516060 301504 516112
rect 301556 516100 301562 516112
rect 512178 516100 512184 516112
rect 301556 516072 512184 516100
rect 301556 516060 301562 516072
rect 512178 516060 512184 516072
rect 512236 516060 512242 516112
rect 316954 515992 316960 516044
rect 317012 516032 317018 516044
rect 500954 516032 500960 516044
rect 317012 516004 500960 516032
rect 317012 515992 317018 516004
rect 500954 515992 500960 516004
rect 501012 515992 501018 516044
rect 314010 515924 314016 515976
rect 314068 515964 314074 515976
rect 488534 515964 488540 515976
rect 314068 515936 488540 515964
rect 314068 515924 314074 515936
rect 488534 515924 488540 515936
rect 488592 515924 488598 515976
rect 314102 515856 314108 515908
rect 314160 515896 314166 515908
rect 470594 515896 470600 515908
rect 314160 515868 470600 515896
rect 314160 515856 314166 515868
rect 470594 515856 470600 515868
rect 470652 515856 470658 515908
rect 314286 515788 314292 515840
rect 314344 515828 314350 515840
rect 465074 515828 465080 515840
rect 314344 515800 465080 515828
rect 314344 515788 314350 515800
rect 465074 515788 465080 515800
rect 465132 515788 465138 515840
rect 313918 515720 313924 515772
rect 313976 515760 313982 515772
rect 457622 515760 457628 515772
rect 313976 515732 457628 515760
rect 313976 515720 313982 515732
rect 457622 515720 457628 515732
rect 457680 515720 457686 515772
rect 316862 515652 316868 515704
rect 316920 515692 316926 515704
rect 429470 515692 429476 515704
rect 316920 515664 429476 515692
rect 316920 515652 316926 515664
rect 429470 515652 429476 515664
rect 429528 515652 429534 515704
rect 304350 515380 304356 515432
rect 304408 515420 304414 515432
rect 580258 515420 580264 515432
rect 304408 515392 580264 515420
rect 304408 515380 304414 515392
rect 580258 515380 580264 515392
rect 580316 515380 580322 515432
rect 316678 514700 316684 514752
rect 316736 514740 316742 514752
rect 428366 514740 428372 514752
rect 316736 514712 428372 514740
rect 316736 514700 316742 514712
rect 428366 514700 428372 514712
rect 428424 514700 428430 514752
rect 316770 514632 316776 514684
rect 316828 514672 316834 514684
rect 427814 514672 427820 514684
rect 316828 514644 427820 514672
rect 316828 514632 316834 514644
rect 427814 514632 427820 514644
rect 427872 514632 427878 514684
rect 560938 511912 560944 511964
rect 560996 511952 561002 511964
rect 580166 511952 580172 511964
rect 560996 511924 580172 511952
rect 560996 511912 561002 511924
rect 580166 511912 580172 511924
rect 580224 511912 580230 511964
rect 42702 509872 42708 509924
rect 42760 509912 42766 509924
rect 57698 509912 57704 509924
rect 42760 509884 57704 509912
rect 42760 509872 42766 509884
rect 57698 509872 57704 509884
rect 57756 509872 57762 509924
rect 302878 487160 302884 487212
rect 302936 487200 302942 487212
rect 520918 487200 520924 487212
rect 302936 487172 520924 487200
rect 302936 487160 302942 487172
rect 520918 487160 520924 487172
rect 520976 487160 520982 487212
rect 158714 480020 158720 480072
rect 158772 480060 158778 480072
rect 158990 480060 158996 480072
rect 158772 480032 158996 480060
rect 158772 480020 158778 480032
rect 158990 480020 158996 480032
rect 159048 480020 159054 480072
rect 187786 480020 187792 480072
rect 187844 480060 187850 480072
rect 188062 480060 188068 480072
rect 187844 480032 188068 480060
rect 187844 480020 187850 480032
rect 188062 480020 188068 480032
rect 188120 480020 188126 480072
rect 248414 480020 248420 480072
rect 248472 480060 248478 480072
rect 248782 480060 248788 480072
rect 248472 480032 248788 480060
rect 248472 480020 248478 480032
rect 248782 480020 248788 480032
rect 248840 480020 248846 480072
rect 161490 479816 161496 479868
rect 161548 479856 161554 479868
rect 162026 479856 162032 479868
rect 161548 479828 162032 479856
rect 161548 479816 161554 479828
rect 162026 479816 162032 479828
rect 162084 479816 162090 479868
rect 223590 479816 223596 479868
rect 223648 479856 223654 479868
rect 223758 479856 223764 479868
rect 223648 479828 223764 479856
rect 223648 479816 223654 479828
rect 223758 479816 223764 479828
rect 223816 479816 223822 479868
rect 295350 479816 295356 479868
rect 295408 479856 295414 479868
rect 295978 479856 295984 479868
rect 295408 479828 295984 479856
rect 295408 479816 295414 479828
rect 295978 479816 295984 479828
rect 296036 479816 296042 479868
rect 50982 478932 50988 478984
rect 51040 478972 51046 478984
rect 84378 478972 84384 478984
rect 51040 478944 84384 478972
rect 51040 478932 51046 478944
rect 84378 478932 84384 478944
rect 84436 478932 84442 478984
rect 140774 478932 140780 478984
rect 140832 478972 140838 478984
rect 197722 478972 197728 478984
rect 140832 478944 197728 478972
rect 140832 478932 140838 478944
rect 197722 478932 197728 478944
rect 197780 478932 197786 478984
rect 52086 478864 52092 478916
rect 52144 478904 52150 478916
rect 99374 478904 99380 478916
rect 52144 478876 99380 478904
rect 52144 478864 52150 478876
rect 99374 478864 99380 478876
rect 99432 478864 99438 478916
rect 109494 478864 109500 478916
rect 109552 478904 109558 478916
rect 207106 478904 207112 478916
rect 109552 478876 207112 478904
rect 109552 478864 109558 478876
rect 207106 478864 207112 478876
rect 207164 478864 207170 478916
rect 54570 478796 54576 478848
rect 54628 478836 54634 478848
rect 63678 478836 63684 478848
rect 54628 478808 63684 478836
rect 54628 478796 54634 478808
rect 63678 478796 63684 478808
rect 63736 478796 63742 478848
rect 68278 478796 68284 478848
rect 68336 478836 68342 478848
rect 91830 478836 91836 478848
rect 68336 478808 91836 478836
rect 68336 478796 68342 478808
rect 91830 478796 91836 478808
rect 91888 478796 91894 478848
rect 149974 478796 149980 478848
rect 150032 478836 150038 478848
rect 212534 478836 212540 478848
rect 150032 478808 212540 478836
rect 150032 478796 150038 478808
rect 212534 478796 212540 478808
rect 212592 478796 212598 478848
rect 236270 478796 236276 478848
rect 236328 478836 236334 478848
rect 357434 478836 357440 478848
rect 236328 478808 357440 478836
rect 236328 478796 236334 478808
rect 357434 478796 357440 478808
rect 357492 478796 357498 478848
rect 50890 478728 50896 478780
rect 50948 478768 50954 478780
rect 73154 478768 73160 478780
rect 50948 478740 73160 478768
rect 50948 478728 50954 478740
rect 73154 478728 73160 478740
rect 73212 478728 73218 478780
rect 156138 478728 156144 478780
rect 156196 478768 156202 478780
rect 213914 478768 213920 478780
rect 156196 478740 213920 478768
rect 156196 478728 156202 478740
rect 213914 478728 213920 478740
rect 213972 478728 213978 478780
rect 56410 478660 56416 478712
rect 56468 478700 56474 478712
rect 81710 478700 81716 478712
rect 56468 478672 81716 478700
rect 56468 478660 56474 478672
rect 81710 478660 81716 478672
rect 81768 478660 81774 478712
rect 149514 478660 149520 478712
rect 149572 478700 149578 478712
rect 205634 478700 205640 478712
rect 149572 478672 205640 478700
rect 149572 478660 149578 478672
rect 205634 478660 205640 478672
rect 205692 478660 205698 478712
rect 50062 478592 50068 478644
rect 50120 478632 50126 478644
rect 77294 478632 77300 478644
rect 50120 478604 77300 478632
rect 50120 478592 50126 478604
rect 77294 478592 77300 478604
rect 77352 478592 77358 478644
rect 153470 478592 153476 478644
rect 153528 478632 153534 478644
rect 208486 478632 208492 478644
rect 153528 478604 208492 478632
rect 153528 478592 153534 478604
rect 208486 478592 208492 478604
rect 208544 478592 208550 478644
rect 59170 478524 59176 478576
rect 59228 478564 59234 478576
rect 91002 478564 91008 478576
rect 59228 478536 91008 478564
rect 59228 478524 59234 478536
rect 91002 478524 91008 478536
rect 91060 478524 91066 478576
rect 152182 478524 152188 478576
rect 152240 478564 152246 478576
rect 204346 478564 204352 478576
rect 152240 478536 204352 478564
rect 152240 478524 152246 478536
rect 204346 478524 204352 478536
rect 204404 478524 204410 478576
rect 239398 478524 239404 478576
rect 239456 478564 239462 478576
rect 356698 478564 356704 478576
rect 239456 478536 356704 478564
rect 239456 478524 239462 478536
rect 356698 478524 356704 478536
rect 356756 478524 356762 478576
rect 52822 478456 52828 478508
rect 52880 478496 52886 478508
rect 74258 478496 74264 478508
rect 52880 478468 74264 478496
rect 52880 478456 52886 478468
rect 74258 478456 74264 478468
rect 74316 478456 74322 478508
rect 74350 478456 74356 478508
rect 74408 478496 74414 478508
rect 105078 478496 105084 478508
rect 74408 478468 105084 478496
rect 74408 478456 74414 478468
rect 105078 478456 105084 478468
rect 105136 478456 105142 478508
rect 154850 478456 154856 478508
rect 154908 478496 154914 478508
rect 205634 478496 205640 478508
rect 154908 478468 205640 478496
rect 154908 478456 154914 478468
rect 205634 478456 205640 478468
rect 205692 478456 205698 478508
rect 240226 478456 240232 478508
rect 240284 478496 240290 478508
rect 358354 478496 358360 478508
rect 240284 478468 358360 478496
rect 240284 478456 240290 478468
rect 358354 478456 358360 478468
rect 358412 478456 358418 478508
rect 56318 478388 56324 478440
rect 56376 478428 56382 478440
rect 89162 478428 89168 478440
rect 56376 478400 89168 478428
rect 56376 478388 56382 478400
rect 89162 478388 89168 478400
rect 89220 478388 89226 478440
rect 151262 478388 151268 478440
rect 151320 478428 151326 478440
rect 200666 478428 200672 478440
rect 151320 478400 200672 478428
rect 151320 478388 151326 478400
rect 200666 478388 200672 478400
rect 200724 478388 200730 478440
rect 239858 478388 239864 478440
rect 239916 478428 239922 478440
rect 358262 478428 358268 478440
rect 239916 478400 358268 478428
rect 239916 478388 239922 478400
rect 358262 478388 358268 478400
rect 358320 478388 358326 478440
rect 53466 478320 53472 478372
rect 53524 478360 53530 478372
rect 73154 478360 73160 478372
rect 53524 478332 73160 478360
rect 53524 478320 53530 478332
rect 73154 478320 73160 478332
rect 73212 478320 73218 478372
rect 73890 478320 73896 478372
rect 73948 478360 73954 478372
rect 110322 478360 110328 478372
rect 73948 478332 110328 478360
rect 73948 478320 73954 478332
rect 110322 478320 110328 478332
rect 110380 478320 110386 478372
rect 149146 478320 149152 478372
rect 149204 478360 149210 478372
rect 197354 478360 197360 478372
rect 149204 478332 197360 478360
rect 149204 478320 149210 478332
rect 197354 478320 197360 478332
rect 197412 478320 197418 478372
rect 232774 478320 232780 478372
rect 232832 478360 232838 478372
rect 366450 478360 366456 478372
rect 232832 478332 366456 478360
rect 232832 478320 232838 478332
rect 366450 478320 366456 478332
rect 366508 478320 366514 478372
rect 51994 478252 52000 478304
rect 52052 478292 52058 478304
rect 100202 478292 100208 478304
rect 52052 478264 100208 478292
rect 52052 478252 52058 478264
rect 100202 478252 100208 478264
rect 100260 478252 100266 478304
rect 157058 478252 157064 478304
rect 157116 478292 157122 478304
rect 200114 478292 200120 478304
rect 157116 478264 200120 478292
rect 157116 478252 157122 478264
rect 200114 478252 200120 478264
rect 200172 478252 200178 478304
rect 200206 478252 200212 478304
rect 200264 478292 200270 478304
rect 217502 478292 217508 478304
rect 200264 478264 217508 478292
rect 200264 478252 200270 478264
rect 217502 478252 217508 478264
rect 217560 478252 217566 478304
rect 224402 478252 224408 478304
rect 224460 478292 224466 478304
rect 362218 478292 362224 478304
rect 224460 478264 362224 478292
rect 224460 478252 224466 478264
rect 362218 478252 362224 478264
rect 362276 478252 362282 478304
rect 62758 478184 62764 478236
rect 62816 478224 62822 478236
rect 116302 478224 116308 478236
rect 62816 478196 116308 478224
rect 62816 478184 62822 478196
rect 116302 478184 116308 478196
rect 116360 478184 116366 478236
rect 158346 478184 158352 478236
rect 158404 478224 158410 478236
rect 201494 478224 201500 478236
rect 158404 478196 201500 478224
rect 158404 478184 158410 478196
rect 201494 478184 201500 478196
rect 201552 478184 201558 478236
rect 205450 478184 205456 478236
rect 205508 478224 205514 478236
rect 221734 478224 221740 478236
rect 205508 478196 221740 478224
rect 205508 478184 205514 478196
rect 221734 478184 221740 478196
rect 221792 478184 221798 478236
rect 225690 478184 225696 478236
rect 225748 478224 225754 478236
rect 363598 478224 363604 478236
rect 225748 478196 363604 478224
rect 225748 478184 225754 478196
rect 363598 478184 363604 478196
rect 363656 478184 363662 478236
rect 43806 478116 43812 478168
rect 43864 478156 43870 478168
rect 102410 478156 102416 478168
rect 43864 478128 102416 478156
rect 43864 478116 43870 478128
rect 102410 478116 102416 478128
rect 102468 478116 102474 478168
rect 138934 478116 138940 478168
rect 138992 478156 138998 478168
rect 185578 478156 185584 478168
rect 138992 478128 185584 478156
rect 138992 478116 138998 478128
rect 185578 478116 185584 478128
rect 185636 478116 185642 478168
rect 198458 478116 198464 478168
rect 198516 478156 198522 478168
rect 217318 478156 217324 478168
rect 198516 478128 217324 478156
rect 198516 478116 198522 478128
rect 217318 478116 217324 478128
rect 217376 478116 217382 478168
rect 225322 478116 225328 478168
rect 225380 478156 225386 478168
rect 373258 478156 373264 478168
rect 225380 478128 373264 478156
rect 225380 478116 225386 478128
rect 373258 478116 373264 478128
rect 373316 478116 373322 478168
rect 64138 478048 64144 478100
rect 64196 478088 64202 478100
rect 72418 478088 72424 478100
rect 64196 478060 72424 478088
rect 64196 478048 64202 478060
rect 72418 478048 72424 478060
rect 72476 478048 72482 478100
rect 74074 478048 74080 478100
rect 74132 478088 74138 478100
rect 95326 478088 95332 478100
rect 74132 478060 95332 478088
rect 74132 478048 74138 478060
rect 95326 478048 95332 478060
rect 95384 478048 95390 478100
rect 166258 478048 166264 478100
rect 166316 478088 166322 478100
rect 204898 478088 204904 478100
rect 166316 478060 204904 478088
rect 166316 478048 166322 478060
rect 204898 478048 204904 478060
rect 204956 478048 204962 478100
rect 74166 477980 74172 478032
rect 74224 478020 74230 478032
rect 94958 478020 94964 478032
rect 74224 477992 94964 478020
rect 74224 477980 74230 477992
rect 94958 477980 94964 477992
rect 95016 477980 95022 478032
rect 139394 477980 139400 478032
rect 139452 478020 139458 478032
rect 169018 478020 169024 478032
rect 139452 477992 169024 478020
rect 139452 477980 139458 477992
rect 169018 477980 169024 477992
rect 169076 477980 169082 478032
rect 186130 477980 186136 478032
rect 186188 478020 186194 478032
rect 186498 478020 186504 478032
rect 186188 477992 186504 478020
rect 186188 477980 186194 477992
rect 186498 477980 186504 477992
rect 186556 477980 186562 478032
rect 186958 477980 186964 478032
rect 187016 478020 187022 478032
rect 197998 478020 198004 478032
rect 187016 477992 198004 478020
rect 187016 477980 187022 477992
rect 197998 477980 198004 477992
rect 198056 477980 198062 478032
rect 73982 477912 73988 477964
rect 74040 477952 74046 477964
rect 91370 477952 91376 477964
rect 74040 477924 91376 477952
rect 74040 477912 74046 477924
rect 91370 477912 91376 477924
rect 91428 477912 91434 477964
rect 71314 477844 71320 477896
rect 71372 477884 71378 477896
rect 84838 477884 84844 477896
rect 71372 477856 84844 477884
rect 71372 477844 71378 477856
rect 84838 477844 84844 477856
rect 84896 477844 84902 477896
rect 195330 477572 195336 477624
rect 195388 477612 195394 477624
rect 199378 477612 199384 477624
rect 195388 477584 199384 477612
rect 195388 477572 195394 477584
rect 199378 477572 199384 477584
rect 199436 477572 199442 477624
rect 73798 477504 73804 477556
rect 73856 477544 73862 477556
rect 74350 477544 74356 477556
rect 73856 477516 74356 477544
rect 73856 477504 73862 477516
rect 74350 477504 74356 477516
rect 74408 477504 74414 477556
rect 194870 477504 194876 477556
rect 194928 477544 194934 477556
rect 196986 477544 196992 477556
rect 194928 477516 196992 477544
rect 194928 477504 194934 477516
rect 196986 477504 196992 477516
rect 197044 477504 197050 477556
rect 209406 477504 209412 477556
rect 209464 477544 209470 477556
rect 210326 477544 210332 477556
rect 209464 477516 210332 477544
rect 209464 477504 209470 477516
rect 210326 477504 210332 477516
rect 210384 477504 210390 477556
rect 212074 477504 212080 477556
rect 212132 477544 212138 477556
rect 215938 477544 215944 477556
rect 212132 477516 215944 477544
rect 212132 477504 212138 477516
rect 215938 477504 215944 477516
rect 215996 477504 216002 477556
rect 217410 477504 217416 477556
rect 217468 477544 217474 477556
rect 219710 477544 219716 477556
rect 217468 477516 219716 477544
rect 217468 477504 217474 477516
rect 219710 477504 219716 477516
rect 219768 477504 219774 477556
rect 219986 477504 219992 477556
rect 220044 477544 220050 477556
rect 222654 477544 222660 477556
rect 220044 477516 222660 477544
rect 220044 477504 220050 477516
rect 222654 477504 222660 477516
rect 222712 477504 222718 477556
rect 283006 477436 283012 477488
rect 283064 477476 283070 477488
rect 359826 477476 359832 477488
rect 283064 477448 359832 477476
rect 283064 477436 283070 477448
rect 359826 477436 359832 477448
rect 359884 477436 359890 477488
rect 294414 477368 294420 477420
rect 294472 477408 294478 477420
rect 375190 477408 375196 477420
rect 294472 477380 375196 477408
rect 294472 477368 294478 477380
rect 375190 477368 375196 477380
rect 375248 477368 375254 477420
rect 275922 477300 275928 477352
rect 275980 477340 275986 477352
rect 377306 477340 377312 477352
rect 275980 477312 377312 477340
rect 275980 477300 275986 477312
rect 377306 477300 377312 477312
rect 377364 477300 377370 477352
rect 254762 477232 254768 477284
rect 254820 477272 254826 477284
rect 356790 477272 356796 477284
rect 254820 477244 356796 477272
rect 254820 477232 254826 477244
rect 356790 477232 356796 477244
rect 356848 477232 356854 477284
rect 267550 477164 267556 477216
rect 267608 477204 267614 477216
rect 371050 477204 371056 477216
rect 267608 477176 371056 477204
rect 267608 477164 267614 477176
rect 371050 477164 371056 477176
rect 371108 477164 371114 477216
rect 255682 477096 255688 477148
rect 255740 477136 255746 477148
rect 361022 477136 361028 477148
rect 255740 477108 361028 477136
rect 255740 477096 255746 477108
rect 361022 477096 361028 477108
rect 361080 477096 361086 477148
rect 269758 477028 269764 477080
rect 269816 477068 269822 477080
rect 377950 477068 377956 477080
rect 269816 477040 377956 477068
rect 269816 477028 269822 477040
rect 377950 477028 377956 477040
rect 378008 477028 378014 477080
rect 167638 476960 167644 477012
rect 167696 477000 167702 477012
rect 214558 477000 214564 477012
rect 167696 476972 214564 477000
rect 167696 476960 167702 476972
rect 214558 476960 214564 476972
rect 214616 476960 214622 477012
rect 260558 476960 260564 477012
rect 260616 477000 260622 477012
rect 369486 477000 369492 477012
rect 260616 476972 369492 477000
rect 260616 476960 260622 476972
rect 369486 476960 369492 476972
rect 369544 476960 369550 477012
rect 163222 476892 163228 476944
rect 163280 476932 163286 476944
rect 210234 476932 210240 476944
rect 163280 476904 210240 476932
rect 163280 476892 163286 476904
rect 210234 476892 210240 476904
rect 210292 476892 210298 476944
rect 256602 476892 256608 476944
rect 256660 476932 256666 476944
rect 368106 476932 368112 476944
rect 256660 476904 368112 476932
rect 256660 476892 256666 476904
rect 368106 476892 368112 476904
rect 368164 476892 368170 476944
rect 60550 476824 60556 476876
rect 60608 476864 60614 476876
rect 133138 476864 133144 476876
rect 60608 476836 133144 476864
rect 60608 476824 60614 476836
rect 133138 476824 133144 476836
rect 133196 476824 133202 476876
rect 164050 476824 164056 476876
rect 164108 476864 164114 476876
rect 214650 476864 214656 476876
rect 164108 476836 214656 476864
rect 164108 476824 164114 476836
rect 214650 476824 214656 476836
rect 214708 476824 214714 476876
rect 242894 476824 242900 476876
rect 242952 476864 242958 476876
rect 363782 476864 363788 476876
rect 242952 476836 363788 476864
rect 242952 476824 242958 476836
rect 363782 476824 363788 476836
rect 363840 476824 363846 476876
rect 14458 476756 14464 476808
rect 14516 476796 14522 476808
rect 378134 476796 378140 476808
rect 14516 476768 378140 476796
rect 14516 476756 14522 476768
rect 378134 476756 378140 476768
rect 378192 476756 378198 476808
rect 70394 476076 70400 476128
rect 70452 476116 70458 476128
rect 70854 476116 70860 476128
rect 70452 476088 70860 476116
rect 70452 476076 70458 476088
rect 70854 476076 70860 476088
rect 70912 476076 70918 476128
rect 85574 476076 85580 476128
rect 85632 476116 85638 476128
rect 85758 476116 85764 476128
rect 85632 476088 85764 476116
rect 85632 476076 85638 476088
rect 85758 476076 85764 476088
rect 85816 476076 85822 476128
rect 51902 476008 51908 476060
rect 51960 476048 51966 476060
rect 98454 476048 98460 476060
rect 51960 476020 98460 476048
rect 51960 476008 51966 476020
rect 98454 476008 98460 476020
rect 98512 476008 98518 476060
rect 183526 476020 193214 476048
rect 48038 475940 48044 475992
rect 48096 475980 48102 475992
rect 97166 475980 97172 475992
rect 48096 475952 97172 475980
rect 48096 475940 48102 475952
rect 97166 475940 97172 475952
rect 97224 475940 97230 475992
rect 178126 475940 178132 475992
rect 178184 475980 178190 475992
rect 183526 475980 183554 476020
rect 178184 475952 183554 475980
rect 193186 475980 193214 476020
rect 203518 475980 203524 475992
rect 193186 475952 203524 475980
rect 178184 475940 178190 475952
rect 203518 475940 203524 475952
rect 203576 475940 203582 475992
rect 49050 475872 49056 475924
rect 49108 475912 49114 475924
rect 97994 475912 98000 475924
rect 49108 475884 98000 475912
rect 49108 475872 49114 475884
rect 97994 475872 98000 475884
rect 98052 475872 98058 475924
rect 186498 475872 186504 475924
rect 186556 475912 186562 475924
rect 212074 475912 212080 475924
rect 186556 475884 212080 475912
rect 186556 475872 186562 475884
rect 212074 475872 212080 475884
rect 212132 475872 212138 475924
rect 283834 475872 283840 475924
rect 283892 475912 283898 475924
rect 359918 475912 359924 475924
rect 283892 475884 359924 475912
rect 283892 475872 283898 475884
rect 359918 475872 359924 475884
rect 359976 475872 359982 475924
rect 59814 475804 59820 475856
rect 59872 475844 59878 475856
rect 119614 475844 119620 475856
rect 59872 475816 119620 475844
rect 59872 475804 59878 475816
rect 119614 475804 119620 475816
rect 119672 475804 119678 475856
rect 165430 475804 165436 475856
rect 165488 475844 165494 475856
rect 211798 475844 211804 475856
rect 165488 475816 211804 475844
rect 165488 475804 165494 475816
rect 211798 475804 211804 475816
rect 211856 475804 211862 475856
rect 294874 475804 294880 475856
rect 294932 475844 294938 475856
rect 379146 475844 379152 475856
rect 294932 475816 379152 475844
rect 294932 475804 294938 475816
rect 379146 475804 379152 475816
rect 379204 475804 379210 475856
rect 48130 475736 48136 475788
rect 48188 475776 48194 475788
rect 111702 475776 111708 475788
rect 48188 475748 111708 475776
rect 48188 475736 48194 475748
rect 111702 475736 111708 475748
rect 111760 475736 111766 475788
rect 160094 475736 160100 475788
rect 160152 475776 160158 475788
rect 210418 475776 210424 475788
rect 160152 475748 210424 475776
rect 160152 475736 160158 475748
rect 210418 475736 210424 475748
rect 210476 475736 210482 475788
rect 272426 475736 272432 475788
rect 272484 475776 272490 475788
rect 367002 475776 367008 475788
rect 272484 475748 367008 475776
rect 272484 475736 272490 475748
rect 367002 475736 367008 475748
rect 367060 475736 367066 475788
rect 47854 475668 47860 475720
rect 47912 475708 47918 475720
rect 112070 475708 112076 475720
rect 47912 475680 112076 475708
rect 47912 475668 47918 475680
rect 112070 475668 112076 475680
rect 112128 475668 112134 475720
rect 137646 475668 137652 475720
rect 137704 475708 137710 475720
rect 198090 475708 198096 475720
rect 137704 475680 198096 475708
rect 137704 475668 137710 475680
rect 198090 475668 198096 475680
rect 198148 475668 198154 475720
rect 271506 475668 271512 475720
rect 271564 475708 271570 475720
rect 371786 475708 371792 475720
rect 271564 475680 371792 475708
rect 271564 475668 271570 475680
rect 371786 475668 371792 475680
rect 371844 475668 371850 475720
rect 46382 475600 46388 475652
rect 46440 475640 46446 475652
rect 111242 475640 111248 475652
rect 46440 475612 111248 475640
rect 46440 475600 46446 475612
rect 111242 475600 111248 475612
rect 111300 475600 111306 475652
rect 138566 475600 138572 475652
rect 138624 475640 138630 475652
rect 200390 475640 200396 475652
rect 138624 475612 200396 475640
rect 138624 475600 138630 475612
rect 200390 475600 200396 475612
rect 200448 475600 200454 475652
rect 270218 475600 270224 475652
rect 270276 475640 270282 475652
rect 376478 475640 376484 475652
rect 270276 475612 376484 475640
rect 270276 475600 270282 475612
rect 376478 475600 376484 475612
rect 376536 475600 376542 475652
rect 48958 475532 48964 475584
rect 49016 475572 49022 475584
rect 115198 475572 115204 475584
rect 49016 475544 115204 475572
rect 49016 475532 49022 475544
rect 115198 475532 115204 475544
rect 115256 475532 115262 475584
rect 138106 475532 138112 475584
rect 138164 475572 138170 475584
rect 200298 475572 200304 475584
rect 138164 475544 200304 475572
rect 138164 475532 138170 475544
rect 200298 475532 200304 475544
rect 200356 475532 200362 475584
rect 260926 475532 260932 475584
rect 260984 475572 260990 475584
rect 374914 475572 374920 475584
rect 260984 475544 374920 475572
rect 260984 475532 260990 475544
rect 374914 475532 374920 475544
rect 374972 475532 374978 475584
rect 46750 475464 46756 475516
rect 46808 475504 46814 475516
rect 115658 475504 115664 475516
rect 46808 475476 115664 475504
rect 46808 475464 46814 475476
rect 115658 475464 115664 475476
rect 115716 475464 115722 475516
rect 135898 475464 135904 475516
rect 135956 475504 135962 475516
rect 197814 475504 197820 475516
rect 135956 475476 197820 475504
rect 135956 475464 135962 475476
rect 197814 475464 197820 475476
rect 197872 475464 197878 475516
rect 209958 475464 209964 475516
rect 210016 475504 210022 475516
rect 210142 475504 210148 475516
rect 210016 475476 210148 475504
rect 210016 475464 210022 475476
rect 210142 475464 210148 475476
rect 210200 475464 210206 475516
rect 211246 475464 211252 475516
rect 211304 475464 211310 475516
rect 246390 475464 246396 475516
rect 246448 475504 246454 475516
rect 365162 475504 365168 475516
rect 246448 475476 365168 475504
rect 246448 475464 246454 475476
rect 365162 475464 365168 475476
rect 365220 475464 365226 475516
rect 49142 475396 49148 475448
rect 49200 475436 49206 475448
rect 120074 475436 120080 475448
rect 49200 475408 120080 475436
rect 49200 475396 49206 475408
rect 120074 475396 120080 475408
rect 120132 475396 120138 475448
rect 122834 475396 122840 475448
rect 122892 475436 122898 475448
rect 123662 475436 123668 475448
rect 122892 475408 123668 475436
rect 122892 475396 122898 475408
rect 123662 475396 123668 475408
rect 123720 475396 123726 475448
rect 136726 475396 136732 475448
rect 136784 475436 136790 475448
rect 199654 475436 199660 475448
rect 136784 475408 199660 475436
rect 136784 475396 136790 475408
rect 199654 475396 199660 475408
rect 199712 475396 199718 475448
rect 60734 475328 60740 475380
rect 60792 475368 60798 475380
rect 61102 475368 61108 475380
rect 60792 475340 61108 475368
rect 60792 475328 60798 475340
rect 61102 475328 61108 475340
rect 61160 475328 61166 475380
rect 62114 475328 62120 475380
rect 62172 475368 62178 475380
rect 62942 475368 62948 475380
rect 62172 475340 62948 475368
rect 62172 475328 62178 475340
rect 62942 475328 62948 475340
rect 63000 475328 63006 475380
rect 63034 475328 63040 475380
rect 63092 475368 63098 475380
rect 134978 475368 134984 475380
rect 63092 475340 134984 475368
rect 63092 475328 63098 475340
rect 134978 475328 134984 475340
rect 135036 475328 135042 475380
rect 139394 475328 139400 475380
rect 139452 475368 139458 475380
rect 140038 475368 140044 475380
rect 139452 475340 140044 475368
rect 139452 475328 139458 475340
rect 140038 475328 140044 475340
rect 140096 475328 140102 475380
rect 140866 475328 140872 475380
rect 140924 475368 140930 475380
rect 141694 475368 141700 475380
rect 140924 475340 141700 475368
rect 140924 475328 140930 475340
rect 141694 475328 141700 475340
rect 141752 475328 141758 475380
rect 142126 475340 180794 475368
rect 54754 475260 54760 475312
rect 54812 475300 54818 475312
rect 96706 475300 96712 475312
rect 54812 475272 96712 475300
rect 54812 475260 54818 475272
rect 96706 475260 96712 475272
rect 96764 475260 96770 475312
rect 100846 475260 100852 475312
rect 100904 475300 100910 475312
rect 101582 475300 101588 475312
rect 100904 475272 101588 475300
rect 100904 475260 100910 475272
rect 101582 475260 101588 475272
rect 101640 475260 101646 475312
rect 103606 475260 103612 475312
rect 103664 475300 103670 475312
rect 103790 475300 103796 475312
rect 103664 475272 103796 475300
rect 103664 475260 103670 475272
rect 103790 475260 103796 475272
rect 103848 475260 103854 475312
rect 104986 475260 104992 475312
rect 105044 475300 105050 475312
rect 105630 475300 105636 475312
rect 105044 475272 105636 475300
rect 105044 475260 105050 475272
rect 105630 475260 105636 475272
rect 105688 475260 105694 475312
rect 106366 475260 106372 475312
rect 106424 475300 106430 475312
rect 106550 475300 106556 475312
rect 106424 475272 106556 475300
rect 106424 475260 106430 475272
rect 106550 475260 106556 475272
rect 106608 475260 106614 475312
rect 113266 475260 113272 475312
rect 113324 475300 113330 475312
rect 113542 475300 113548 475312
rect 113324 475272 113548 475300
rect 113324 475260 113330 475272
rect 113542 475260 113548 475272
rect 113600 475260 113606 475312
rect 122926 475260 122932 475312
rect 122984 475300 122990 475312
rect 123294 475300 123300 475312
rect 122984 475272 123300 475300
rect 122984 475260 122990 475272
rect 123294 475260 123300 475272
rect 123352 475260 123358 475312
rect 124214 475260 124220 475312
rect 124272 475300 124278 475312
rect 124950 475300 124956 475312
rect 124272 475272 124956 475300
rect 124272 475260 124278 475272
rect 124950 475260 124956 475272
rect 125008 475260 125014 475312
rect 125594 475260 125600 475312
rect 125652 475300 125658 475312
rect 126330 475300 126336 475312
rect 125652 475272 126336 475300
rect 125652 475260 125658 475272
rect 126330 475260 126336 475272
rect 126388 475260 126394 475312
rect 140774 475260 140780 475312
rect 140832 475300 140838 475312
rect 141326 475300 141332 475312
rect 140832 475272 141332 475300
rect 140832 475260 140838 475272
rect 141326 475260 141332 475272
rect 141384 475260 141390 475312
rect 58802 475192 58808 475244
rect 58860 475232 58866 475244
rect 96246 475232 96252 475244
rect 58860 475204 96252 475232
rect 58860 475192 58866 475204
rect 96246 475192 96252 475204
rect 96304 475192 96310 475244
rect 103514 475192 103520 475244
rect 103572 475232 103578 475244
rect 104342 475232 104348 475244
rect 103572 475204 104348 475232
rect 103572 475192 103578 475204
rect 104342 475192 104348 475204
rect 104400 475192 104406 475244
rect 106274 475192 106280 475244
rect 106332 475232 106338 475244
rect 106918 475232 106924 475244
rect 106332 475204 106924 475232
rect 106332 475192 106338 475204
rect 106918 475192 106924 475204
rect 106976 475192 106982 475244
rect 135438 475192 135444 475244
rect 135496 475232 135502 475244
rect 142126 475232 142154 475340
rect 143626 475260 143632 475312
rect 143684 475300 143690 475312
rect 144454 475300 144460 475312
rect 143684 475272 144460 475300
rect 143684 475260 143690 475272
rect 144454 475260 144460 475272
rect 144512 475260 144518 475312
rect 146294 475260 146300 475312
rect 146352 475300 146358 475312
rect 146662 475300 146668 475312
rect 146352 475272 146668 475300
rect 146352 475260 146358 475272
rect 146662 475260 146668 475272
rect 146720 475260 146726 475312
rect 165614 475260 165620 475312
rect 165672 475300 165678 475312
rect 166350 475300 166356 475312
rect 165672 475272 166356 475300
rect 165672 475260 165678 475272
rect 166350 475260 166356 475272
rect 166408 475260 166414 475312
rect 168374 475260 168380 475312
rect 168432 475300 168438 475312
rect 169110 475300 169116 475312
rect 168432 475272 169116 475300
rect 168432 475260 168438 475272
rect 169110 475260 169116 475272
rect 169168 475260 169174 475312
rect 172514 475260 172520 475312
rect 172572 475300 172578 475312
rect 173526 475300 173532 475312
rect 172572 475272 173532 475300
rect 172572 475260 172578 475272
rect 173526 475260 173532 475272
rect 173584 475260 173590 475312
rect 173894 475260 173900 475312
rect 173952 475300 173958 475312
rect 174262 475300 174268 475312
rect 173952 475272 174268 475300
rect 173952 475260 173958 475272
rect 174262 475260 174268 475272
rect 174320 475260 174326 475312
rect 175274 475260 175280 475312
rect 175332 475300 175338 475312
rect 176102 475300 176108 475312
rect 175332 475272 176108 475300
rect 175332 475260 175338 475272
rect 176102 475260 176108 475272
rect 176160 475260 176166 475312
rect 135496 475204 142154 475232
rect 180766 475232 180794 475340
rect 205726 475328 205732 475380
rect 205784 475368 205790 475380
rect 206462 475368 206468 475380
rect 205784 475340 206468 475368
rect 205784 475328 205790 475340
rect 206462 475328 206468 475340
rect 206520 475328 206526 475380
rect 207198 475328 207204 475380
rect 207256 475368 207262 475380
rect 207750 475368 207756 475380
rect 207256 475340 207756 475368
rect 207256 475328 207262 475340
rect 207750 475328 207756 475340
rect 207808 475328 207814 475380
rect 209774 475328 209780 475380
rect 209832 475368 209838 475380
rect 210510 475368 210516 475380
rect 209832 475340 210516 475368
rect 209832 475328 209838 475340
rect 210510 475328 210516 475340
rect 210568 475328 210574 475380
rect 211264 475312 211292 475464
rect 238110 475396 238116 475448
rect 238168 475436 238174 475448
rect 362402 475436 362408 475448
rect 238168 475408 362408 475436
rect 238168 475396 238174 475408
rect 362402 475396 362408 475408
rect 362460 475396 362466 475448
rect 212718 475328 212724 475380
rect 212776 475368 212782 475380
rect 213086 475368 213092 475380
rect 212776 475340 213092 475368
rect 212776 475328 212782 475340
rect 213086 475328 213092 475340
rect 213144 475328 213150 475380
rect 213914 475328 213920 475380
rect 213972 475368 213978 475380
rect 214926 475368 214932 475380
rect 213972 475340 214932 475368
rect 213972 475328 213978 475340
rect 214926 475328 214932 475340
rect 214984 475328 214990 475380
rect 215386 475328 215392 475380
rect 215444 475368 215450 475380
rect 216214 475368 216220 475380
rect 215444 475340 216220 475368
rect 215444 475328 215450 475340
rect 216214 475328 216220 475340
rect 216272 475328 216278 475380
rect 218054 475328 218060 475380
rect 218112 475368 218118 475380
rect 218790 475368 218796 475380
rect 218112 475340 218796 475368
rect 218112 475328 218118 475340
rect 218790 475328 218796 475340
rect 218848 475328 218854 475380
rect 219434 475328 219440 475380
rect 219492 475368 219498 475380
rect 220078 475368 220084 475380
rect 219492 475340 220084 475368
rect 219492 475328 219498 475340
rect 220078 475328 220084 475340
rect 220136 475328 220142 475380
rect 223574 475328 223580 475380
rect 223632 475368 223638 475380
rect 224494 475368 224500 475380
rect 223632 475340 224500 475368
rect 223632 475328 223638 475340
rect 224494 475328 224500 475340
rect 224552 475328 224558 475380
rect 226334 475328 226340 475380
rect 226392 475368 226398 475380
rect 226702 475368 226708 475380
rect 226392 475340 226708 475368
rect 226392 475328 226398 475340
rect 226702 475328 226708 475340
rect 226760 475328 226766 475380
rect 227714 475328 227720 475380
rect 227772 475368 227778 475380
rect 228542 475368 228548 475380
rect 227772 475340 228548 475368
rect 227772 475328 227778 475340
rect 228542 475328 228548 475340
rect 228600 475328 228606 475380
rect 229094 475328 229100 475380
rect 229152 475368 229158 475380
rect 229462 475368 229468 475380
rect 229152 475340 229468 475368
rect 229152 475328 229158 475340
rect 229462 475328 229468 475340
rect 229520 475328 229526 475380
rect 240134 475328 240140 475380
rect 240192 475368 240198 475380
rect 240870 475368 240876 475380
rect 240192 475340 240876 475368
rect 240192 475328 240198 475340
rect 240870 475328 240876 475340
rect 240928 475328 240934 475380
rect 244274 475328 244280 475380
rect 244332 475368 244338 475380
rect 244734 475368 244740 475380
rect 244332 475340 244740 475368
rect 244332 475328 244338 475340
rect 244734 475328 244740 475340
rect 244792 475328 244798 475380
rect 247126 475328 247132 475380
rect 247184 475368 247190 475380
rect 247494 475368 247500 475380
rect 247184 475340 247500 475368
rect 247184 475328 247190 475340
rect 247494 475328 247500 475340
rect 247552 475328 247558 475380
rect 369118 475368 369124 475380
rect 248386 475340 369124 475368
rect 203702 475260 203708 475312
rect 203760 475300 203766 475312
rect 209498 475300 209504 475312
rect 203760 475272 209504 475300
rect 203760 475260 203766 475272
rect 209498 475260 209504 475272
rect 209556 475260 209562 475312
rect 211246 475260 211252 475312
rect 211304 475260 211310 475312
rect 212534 475260 212540 475312
rect 212592 475300 212598 475312
rect 213454 475300 213460 475312
rect 212592 475272 213460 475300
rect 212592 475260 212598 475272
rect 213454 475260 213460 475272
rect 213512 475260 213518 475312
rect 215294 475260 215300 475312
rect 215352 475300 215358 475312
rect 215662 475300 215668 475312
rect 215352 475272 215668 475300
rect 215352 475260 215358 475272
rect 215662 475260 215668 475272
rect 215720 475260 215726 475312
rect 244366 475260 244372 475312
rect 244424 475300 244430 475312
rect 244550 475300 244556 475312
rect 244424 475272 244556 475300
rect 244424 475260 244430 475272
rect 244550 475260 244556 475272
rect 244608 475260 244614 475312
rect 247034 475260 247040 475312
rect 247092 475300 247098 475312
rect 247862 475300 247868 475312
rect 247092 475272 247868 475300
rect 247092 475260 247098 475272
rect 247862 475260 247868 475272
rect 247920 475260 247926 475312
rect 198182 475232 198188 475244
rect 180766 475204 198188 475232
rect 135496 475192 135502 475204
rect 198182 475192 198188 475204
rect 198240 475192 198246 475244
rect 210326 475192 210332 475244
rect 210384 475192 210390 475244
rect 220814 475192 220820 475244
rect 220872 475232 220878 475244
rect 220998 475232 221004 475244
rect 220872 475204 221004 475232
rect 220872 475192 220878 475204
rect 220998 475192 221004 475204
rect 221056 475192 221062 475244
rect 242066 475192 242072 475244
rect 242124 475232 242130 475244
rect 248386 475232 248414 475340
rect 369118 475328 369124 475340
rect 369176 475328 369182 475380
rect 248506 475260 248512 475312
rect 248564 475300 248570 475312
rect 249150 475300 249156 475312
rect 248564 475272 249156 475300
rect 248564 475260 248570 475272
rect 249150 475260 249156 475272
rect 249208 475260 249214 475312
rect 262214 475260 262220 475312
rect 262272 475300 262278 475312
rect 262398 475300 262404 475312
rect 262272 475272 262404 475300
rect 262272 475260 262278 475272
rect 262398 475260 262404 475272
rect 262456 475260 262462 475312
rect 263594 475260 263600 475312
rect 263652 475300 263658 475312
rect 264238 475300 264244 475312
rect 263652 475272 264244 475300
rect 263652 475260 263658 475272
rect 264238 475260 264244 475272
rect 264296 475260 264302 475312
rect 264974 475260 264980 475312
rect 265032 475300 265038 475312
rect 265894 475300 265900 475312
rect 265032 475272 265900 475300
rect 265032 475260 265038 475272
rect 265894 475260 265900 475272
rect 265952 475260 265958 475312
rect 292574 475260 292580 475312
rect 292632 475300 292638 475312
rect 293310 475300 293316 475312
rect 292632 475272 293316 475300
rect 292632 475260 292638 475272
rect 293310 475260 293316 475272
rect 293368 475260 293374 475312
rect 296714 475260 296720 475312
rect 296772 475300 296778 475312
rect 297726 475300 297732 475312
rect 296772 475272 297732 475300
rect 296772 475260 296778 475272
rect 297726 475260 297732 475272
rect 297784 475260 297790 475312
rect 242124 475204 248414 475232
rect 242124 475192 242130 475204
rect 59722 475124 59728 475176
rect 59780 475164 59786 475176
rect 97534 475164 97540 475176
rect 59780 475136 97540 475164
rect 59780 475124 59786 475136
rect 97534 475124 97540 475136
rect 97592 475124 97598 475176
rect 142154 475124 142160 475176
rect 142212 475164 142218 475176
rect 142614 475164 142620 475176
rect 142212 475136 142620 475164
rect 142212 475124 142218 475136
rect 142614 475124 142620 475136
rect 142672 475124 142678 475176
rect 57330 475056 57336 475108
rect 57388 475096 57394 475108
rect 63034 475096 63040 475108
rect 57388 475068 63040 475096
rect 57388 475056 57394 475068
rect 63034 475056 63040 475068
rect 63092 475056 63098 475108
rect 66254 475056 66260 475108
rect 66312 475096 66318 475108
rect 66806 475096 66812 475108
rect 66312 475068 66812 475096
rect 66312 475056 66318 475068
rect 66806 475056 66812 475068
rect 66864 475056 66870 475108
rect 67818 475056 67824 475108
rect 67876 475096 67882 475108
rect 68646 475096 68652 475108
rect 67876 475068 68652 475096
rect 67876 475056 67882 475068
rect 68646 475056 68652 475068
rect 68704 475056 68710 475108
rect 71774 475056 71780 475108
rect 71832 475096 71838 475108
rect 72602 475096 72608 475108
rect 71832 475068 72608 475096
rect 71832 475056 71838 475068
rect 72602 475056 72608 475068
rect 72660 475056 72666 475108
rect 74534 475056 74540 475108
rect 74592 475096 74598 475108
rect 75270 475096 75276 475108
rect 74592 475068 75276 475096
rect 74592 475056 74598 475068
rect 75270 475056 75276 475068
rect 75328 475056 75334 475108
rect 78766 475056 78772 475108
rect 78824 475096 78830 475108
rect 79686 475096 79692 475108
rect 78824 475068 79692 475096
rect 78824 475056 78830 475068
rect 79686 475056 79692 475068
rect 79744 475056 79750 475108
rect 92566 475056 92572 475108
rect 92624 475096 92630 475108
rect 93302 475096 93308 475108
rect 92624 475068 93308 475096
rect 92624 475056 92630 475068
rect 93302 475056 93308 475068
rect 93360 475056 93366 475108
rect 210344 475040 210372 475192
rect 67634 474988 67640 475040
rect 67692 475028 67698 475040
rect 67910 475028 67916 475040
rect 67692 475000 67916 475028
rect 67692 474988 67698 475000
rect 67910 474988 67916 475000
rect 67968 474988 67974 475040
rect 210326 474988 210332 475040
rect 210384 474988 210390 475040
rect 297082 474580 297088 474632
rect 297140 474620 297146 474632
rect 362770 474620 362776 474632
rect 297140 474592 362776 474620
rect 297140 474580 297146 474592
rect 362770 474580 362776 474592
rect 362828 474580 362834 474632
rect 282546 474512 282552 474564
rect 282604 474552 282610 474564
rect 375098 474552 375104 474564
rect 282604 474524 375104 474552
rect 282604 474512 282610 474524
rect 375098 474512 375104 474524
rect 375156 474512 375162 474564
rect 272886 474444 272892 474496
rect 272944 474484 272950 474496
rect 369670 474484 369676 474496
rect 272944 474456 369676 474484
rect 272944 474444 272950 474456
rect 369670 474444 369676 474456
rect 369728 474444 369734 474496
rect 282086 474376 282092 474428
rect 282144 474416 282150 474428
rect 379974 474416 379980 474428
rect 282144 474388 379980 474416
rect 282144 474376 282150 474388
rect 379974 474376 379980 474388
rect 380032 474376 380038 474428
rect 265250 474308 265256 474360
rect 265308 474348 265314 474360
rect 369578 474348 369584 474360
rect 265308 474320 369584 474348
rect 265308 474308 265314 474320
rect 369578 474308 369584 474320
rect 369636 474308 369642 474360
rect 254394 474240 254400 474292
rect 254452 474280 254458 474292
rect 358446 474280 358452 474292
rect 254452 474252 358452 474280
rect 254452 474240 254458 474252
rect 358446 474240 358452 474252
rect 358504 474240 358510 474292
rect 265342 474172 265348 474224
rect 265400 474212 265406 474224
rect 372154 474212 372160 474224
rect 265400 474184 372160 474212
rect 265400 474172 265406 474184
rect 372154 474172 372160 474184
rect 372212 474172 372218 474224
rect 205910 474104 205916 474156
rect 205968 474144 205974 474156
rect 217318 474144 217324 474156
rect 205968 474116 217324 474144
rect 205968 474104 205974 474116
rect 217318 474104 217324 474116
rect 217376 474104 217382 474156
rect 260098 474104 260104 474156
rect 260156 474144 260162 474156
rect 368198 474144 368204 474156
rect 260156 474116 368204 474144
rect 260156 474104 260162 474116
rect 368198 474104 368204 474116
rect 368256 474104 368262 474156
rect 176010 474036 176016 474088
rect 176068 474076 176074 474088
rect 206554 474076 206560 474088
rect 176068 474048 206560 474076
rect 176068 474036 176074 474048
rect 206554 474036 206560 474048
rect 206612 474036 206618 474088
rect 246022 474036 246028 474088
rect 246080 474076 246086 474088
rect 369210 474076 369216 474088
rect 246080 474048 369216 474076
rect 246080 474036 246086 474048
rect 369210 474036 369216 474048
rect 369268 474036 369274 474088
rect 57882 473968 57888 474020
rect 57940 474008 57946 474020
rect 114278 474008 114284 474020
rect 57940 473980 114284 474008
rect 57940 473968 57946 473980
rect 114278 473968 114284 473980
rect 114336 473968 114342 474020
rect 159634 473968 159640 474020
rect 159692 474008 159698 474020
rect 216030 474008 216036 474020
rect 159692 473980 216036 474008
rect 159692 473968 159698 473980
rect 216030 473968 216036 473980
rect 216088 473968 216094 474020
rect 237190 473968 237196 474020
rect 237248 474008 237254 474020
rect 366726 474008 366732 474020
rect 237248 473980 366732 474008
rect 237248 473968 237254 473980
rect 366726 473968 366732 473980
rect 366784 473968 366790 474020
rect 48222 473288 48228 473340
rect 48280 473328 48286 473340
rect 117866 473328 117872 473340
rect 48280 473300 117872 473328
rect 48280 473288 48286 473300
rect 117866 473288 117872 473300
rect 117924 473288 117930 473340
rect 46566 473220 46572 473272
rect 46624 473260 46630 473272
rect 116486 473260 116492 473272
rect 46624 473232 116492 473260
rect 46624 473220 46630 473232
rect 116486 473220 116492 473232
rect 116544 473220 116550 473272
rect 49234 473152 49240 473204
rect 49292 473192 49298 473204
rect 119154 473192 119160 473204
rect 49292 473164 119160 473192
rect 49292 473152 49298 473164
rect 119154 473152 119160 473164
rect 119212 473152 119218 473204
rect 284754 473152 284760 473204
rect 284812 473192 284818 473204
rect 360010 473192 360016 473204
rect 284812 473164 360016 473192
rect 284812 473152 284818 473164
rect 360010 473152 360016 473164
rect 360068 473152 360074 473204
rect 45462 473084 45468 473136
rect 45520 473124 45526 473136
rect 118234 473124 118240 473136
rect 45520 473096 118240 473124
rect 45520 473084 45526 473096
rect 118234 473084 118240 473096
rect 118292 473084 118298 473136
rect 295978 473084 295984 473136
rect 296036 473124 296042 473136
rect 372614 473124 372620 473136
rect 296036 473096 372620 473124
rect 296036 473084 296042 473096
rect 372614 473084 372620 473096
rect 372672 473084 372678 473136
rect 53558 473016 53564 473068
rect 53616 473056 53622 473068
rect 131942 473056 131948 473068
rect 53616 473028 131948 473056
rect 53616 473016 53622 473028
rect 131942 473016 131948 473028
rect 132000 473016 132006 473068
rect 274174 473016 274180 473068
rect 274232 473056 274238 473068
rect 362862 473056 362868 473068
rect 274232 473028 362868 473056
rect 274232 473016 274238 473028
rect 362862 473016 362868 473028
rect 362920 473016 362926 473068
rect 57054 472948 57060 473000
rect 57112 472988 57118 473000
rect 136358 472988 136364 473000
rect 57112 472960 136364 472988
rect 57112 472948 57118 472960
rect 136358 472948 136364 472960
rect 136416 472948 136422 473000
rect 192110 472948 192116 473000
rect 192168 472988 192174 473000
rect 192662 472988 192668 473000
rect 192168 472960 192668 472988
rect 192168 472948 192174 472960
rect 192662 472948 192668 472960
rect 192720 472948 192726 473000
rect 261846 472948 261852 473000
rect 261904 472988 261910 473000
rect 372246 472988 372252 473000
rect 261904 472960 372252 472988
rect 261904 472948 261910 472960
rect 372246 472948 372252 472960
rect 372304 472948 372310 473000
rect 50154 472880 50160 472932
rect 50212 472920 50218 472932
rect 131482 472920 131488 472932
rect 50212 472892 131488 472920
rect 50212 472880 50218 472892
rect 131482 472880 131488 472892
rect 131540 472880 131546 472932
rect 182266 472880 182272 472932
rect 182324 472920 182330 472932
rect 183094 472920 183100 472932
rect 182324 472892 183100 472920
rect 182324 472880 182330 472892
rect 183094 472880 183100 472892
rect 183152 472880 183158 472932
rect 242434 472880 242440 472932
rect 242492 472920 242498 472932
rect 360930 472920 360936 472932
rect 242492 472892 360936 472920
rect 242492 472880 242498 472892
rect 360930 472880 360936 472892
rect 360988 472880 360994 472932
rect 48866 472812 48872 472864
rect 48924 472852 48930 472864
rect 129734 472852 129740 472864
rect 48924 472824 129740 472852
rect 48924 472812 48930 472824
rect 129734 472812 129740 472824
rect 129792 472812 129798 472864
rect 245562 472812 245568 472864
rect 245620 472852 245626 472864
rect 370682 472852 370688 472864
rect 245620 472824 370688 472852
rect 245620 472812 245626 472824
rect 370682 472812 370688 472824
rect 370740 472812 370746 472864
rect 47762 472744 47768 472796
rect 47820 472784 47826 472796
rect 131022 472784 131028 472796
rect 47820 472756 131028 472784
rect 47820 472744 47826 472756
rect 131022 472744 131028 472756
rect 131080 472744 131086 472796
rect 234982 472744 234988 472796
rect 235040 472784 235046 472796
rect 364978 472784 364984 472796
rect 235040 472756 364984 472784
rect 235040 472744 235046 472756
rect 364978 472744 364984 472756
rect 365036 472744 365042 472796
rect 46290 472676 46296 472728
rect 46348 472716 46354 472728
rect 130562 472716 130568 472728
rect 46348 472688 130568 472716
rect 46348 472676 46354 472688
rect 130562 472676 130568 472688
rect 130620 472676 130626 472728
rect 172422 472676 172428 472728
rect 172480 472716 172486 472728
rect 210602 472716 210608 472728
rect 172480 472688 210608 472716
rect 172480 472676 172486 472688
rect 210602 472676 210608 472688
rect 210660 472676 210666 472728
rect 238938 472676 238944 472728
rect 238996 472716 239002 472728
rect 378778 472716 378784 472728
rect 238996 472688 378784 472716
rect 238996 472676 239002 472688
rect 378778 472676 378784 472688
rect 378836 472676 378842 472728
rect 46106 472608 46112 472660
rect 46164 472648 46170 472660
rect 143810 472648 143816 472660
rect 46164 472620 143816 472648
rect 46164 472608 46170 472620
rect 143810 472608 143816 472620
rect 143868 472608 143874 472660
rect 147766 472608 147772 472660
rect 147824 472648 147830 472660
rect 218698 472648 218704 472660
rect 147824 472620 218704 472648
rect 147824 472608 147830 472620
rect 218698 472608 218704 472620
rect 218756 472608 218762 472660
rect 227530 472608 227536 472660
rect 227588 472648 227594 472660
rect 371878 472648 371884 472660
rect 227588 472620 371884 472648
rect 227588 472608 227594 472620
rect 371878 472608 371884 472620
rect 371936 472608 371942 472660
rect 46658 472540 46664 472592
rect 46716 472580 46722 472592
rect 116946 472580 116952 472592
rect 46716 472552 116952 472580
rect 46716 472540 46722 472552
rect 116946 472540 116952 472552
rect 117004 472540 117010 472592
rect 50430 472472 50436 472524
rect 50488 472512 50494 472524
rect 116026 472512 116032 472524
rect 50488 472484 116032 472512
rect 50488 472472 50494 472484
rect 116026 472472 116032 472484
rect 116084 472472 116090 472524
rect 58618 472404 58624 472456
rect 58676 472444 58682 472456
rect 118694 472444 118700 472456
rect 58676 472416 118700 472444
rect 58676 472404 58682 472416
rect 118694 472404 118700 472416
rect 118752 472404 118758 472456
rect 258074 472064 258080 472116
rect 258132 472104 258138 472116
rect 258902 472104 258908 472116
rect 258132 472076 258908 472104
rect 258132 472064 258138 472076
rect 258902 472064 258908 472076
rect 258960 472064 258966 472116
rect 280246 471928 280252 471980
rect 280304 471968 280310 471980
rect 280430 471968 280436 471980
rect 280304 471940 280436 471968
rect 280304 471928 280310 471940
rect 280430 471928 280436 471940
rect 280488 471928 280494 471980
rect 292206 471928 292212 471980
rect 292264 471968 292270 471980
rect 368290 471968 368296 471980
rect 292264 471940 368296 471968
rect 292264 471928 292270 471940
rect 368290 471928 368296 471940
rect 368348 471928 368354 471980
rect 269298 471860 269304 471912
rect 269356 471900 269362 471912
rect 356882 471900 356888 471912
rect 269356 471872 356888 471900
rect 269356 471860 269362 471872
rect 356882 471860 356888 471872
rect 356940 471860 356946 471912
rect 263778 471792 263784 471844
rect 263836 471832 263842 471844
rect 365346 471832 365352 471844
rect 263836 471804 365352 471832
rect 263836 471792 263842 471804
rect 365346 471792 365352 471804
rect 365404 471792 365410 471844
rect 258350 471724 258356 471776
rect 258408 471764 258414 471776
rect 362586 471764 362592 471776
rect 258408 471736 362592 471764
rect 258408 471724 258414 471736
rect 362586 471724 362592 471736
rect 362644 471724 362650 471776
rect 273714 471656 273720 471708
rect 273772 471696 273778 471708
rect 378042 471696 378048 471708
rect 273772 471668 378048 471696
rect 273772 471656 273778 471668
rect 378042 471656 378048 471668
rect 378100 471656 378106 471708
rect 270678 471588 270684 471640
rect 270736 471628 270742 471640
rect 377674 471628 377680 471640
rect 270736 471600 377680 471628
rect 270736 471588 270742 471600
rect 377674 471588 377680 471600
rect 377732 471588 377738 471640
rect 252186 471520 252192 471572
rect 252244 471560 252250 471572
rect 361206 471560 361212 471572
rect 252244 471532 361212 471560
rect 252244 471520 252250 471532
rect 361206 471520 361212 471532
rect 361264 471520 361270 471572
rect 198918 471452 198924 471504
rect 198976 471492 198982 471504
rect 199102 471492 199108 471504
rect 198976 471464 199108 471492
rect 198976 471452 198982 471464
rect 199102 471452 199108 471464
rect 199160 471452 199166 471504
rect 263134 471452 263140 471504
rect 263192 471492 263198 471504
rect 375006 471492 375012 471504
rect 263192 471464 375012 471492
rect 263192 471452 263198 471464
rect 375006 471452 375012 471464
rect 375064 471452 375070 471504
rect 180334 471384 180340 471436
rect 180392 471424 180398 471436
rect 209222 471424 209228 471436
rect 180392 471396 209228 471424
rect 180392 471384 180398 471396
rect 209222 471384 209228 471396
rect 209280 471384 209286 471436
rect 237650 471384 237656 471436
rect 237708 471424 237714 471436
rect 367738 471424 367744 471436
rect 237708 471396 367744 471424
rect 237708 471384 237714 471396
rect 367738 471384 367744 471396
rect 367796 471384 367802 471436
rect 57238 471316 57244 471368
rect 57296 471356 57302 471368
rect 129274 471356 129280 471368
rect 57296 471328 129280 471356
rect 57296 471316 57302 471328
rect 129274 471316 129280 471328
rect 129332 471316 129338 471368
rect 162026 471316 162032 471368
rect 162084 471356 162090 471368
rect 211890 471356 211896 471368
rect 162084 471328 211896 471356
rect 162084 471316 162090 471328
rect 211890 471316 211896 471328
rect 211948 471316 211954 471368
rect 246850 471316 246856 471368
rect 246908 471356 246914 471368
rect 378870 471356 378876 471368
rect 246908 471328 378876 471356
rect 246908 471316 246914 471328
rect 378870 471316 378876 471328
rect 378928 471316 378934 471368
rect 61930 471248 61936 471300
rect 61988 471288 61994 471300
rect 61988 471260 195974 471288
rect 61988 471248 61994 471260
rect 81526 471180 81532 471232
rect 81584 471220 81590 471232
rect 82262 471220 82268 471232
rect 81584 471192 82268 471220
rect 81584 471180 81590 471192
rect 82262 471180 82268 471192
rect 82320 471180 82326 471232
rect 82814 471180 82820 471232
rect 82872 471220 82878 471232
rect 82998 471220 83004 471232
rect 82872 471192 83004 471220
rect 82872 471180 82878 471192
rect 82998 471180 83004 471192
rect 83056 471180 83062 471232
rect 85666 471180 85672 471232
rect 85724 471220 85730 471232
rect 86310 471220 86316 471232
rect 85724 471192 86316 471220
rect 85724 471180 85730 471192
rect 86310 471180 86316 471192
rect 86368 471180 86374 471232
rect 189166 471180 189172 471232
rect 189224 471220 189230 471232
rect 189718 471220 189724 471232
rect 189224 471192 189724 471220
rect 189224 471180 189230 471192
rect 189718 471180 189724 471192
rect 189776 471180 189782 471232
rect 192018 471180 192024 471232
rect 192076 471220 192082 471232
rect 192846 471220 192852 471232
rect 192076 471192 192852 471220
rect 192076 471180 192082 471192
rect 192846 471180 192852 471192
rect 192904 471180 192910 471232
rect 193214 471180 193220 471232
rect 193272 471220 193278 471232
rect 193766 471220 193772 471232
rect 193272 471192 193772 471220
rect 193272 471180 193278 471192
rect 193766 471180 193772 471192
rect 193824 471180 193830 471232
rect 195946 471220 195974 471260
rect 196710 471248 196716 471300
rect 196768 471288 196774 471300
rect 196894 471288 196900 471300
rect 196768 471260 196900 471288
rect 196768 471248 196774 471260
rect 196894 471248 196900 471260
rect 196952 471248 196958 471300
rect 197354 471248 197360 471300
rect 197412 471288 197418 471300
rect 197630 471288 197636 471300
rect 197412 471260 197636 471288
rect 197412 471248 197418 471260
rect 197630 471248 197636 471260
rect 197688 471248 197694 471300
rect 198734 471248 198740 471300
rect 198792 471288 198798 471300
rect 199470 471288 199476 471300
rect 198792 471260 199476 471288
rect 198792 471248 198798 471260
rect 199470 471248 199476 471260
rect 199528 471248 199534 471300
rect 201494 471248 201500 471300
rect 201552 471288 201558 471300
rect 201678 471288 201684 471300
rect 201552 471260 201684 471288
rect 201552 471248 201558 471260
rect 201678 471248 201684 471260
rect 201736 471248 201742 471300
rect 203058 471248 203064 471300
rect 203116 471288 203122 471300
rect 203886 471288 203892 471300
rect 203116 471260 203892 471288
rect 203116 471248 203122 471260
rect 203886 471248 203892 471260
rect 203944 471248 203950 471300
rect 204346 471248 204352 471300
rect 204404 471288 204410 471300
rect 205174 471288 205180 471300
rect 204404 471260 205180 471288
rect 204404 471248 204410 471260
rect 205174 471248 205180 471260
rect 205232 471248 205238 471300
rect 217686 471288 217692 471300
rect 205606 471260 217692 471288
rect 199194 471220 199200 471232
rect 195946 471192 199200 471220
rect 199194 471180 199200 471192
rect 199252 471180 199258 471232
rect 202874 471180 202880 471232
rect 202932 471220 202938 471232
rect 203150 471220 203156 471232
rect 202932 471192 203156 471220
rect 202932 471180 202938 471192
rect 203150 471180 203156 471192
rect 203208 471180 203214 471232
rect 204990 471180 204996 471232
rect 205048 471220 205054 471232
rect 205606 471220 205634 471260
rect 217686 471248 217692 471260
rect 217744 471248 217750 471300
rect 227898 471248 227904 471300
rect 227956 471288 227962 471300
rect 362310 471288 362316 471300
rect 227956 471260 362316 471288
rect 227956 471248 227962 471260
rect 362310 471248 362316 471260
rect 362368 471248 362374 471300
rect 205048 471192 205634 471220
rect 205048 471180 205054 471192
rect 277394 471180 277400 471232
rect 277452 471220 277458 471232
rect 277854 471220 277860 471232
rect 277452 471192 277860 471220
rect 277452 471180 277458 471192
rect 277854 471180 277860 471192
rect 277912 471180 277918 471232
rect 278774 471180 278780 471232
rect 278832 471220 278838 471232
rect 279142 471220 279148 471232
rect 278832 471192 279148 471220
rect 278832 471180 278838 471192
rect 279142 471180 279148 471192
rect 279200 471180 279206 471232
rect 287054 471180 287060 471232
rect 287112 471220 287118 471232
rect 287974 471220 287980 471232
rect 287112 471192 287980 471220
rect 287112 471180 287118 471192
rect 287974 471180 287980 471192
rect 288032 471180 288038 471232
rect 361298 471220 361304 471232
rect 292546 471192 361304 471220
rect 191834 471112 191840 471164
rect 191892 471152 191898 471164
rect 192386 471152 192392 471164
rect 191892 471124 192392 471152
rect 191892 471112 191898 471124
rect 192386 471112 192392 471124
rect 192444 471112 192450 471164
rect 193306 471112 193312 471164
rect 193364 471152 193370 471164
rect 194134 471152 194140 471164
rect 193364 471124 194140 471152
rect 193364 471112 193370 471124
rect 194134 471112 194140 471124
rect 194192 471112 194198 471164
rect 287422 471112 287428 471164
rect 287480 471152 287486 471164
rect 292546 471152 292574 471192
rect 361298 471180 361304 471192
rect 361356 471180 361362 471232
rect 287480 471124 292574 471152
rect 287480 471112 287486 471124
rect 82814 471044 82820 471096
rect 82872 471084 82878 471096
rect 83550 471084 83556 471096
rect 82872 471056 83556 471084
rect 82872 471044 82878 471056
rect 83550 471044 83556 471056
rect 83608 471044 83614 471096
rect 55674 470500 55680 470552
rect 55732 470540 55738 470552
rect 128354 470540 128360 470552
rect 55732 470512 128360 470540
rect 55732 470500 55738 470512
rect 128354 470500 128360 470512
rect 128412 470500 128418 470552
rect 54386 470432 54392 470484
rect 54444 470472 54450 470484
rect 127066 470472 127072 470484
rect 54444 470444 127072 470472
rect 54444 470432 54450 470444
rect 127066 470432 127072 470444
rect 127124 470432 127130 470484
rect 57146 470364 57152 470416
rect 57204 470404 57210 470416
rect 132770 470404 132776 470416
rect 57204 470376 132776 470404
rect 57204 470364 57210 470376
rect 132770 470364 132776 470376
rect 132828 470364 132834 470416
rect 275186 470364 275192 470416
rect 275244 470404 275250 470416
rect 359458 470404 359464 470416
rect 275244 470376 359464 470404
rect 275244 470364 275250 470376
rect 359458 470364 359464 470376
rect 359516 470364 359522 470416
rect 43898 470296 43904 470348
rect 43956 470336 43962 470348
rect 122834 470336 122840 470348
rect 43956 470308 122840 470336
rect 43956 470296 43962 470308
rect 122834 470296 122840 470308
rect 122892 470296 122898 470348
rect 187694 470296 187700 470348
rect 187752 470336 187758 470348
rect 188430 470336 188436 470348
rect 187752 470308 188436 470336
rect 187752 470296 187758 470308
rect 188430 470296 188436 470308
rect 188488 470296 188494 470348
rect 274726 470296 274732 470348
rect 274784 470336 274790 470348
rect 364150 470336 364156 470348
rect 274784 470308 364156 470336
rect 274784 470296 274790 470308
rect 364150 470296 364156 470308
rect 364208 470296 364214 470348
rect 42426 470228 42432 470280
rect 42484 470268 42490 470280
rect 122926 470268 122932 470280
rect 42484 470240 122932 470268
rect 42484 470228 42490 470240
rect 122926 470228 122932 470240
rect 122984 470228 122990 470280
rect 286042 470228 286048 470280
rect 286100 470268 286106 470280
rect 376754 470268 376760 470280
rect 286100 470240 376760 470268
rect 286100 470228 286106 470240
rect 376754 470228 376760 470240
rect 376812 470228 376818 470280
rect 43714 470160 43720 470212
rect 43772 470200 43778 470212
rect 124398 470200 124404 470212
rect 43772 470172 124404 470200
rect 43772 470160 43778 470172
rect 124398 470160 124404 470172
rect 124456 470160 124462 470212
rect 265066 470160 265072 470212
rect 265124 470200 265130 470212
rect 362678 470200 362684 470212
rect 265124 470172 362684 470200
rect 265124 470160 265130 470172
rect 362678 470160 362684 470172
rect 362736 470160 362742 470212
rect 42334 470092 42340 470144
rect 42392 470132 42398 470144
rect 123018 470132 123024 470144
rect 42392 470104 123024 470132
rect 42392 470092 42398 470104
rect 123018 470092 123024 470104
rect 123076 470092 123082 470144
rect 256878 470092 256884 470144
rect 256936 470132 256942 470144
rect 366818 470132 366824 470144
rect 256936 470104 366824 470132
rect 256936 470092 256942 470104
rect 366818 470092 366824 470104
rect 366876 470092 366882 470144
rect 51534 470024 51540 470076
rect 51592 470064 51598 470076
rect 133966 470064 133972 470076
rect 51592 470036 133972 470064
rect 51592 470024 51598 470036
rect 133966 470024 133972 470036
rect 134024 470024 134030 470076
rect 244458 470024 244464 470076
rect 244516 470064 244522 470076
rect 371970 470064 371976 470076
rect 244516 470036 371976 470064
rect 244516 470024 244522 470036
rect 371970 470024 371976 470036
rect 372028 470024 372034 470076
rect 48774 469956 48780 470008
rect 48832 469996 48838 470008
rect 133414 469996 133420 470008
rect 48832 469968 133420 469996
rect 48832 469956 48838 469968
rect 133414 469956 133420 469968
rect 133472 469956 133478 470008
rect 235994 469956 236000 470008
rect 236052 469996 236058 470008
rect 365070 469996 365076 470008
rect 236052 469968 365076 469996
rect 236052 469956 236058 469968
rect 365070 469956 365076 469968
rect 365128 469956 365134 470008
rect 46198 469888 46204 469940
rect 46256 469928 46262 469940
rect 132862 469928 132868 469940
rect 46256 469900 132868 469928
rect 46256 469888 46262 469900
rect 132862 469888 132868 469900
rect 132920 469888 132926 469940
rect 178126 469888 178132 469940
rect 178184 469928 178190 469940
rect 214834 469928 214840 469940
rect 178184 469900 214840 469928
rect 178184 469888 178190 469900
rect 214834 469888 214840 469900
rect 214892 469888 214898 469940
rect 227806 469888 227812 469940
rect 227864 469928 227870 469940
rect 358170 469928 358176 469940
rect 227864 469900 358176 469928
rect 227864 469888 227870 469900
rect 358170 469888 358176 469900
rect 358228 469888 358234 469940
rect 43438 469820 43444 469872
rect 43496 469860 43502 469872
rect 132126 469860 132132 469872
rect 43496 469832 132132 469860
rect 43496 469820 43502 469832
rect 132126 469820 132132 469832
rect 132184 469820 132190 469872
rect 158806 469820 158812 469872
rect 158864 469860 158870 469872
rect 207658 469860 207664 469872
rect 158864 469832 207664 469860
rect 158864 469820 158870 469832
rect 207658 469820 207664 469832
rect 207716 469820 207722 469872
rect 229278 469820 229284 469872
rect 229336 469860 229342 469872
rect 374638 469860 374644 469872
rect 229336 469832 374644 469860
rect 229336 469820 229342 469832
rect 374638 469820 374644 469832
rect 374696 469820 374702 469872
rect 58526 469752 58532 469804
rect 58584 469792 58590 469804
rect 127158 469792 127164 469804
rect 58584 469764 127164 469792
rect 58584 469752 58590 469764
rect 127158 469752 127164 469764
rect 127216 469752 127222 469804
rect 58434 469684 58440 469736
rect 58492 469724 58498 469736
rect 126974 469724 126980 469736
rect 58492 469696 126980 469724
rect 58492 469684 58498 469696
rect 126974 469684 126980 469696
rect 127032 469684 127038 469736
rect 280890 469140 280896 469192
rect 280948 469180 280954 469192
rect 364058 469180 364064 469192
rect 280948 469152 364064 469180
rect 280948 469140 280954 469152
rect 364058 469140 364064 469152
rect 364116 469140 364122 469192
rect 264974 469072 264980 469124
rect 265032 469112 265038 469124
rect 358538 469112 358544 469124
rect 265032 469084 358544 469112
rect 265032 469072 265038 469084
rect 358538 469072 358544 469084
rect 358596 469072 358602 469124
rect 42150 469004 42156 469056
rect 42208 469044 42214 469056
rect 62206 469044 62212 469056
rect 42208 469016 62212 469044
rect 42208 469004 42214 469016
rect 62206 469004 62212 469016
rect 62264 469004 62270 469056
rect 273254 469004 273260 469056
rect 273312 469044 273318 469056
rect 372430 469044 372436 469056
rect 273312 469016 372436 469044
rect 273312 469004 273318 469016
rect 372430 469004 372436 469016
rect 372488 469004 372494 469056
rect 47946 468936 47952 468988
rect 48004 468976 48010 468988
rect 73890 468976 73896 468988
rect 48004 468948 73896 468976
rect 48004 468936 48010 468948
rect 73890 468936 73896 468948
rect 73948 468936 73954 468988
rect 270494 468936 270500 468988
rect 270552 468976 270558 468988
rect 373166 468976 373172 468988
rect 270552 468948 373172 468976
rect 270552 468936 270558 468948
rect 373166 468936 373172 468948
rect 373224 468936 373230 468988
rect 42518 468868 42524 468920
rect 42576 468908 42582 468920
rect 73982 468908 73988 468920
rect 42576 468880 73988 468908
rect 42576 468868 42582 468880
rect 73982 468868 73988 468880
rect 74040 468868 74046 468920
rect 259454 468868 259460 468920
rect 259512 468908 259518 468920
rect 370866 468908 370872 468920
rect 259512 468880 370872 468908
rect 259512 468868 259518 468880
rect 370866 468868 370872 468880
rect 370924 468868 370930 468920
rect 41322 468800 41328 468852
rect 41380 468840 41386 468852
rect 74074 468840 74080 468852
rect 41380 468812 74080 468840
rect 41380 468800 41386 468812
rect 74074 468800 74080 468812
rect 74132 468800 74138 468852
rect 256786 468800 256792 468852
rect 256844 468840 256850 468852
rect 370958 468840 370964 468852
rect 256844 468812 370964 468840
rect 256844 468800 256850 468812
rect 370958 468800 370964 468812
rect 371016 468800 371022 468852
rect 39850 468732 39856 468784
rect 39908 468772 39914 468784
rect 74166 468772 74172 468784
rect 39908 468744 74172 468772
rect 39908 468732 39914 468744
rect 74166 468732 74172 468744
rect 74224 468732 74230 468784
rect 175366 468732 175372 468784
rect 175424 468772 175430 468784
rect 207842 468772 207848 468784
rect 175424 468744 207848 468772
rect 175424 468732 175430 468744
rect 207842 468732 207848 468744
rect 207900 468732 207906 468784
rect 251266 468732 251272 468784
rect 251324 468772 251330 468784
rect 368014 468772 368020 468784
rect 251324 468744 368020 468772
rect 251324 468732 251330 468744
rect 368014 468732 368020 468744
rect 368072 468732 368078 468784
rect 43622 468664 43628 468716
rect 43680 468704 43686 468716
rect 103698 468704 103704 468716
rect 43680 468676 103704 468704
rect 43680 468664 43686 468676
rect 103698 468664 103704 468676
rect 103756 468664 103762 468716
rect 169018 468664 169024 468716
rect 169076 468704 169082 468716
rect 205910 468704 205916 468716
rect 169076 468676 205916 468704
rect 169076 468664 169082 468676
rect 205910 468664 205916 468676
rect 205968 468664 205974 468716
rect 244366 468664 244372 468716
rect 244424 468704 244430 468716
rect 366542 468704 366548 468716
rect 244424 468676 366548 468704
rect 244424 468664 244430 468676
rect 366542 468664 366548 468676
rect 366600 468664 366606 468716
rect 45370 468596 45376 468648
rect 45428 468636 45434 468648
rect 106458 468636 106464 468648
rect 45428 468608 106464 468636
rect 45428 468596 45434 468608
rect 106458 468596 106464 468608
rect 106516 468596 106522 468648
rect 165706 468596 165712 468648
rect 165764 468636 165770 468648
rect 218790 468636 218796 468648
rect 165764 468608 218796 468636
rect 165764 468596 165770 468608
rect 218790 468596 218796 468608
rect 218848 468596 218854 468648
rect 241514 468596 241520 468648
rect 241572 468636 241578 468648
rect 367830 468636 367836 468648
rect 241572 468608 367836 468636
rect 241572 468596 241578 468608
rect 367830 468596 367836 468608
rect 367888 468596 367894 468648
rect 45278 468528 45284 468580
rect 45336 468568 45342 468580
rect 106366 468568 106372 468580
rect 45336 468540 106372 468568
rect 45336 468528 45342 468540
rect 106366 468528 106372 468540
rect 106424 468528 106430 468580
rect 139486 468528 139492 468580
rect 139544 468568 139550 468580
rect 207474 468568 207480 468580
rect 139544 468540 207480 468568
rect 139544 468528 139550 468540
rect 207474 468528 207480 468540
rect 207532 468528 207538 468580
rect 227714 468528 227720 468580
rect 227772 468568 227778 468580
rect 360838 468568 360844 468580
rect 227772 468540 360844 468568
rect 227772 468528 227778 468540
rect 360838 468528 360844 468540
rect 360896 468528 360902 468580
rect 60826 468460 60832 468512
rect 60884 468500 60890 468512
rect 214190 468500 214196 468512
rect 60884 468472 214196 468500
rect 60884 468460 60890 468472
rect 214190 468460 214196 468472
rect 214248 468460 214254 468512
rect 226426 468460 226432 468512
rect 226484 468500 226490 468512
rect 376018 468500 376024 468512
rect 226484 468472 376024 468500
rect 226484 468460 226490 468472
rect 376018 468460 376024 468472
rect 376076 468460 376082 468512
rect 291470 468392 291476 468444
rect 291528 468432 291534 468444
rect 371694 468432 371700 468444
rect 291528 468404 371700 468432
rect 291528 468392 291534 468404
rect 371694 468392 371700 468404
rect 371752 468392 371758 468444
rect 88518 468120 88524 468172
rect 88576 468160 88582 468172
rect 89254 468160 89260 468172
rect 88576 468132 89260 468160
rect 88576 468120 88582 468132
rect 89254 468120 89260 468132
rect 89312 468120 89318 468172
rect 88426 467984 88432 468036
rect 88484 468024 88490 468036
rect 88702 468024 88708 468036
rect 88484 467996 88708 468024
rect 88484 467984 88490 467996
rect 88702 467984 88708 467996
rect 88760 467984 88766 468036
rect 274634 467712 274640 467764
rect 274692 467752 274698 467764
rect 358722 467752 358728 467764
rect 274692 467724 358728 467752
rect 274692 467712 274698 467724
rect 358722 467712 358728 467724
rect 358780 467712 358786 467764
rect 290182 467644 290188 467696
rect 290240 467684 290246 467696
rect 376662 467684 376668 467696
rect 290240 467656 376668 467684
rect 290240 467644 290246 467656
rect 376662 467644 376668 467656
rect 376720 467644 376726 467696
rect 285766 467576 285772 467628
rect 285824 467616 285830 467628
rect 286686 467616 286692 467628
rect 285824 467588 286692 467616
rect 285824 467576 285830 467588
rect 286686 467576 286692 467588
rect 286744 467576 286750 467628
rect 290550 467576 290556 467628
rect 290608 467616 290614 467628
rect 379238 467616 379244 467628
rect 290608 467588 379244 467616
rect 290608 467576 290614 467588
rect 379238 467576 379244 467588
rect 379296 467576 379302 467628
rect 266446 467508 266452 467560
rect 266504 467548 266510 467560
rect 359642 467548 359648 467560
rect 266504 467520 359648 467548
rect 266504 467508 266510 467520
rect 359642 467508 359648 467520
rect 359700 467508 359706 467560
rect 267918 467440 267924 467492
rect 267976 467480 267982 467492
rect 361390 467480 361396 467492
rect 267976 467452 361396 467480
rect 267976 467440 267982 467452
rect 361390 467440 361396 467452
rect 361448 467440 361454 467492
rect 256694 467372 256700 467424
rect 256752 467412 256758 467424
rect 365438 467412 365444 467424
rect 256752 467384 365444 467412
rect 256752 467372 256758 467384
rect 365438 467372 365444 467384
rect 365496 467372 365502 467424
rect 262306 467304 262312 467356
rect 262364 467344 262370 467356
rect 378962 467344 378968 467356
rect 262364 467316 378968 467344
rect 262364 467304 262370 467316
rect 378962 467304 378968 467316
rect 379020 467304 379026 467356
rect 57790 467236 57796 467288
rect 57848 467276 57854 467288
rect 113266 467276 113272 467288
rect 57848 467248 113272 467276
rect 57848 467236 57854 467248
rect 113266 467236 113272 467248
rect 113324 467236 113330 467288
rect 175274 467236 175280 467288
rect 175332 467276 175338 467288
rect 205082 467276 205088 467288
rect 175332 467248 205088 467276
rect 175332 467236 175338 467248
rect 205082 467236 205088 467248
rect 205140 467236 205146 467288
rect 242986 467236 242992 467288
rect 243044 467276 243050 467288
rect 373350 467276 373356 467288
rect 243044 467248 373356 467276
rect 243044 467236 243050 467248
rect 373350 467236 373356 467248
rect 373408 467236 373414 467288
rect 45186 467168 45192 467220
rect 45244 467208 45250 467220
rect 106274 467208 106280 467220
rect 45244 467180 106280 467208
rect 45244 467168 45250 467180
rect 106274 467168 106280 467180
rect 106332 467168 106338 467220
rect 160186 467168 160192 467220
rect 160244 467208 160250 467220
rect 202138 467208 202144 467220
rect 160244 467180 202144 467208
rect 160244 467168 160250 467180
rect 202138 467168 202144 467180
rect 202196 467168 202202 467220
rect 229186 467168 229192 467220
rect 229244 467208 229250 467220
rect 363690 467208 363696 467220
rect 229244 467180 363696 467208
rect 229244 467168 229250 467180
rect 363690 467168 363696 467180
rect 363748 467168 363754 467220
rect 59354 467100 59360 467152
rect 59412 467140 59418 467152
rect 179506 467140 179512 467152
rect 59412 467112 179512 467140
rect 59412 467100 59418 467112
rect 179506 467100 179512 467112
rect 179564 467100 179570 467152
rect 186406 467100 186412 467152
rect 186464 467140 186470 467152
rect 203702 467140 203708 467152
rect 186464 467112 203708 467140
rect 186464 467100 186470 467112
rect 203702 467100 203708 467112
rect 203760 467100 203766 467152
rect 207290 467100 207296 467152
rect 207348 467140 207354 467152
rect 217778 467140 217784 467152
rect 207348 467112 217784 467140
rect 207348 467100 207354 467112
rect 217778 467100 217784 467112
rect 217836 467100 217842 467152
rect 223666 467100 223672 467152
rect 223724 467140 223730 467152
rect 370498 467140 370504 467152
rect 223724 467112 370504 467140
rect 223724 467100 223730 467112
rect 370498 467100 370504 467112
rect 370556 467100 370562 467152
rect 50614 466352 50620 466404
rect 50672 466392 50678 466404
rect 82998 466392 83004 466404
rect 50672 466364 83004 466392
rect 50672 466352 50678 466364
rect 82998 466352 83004 466364
rect 83056 466352 83062 466404
rect 189166 466352 189172 466404
rect 189224 466392 189230 466404
rect 206278 466392 206284 466404
rect 189224 466364 206284 466392
rect 189224 466352 189230 466364
rect 206278 466352 206284 466364
rect 206336 466352 206342 466404
rect 49418 466284 49424 466336
rect 49476 466324 49482 466336
rect 82906 466324 82912 466336
rect 49476 466296 82912 466324
rect 49476 466284 49482 466296
rect 82906 466284 82912 466296
rect 82964 466284 82970 466336
rect 183646 466284 183652 466336
rect 183704 466324 183710 466336
rect 200758 466324 200764 466336
rect 183704 466296 200764 466324
rect 183704 466284 183710 466296
rect 200758 466284 200764 466296
rect 200816 466284 200822 466336
rect 298186 466284 298192 466336
rect 298244 466324 298250 466336
rect 357066 466324 357072 466336
rect 298244 466296 357072 466324
rect 298244 466284 298250 466296
rect 357066 466284 357072 466296
rect 357124 466284 357130 466336
rect 56502 466216 56508 466268
rect 56560 466256 56566 466268
rect 103606 466256 103612 466268
rect 56560 466228 103612 466256
rect 56560 466216 56566 466228
rect 103606 466216 103612 466228
rect 103664 466216 103670 466268
rect 183738 466216 183744 466268
rect 183796 466256 183802 466268
rect 205174 466256 205180 466268
rect 183796 466228 205180 466256
rect 183796 466216 183802 466228
rect 205174 466216 205180 466228
rect 205232 466216 205238 466268
rect 298278 466216 298284 466268
rect 298336 466256 298342 466268
rect 369854 466256 369860 466268
rect 298336 466228 369860 466256
rect 298336 466216 298342 466228
rect 369854 466216 369860 466228
rect 369912 466216 369918 466268
rect 51810 466148 51816 466200
rect 51868 466188 51874 466200
rect 99466 466188 99472 466200
rect 51868 466160 99472 466188
rect 51868 466148 51874 466160
rect 99466 466148 99472 466160
rect 99524 466148 99530 466200
rect 182450 466148 182456 466200
rect 182508 466188 182514 466200
rect 209314 466188 209320 466200
rect 182508 466160 209320 466188
rect 182508 466148 182514 466160
rect 209314 466148 209320 466160
rect 209372 466148 209378 466200
rect 299474 466148 299480 466200
rect 299532 466188 299538 466200
rect 373810 466188 373816 466200
rect 299532 466160 373816 466188
rect 299532 466148 299538 466160
rect 373810 466148 373816 466160
rect 373868 466148 373874 466200
rect 53190 466080 53196 466132
rect 53248 466120 53254 466132
rect 100938 466120 100944 466132
rect 53248 466092 100944 466120
rect 53248 466080 53254 466092
rect 100938 466080 100944 466092
rect 100996 466080 101002 466132
rect 189258 466080 189264 466132
rect 189316 466120 189322 466132
rect 216398 466120 216404 466132
rect 189316 466092 216404 466120
rect 189316 466080 189322 466092
rect 216398 466080 216404 466092
rect 216456 466080 216462 466132
rect 289814 466080 289820 466132
rect 289872 466120 289878 466132
rect 365530 466120 365536 466132
rect 289872 466092 365536 466120
rect 289872 466080 289878 466092
rect 365530 466080 365536 466092
rect 365588 466080 365594 466132
rect 53098 466012 53104 466064
rect 53156 466052 53162 466064
rect 100846 466052 100852 466064
rect 53156 466024 100852 466052
rect 53156 466012 53162 466024
rect 100846 466012 100852 466024
rect 100904 466012 100910 466064
rect 174078 466012 174084 466064
rect 174136 466052 174142 466064
rect 210786 466052 210792 466064
rect 174136 466024 210792 466052
rect 174136 466012 174142 466024
rect 210786 466012 210792 466024
rect 210844 466012 210850 466064
rect 288618 466012 288624 466064
rect 288676 466052 288682 466064
rect 368382 466052 368388 466064
rect 288676 466024 368388 466052
rect 288676 466012 288682 466024
rect 368382 466012 368388 466024
rect 368440 466012 368446 466064
rect 50246 465944 50252 465996
rect 50304 465984 50310 465996
rect 98178 465984 98184 465996
rect 50304 465956 98184 465984
rect 50304 465944 50310 465956
rect 98178 465944 98184 465956
rect 98236 465944 98242 465996
rect 139394 465944 139400 465996
rect 139452 465984 139458 465996
rect 197078 465984 197084 465996
rect 139452 465956 197084 465984
rect 139452 465944 139458 465956
rect 197078 465944 197084 465956
rect 197136 465944 197142 465996
rect 288526 465944 288532 465996
rect 288584 465984 288590 465996
rect 376570 465984 376576 465996
rect 288584 465956 376576 465984
rect 288584 465944 288590 465956
rect 376570 465944 376576 465956
rect 376628 465944 376634 465996
rect 58710 465876 58716 465928
rect 58768 465916 58774 465928
rect 110598 465916 110604 465928
rect 58768 465888 110604 465916
rect 58768 465876 58774 465888
rect 110598 465876 110604 465888
rect 110656 465876 110662 465928
rect 140958 465876 140964 465928
rect 141016 465916 141022 465928
rect 200574 465916 200580 465928
rect 141016 465888 200580 465916
rect 141016 465876 141022 465888
rect 200574 465876 200580 465888
rect 200632 465876 200638 465928
rect 249978 465876 249984 465928
rect 250036 465916 250042 465928
rect 366634 465916 366640 465928
rect 250036 465888 366640 465916
rect 250036 465876 250042 465888
rect 366634 465876 366640 465888
rect 366692 465876 366698 465928
rect 45002 465808 45008 465860
rect 45060 465848 45066 465860
rect 105078 465848 105084 465860
rect 45060 465820 105084 465848
rect 45060 465808 45066 465820
rect 105078 465808 105084 465820
rect 105136 465808 105142 465860
rect 140774 465808 140780 465860
rect 140832 465848 140838 465860
rect 203150 465848 203156 465860
rect 140832 465820 203156 465848
rect 140832 465808 140838 465820
rect 203150 465808 203156 465820
rect 203208 465808 203214 465860
rect 251174 465808 251180 465860
rect 251232 465848 251238 465860
rect 369302 465848 369308 465860
rect 251232 465820 369308 465848
rect 251232 465808 251238 465820
rect 369302 465808 369308 465820
rect 369360 465808 369366 465860
rect 45094 465740 45100 465792
rect 45152 465780 45158 465792
rect 104986 465780 104992 465792
rect 45152 465752 104992 465780
rect 45152 465740 45158 465752
rect 104986 465740 104992 465752
rect 105044 465740 105050 465792
rect 140866 465740 140872 465792
rect 140924 465780 140930 465792
rect 204438 465780 204444 465792
rect 140924 465752 204444 465780
rect 140924 465740 140930 465752
rect 204438 465740 204444 465752
rect 204496 465740 204502 465792
rect 240226 465740 240232 465792
rect 240284 465780 240290 465792
rect 373442 465780 373448 465792
rect 240284 465752 373448 465780
rect 240284 465740 240290 465752
rect 373442 465740 373448 465752
rect 373500 465740 373506 465792
rect 43530 465672 43536 465724
rect 43588 465712 43594 465724
rect 103514 465712 103520 465724
rect 43588 465684 103520 465712
rect 43588 465672 43594 465684
rect 103514 465672 103520 465684
rect 103572 465672 103578 465724
rect 125778 465672 125784 465724
rect 125836 465712 125842 465724
rect 201586 465712 201592 465724
rect 125836 465684 201592 465712
rect 125836 465672 125842 465684
rect 201586 465672 201592 465684
rect 201644 465672 201650 465724
rect 226334 465672 226340 465724
rect 226392 465712 226398 465724
rect 370590 465712 370596 465724
rect 226392 465684 370596 465712
rect 226392 465672 226398 465684
rect 370590 465672 370596 465684
rect 370648 465672 370654 465724
rect 52270 465604 52276 465656
rect 52328 465644 52334 465656
rect 82814 465644 82820 465656
rect 52328 465616 82820 465644
rect 52328 465604 52334 465616
rect 82814 465604 82820 465616
rect 82872 465604 82878 465656
rect 192018 465604 192024 465656
rect 192076 465644 192082 465656
rect 199562 465644 199568 465656
rect 192076 465616 199568 465644
rect 192076 465604 192082 465616
rect 199562 465604 199568 465616
rect 199620 465604 199626 465656
rect 203886 465644 203892 465656
rect 199764 465616 203892 465644
rect 44726 465536 44732 465588
rect 44784 465576 44790 465588
rect 65058 465576 65064 465588
rect 44784 465548 65064 465576
rect 44784 465536 44790 465548
rect 65058 465536 65064 465548
rect 65116 465536 65122 465588
rect 44818 465468 44824 465520
rect 44876 465508 44882 465520
rect 64966 465508 64972 465520
rect 44876 465480 64972 465508
rect 44876 465468 44882 465480
rect 64966 465468 64972 465480
rect 65024 465468 65030 465520
rect 190638 465468 190644 465520
rect 190696 465508 190702 465520
rect 199764 465508 199792 465616
rect 203886 465604 203892 465616
rect 203944 465604 203950 465656
rect 190696 465480 199792 465508
rect 190696 465468 190702 465480
rect 192662 465400 192668 465452
rect 192720 465440 192726 465452
rect 201034 465440 201040 465452
rect 192720 465412 201040 465440
rect 192720 465400 192726 465412
rect 201034 465400 201040 465412
rect 201092 465400 201098 465452
rect 288434 464924 288440 464976
rect 288492 464964 288498 464976
rect 357250 464964 357256 464976
rect 288492 464936 357256 464964
rect 288492 464924 288498 464936
rect 357250 464924 357256 464936
rect 357308 464924 357314 464976
rect 292666 464856 292672 464908
rect 292724 464896 292730 464908
rect 365622 464896 365628 464908
rect 292724 464868 365628 464896
rect 292724 464856 292730 464868
rect 365622 464856 365628 464868
rect 365680 464856 365686 464908
rect 292758 464788 292764 464840
rect 292816 464828 292822 464840
rect 366266 464828 366272 464840
rect 292816 464800 366272 464828
rect 292816 464788 292822 464800
rect 366266 464788 366272 464800
rect 366324 464788 366330 464840
rect 292574 464720 292580 464772
rect 292632 464760 292638 464772
rect 369026 464760 369032 464772
rect 292632 464732 369032 464760
rect 292632 464720 292638 464732
rect 369026 464720 369032 464732
rect 369084 464720 369090 464772
rect 284386 464652 284392 464704
rect 284444 464692 284450 464704
rect 362034 464692 362040 464704
rect 284444 464664 362040 464692
rect 284444 464652 284450 464664
rect 362034 464652 362040 464664
rect 362092 464652 362098 464704
rect 285674 464584 285680 464636
rect 285732 464624 285738 464636
rect 363506 464624 363512 464636
rect 285732 464596 363512 464624
rect 285732 464584 285738 464596
rect 363506 464584 363512 464596
rect 363564 464584 363570 464636
rect 291194 464516 291200 464568
rect 291252 464556 291258 464568
rect 370406 464556 370412 464568
rect 291252 464528 370412 464556
rect 291252 464516 291258 464528
rect 370406 464516 370412 464528
rect 370464 464516 370470 464568
rect 293954 464448 293960 464500
rect 294012 464488 294018 464500
rect 376846 464488 376852 464500
rect 294012 464460 376852 464488
rect 294012 464448 294018 464460
rect 376846 464448 376852 464460
rect 376904 464448 376910 464500
rect 57422 464380 57428 464432
rect 57480 464420 57486 464432
rect 114738 464420 114744 464432
rect 57480 464392 114744 464420
rect 57480 464380 57486 464392
rect 114738 464380 114744 464392
rect 114796 464380 114802 464432
rect 285858 464380 285864 464432
rect 285916 464420 285922 464432
rect 375374 464420 375380 464432
rect 285916 464392 375380 464420
rect 285916 464380 285922 464392
rect 375374 464380 375380 464392
rect 375432 464380 375438 464432
rect 42242 464312 42248 464364
rect 42300 464352 42306 464364
rect 102318 464352 102324 464364
rect 42300 464324 102324 464352
rect 42300 464312 42306 464324
rect 102318 464312 102324 464324
rect 102376 464312 102382 464364
rect 285766 464312 285772 464364
rect 285824 464352 285830 464364
rect 379330 464352 379336 464364
rect 285824 464324 379336 464352
rect 285824 464312 285830 464324
rect 379330 464312 379336 464324
rect 379388 464312 379394 464364
rect 56042 463632 56048 463684
rect 56100 463672 56106 463684
rect 86954 463672 86960 463684
rect 56100 463644 86960 463672
rect 56100 463632 56106 463644
rect 86954 463632 86960 463644
rect 87012 463632 87018 463684
rect 176838 463632 176844 463684
rect 176896 463672 176902 463684
rect 200850 463672 200856 463684
rect 176896 463644 200856 463672
rect 176896 463632 176902 463644
rect 200850 463632 200856 463644
rect 200908 463632 200914 463684
rect 287146 463632 287152 463684
rect 287204 463672 287210 463684
rect 360746 463672 360752 463684
rect 287204 463644 360752 463672
rect 287204 463632 287210 463644
rect 360746 463632 360752 463644
rect 360804 463632 360810 463684
rect 49326 463564 49332 463616
rect 49384 463604 49390 463616
rect 81618 463604 81624 463616
rect 49384 463576 81624 463604
rect 49384 463564 49390 463576
rect 81618 463564 81624 463576
rect 81676 463564 81682 463616
rect 193398 463564 193404 463616
rect 193456 463604 193462 463616
rect 217594 463604 217600 463616
rect 193456 463576 217600 463604
rect 193456 463564 193462 463576
rect 217594 463564 217600 463576
rect 217652 463564 217658 463616
rect 277486 463564 277492 463616
rect 277544 463604 277550 463616
rect 357158 463604 357164 463616
rect 277544 463576 357164 463604
rect 277544 463564 277550 463576
rect 357158 463564 357164 463576
rect 357216 463564 357222 463616
rect 56226 463496 56232 463548
rect 56284 463536 56290 463548
rect 88610 463536 88616 463548
rect 56284 463508 88616 463536
rect 56284 463496 56290 463508
rect 88610 463496 88616 463508
rect 88668 463496 88674 463548
rect 180978 463496 180984 463548
rect 181036 463536 181042 463548
rect 206646 463536 206652 463548
rect 181036 463508 206652 463536
rect 181036 463496 181042 463508
rect 206646 463496 206652 463508
rect 206704 463496 206710 463548
rect 276198 463496 276204 463548
rect 276256 463536 276262 463548
rect 361482 463536 361488 463548
rect 276256 463508 361488 463536
rect 276256 463496 276262 463508
rect 361482 463496 361488 463508
rect 361540 463496 361546 463548
rect 54938 463428 54944 463480
rect 54996 463468 55002 463480
rect 87138 463468 87144 463480
rect 54996 463440 87144 463468
rect 54996 463428 55002 463440
rect 87138 463428 87144 463440
rect 87196 463428 87202 463480
rect 178034 463428 178040 463480
rect 178092 463468 178098 463480
rect 216122 463468 216128 463480
rect 178092 463440 216128 463468
rect 178092 463428 178098 463440
rect 216122 463428 216128 463440
rect 216180 463428 216186 463480
rect 276106 463428 276112 463480
rect 276164 463468 276170 463480
rect 364886 463468 364892 463480
rect 276164 463440 364892 463468
rect 276164 463428 276170 463440
rect 364886 463428 364892 463440
rect 364944 463428 364950 463480
rect 53282 463360 53288 463412
rect 53340 463400 53346 463412
rect 85666 463400 85672 463412
rect 53340 463372 85672 463400
rect 53340 463360 53346 463372
rect 85666 463360 85672 463372
rect 85724 463360 85730 463412
rect 169754 463360 169760 463412
rect 169812 463400 169818 463412
rect 209130 463400 209136 463412
rect 169812 463372 209136 463400
rect 169812 463360 169818 463372
rect 209130 463360 209136 463372
rect 209188 463360 209194 463412
rect 280246 463360 280252 463412
rect 280304 463400 280310 463412
rect 370314 463400 370320 463412
rect 280304 463372 370320 463400
rect 280304 463360 280310 463372
rect 370314 463360 370320 463372
rect 370372 463360 370378 463412
rect 55122 463292 55128 463344
rect 55180 463332 55186 463344
rect 88518 463332 88524 463344
rect 55180 463304 88524 463332
rect 55180 463292 55186 463304
rect 88518 463292 88524 463304
rect 88576 463292 88582 463344
rect 161566 463292 161572 463344
rect 161624 463332 161630 463344
rect 204990 463332 204996 463344
rect 161624 463304 204996 463332
rect 161624 463292 161630 463304
rect 204990 463292 204996 463304
rect 205048 463292 205054 463344
rect 277578 463292 277584 463344
rect 277636 463332 277642 463344
rect 368934 463332 368940 463344
rect 277636 463304 368940 463332
rect 277636 463292 277642 463304
rect 368934 463292 368940 463304
rect 368992 463292 368998 463344
rect 55030 463224 55036 463276
rect 55088 463264 55094 463276
rect 88426 463264 88432 463276
rect 55088 463236 88432 463264
rect 55088 463224 55094 463236
rect 88426 463224 88432 463236
rect 88484 463224 88490 463276
rect 161474 463224 161480 463276
rect 161532 463264 161538 463276
rect 210694 463264 210700 463276
rect 161532 463236 210700 463264
rect 161532 463224 161538 463236
rect 210694 463224 210700 463236
rect 210752 463224 210758 463276
rect 267826 463224 267832 463276
rect 267884 463264 267890 463276
rect 359550 463264 359556 463276
rect 267884 463236 359556 463264
rect 267884 463224 267890 463236
rect 359550 463224 359556 463236
rect 359608 463224 359614 463276
rect 56134 463156 56140 463208
rect 56192 463196 56198 463208
rect 89806 463196 89812 463208
rect 56192 463168 89812 463196
rect 56192 463156 56198 463168
rect 89806 463156 89812 463168
rect 89864 463156 89870 463208
rect 142338 463156 142344 463208
rect 142396 463196 142402 463208
rect 200482 463196 200488 463208
rect 142396 463168 200488 463196
rect 142396 463156 142402 463168
rect 200482 463156 200488 463168
rect 200540 463156 200546 463208
rect 278958 463156 278964 463208
rect 279016 463196 279022 463208
rect 374454 463196 374460 463208
rect 279016 463168 374460 463196
rect 279016 463156 279022 463168
rect 374454 463156 374460 463168
rect 374512 463156 374518 463208
rect 57606 463088 57612 463140
rect 57664 463128 57670 463140
rect 113358 463128 113364 463140
rect 57664 463100 113364 463128
rect 57664 463088 57670 463100
rect 113358 463088 113364 463100
rect 113416 463088 113422 463140
rect 142246 463088 142252 463140
rect 142304 463128 142310 463140
rect 208578 463128 208584 463140
rect 142304 463100 208584 463128
rect 142304 463088 142310 463100
rect 208578 463088 208584 463100
rect 208636 463088 208642 463140
rect 249886 463088 249892 463140
rect 249944 463128 249950 463140
rect 365254 463128 365260 463140
rect 249944 463100 365260 463128
rect 249944 463088 249950 463100
rect 365254 463088 365260 463100
rect 365312 463088 365318 463140
rect 53374 463020 53380 463072
rect 53432 463060 53438 463072
rect 87046 463060 87052 463072
rect 53432 463032 87052 463060
rect 53432 463020 53438 463032
rect 87046 463020 87052 463032
rect 87104 463020 87110 463072
rect 107746 463020 107752 463072
rect 107804 463060 107810 463072
rect 201862 463060 201868 463072
rect 107804 463032 201868 463060
rect 107804 463020 107810 463032
rect 201862 463020 201868 463032
rect 201920 463020 201926 463072
rect 249794 463020 249800 463072
rect 249852 463060 249858 463072
rect 372062 463060 372068 463072
rect 249852 463032 372068 463060
rect 249852 463020 249858 463032
rect 372062 463020 372068 463032
rect 372120 463020 372126 463072
rect 53006 462952 53012 463004
rect 53064 462992 53070 463004
rect 100754 462992 100760 463004
rect 53064 462964 100760 462992
rect 53064 462952 53070 462964
rect 100754 462952 100760 462964
rect 100812 462952 100818 463004
rect 109126 462952 109132 463004
rect 109184 462992 109190 463004
rect 205634 462992 205640 463004
rect 109184 462964 205640 462992
rect 109184 462952 109190 462964
rect 205634 462952 205640 462964
rect 205692 462952 205698 463004
rect 240134 462952 240140 463004
rect 240192 462992 240198 463004
rect 362494 462992 362500 463004
rect 240192 462964 362500 462992
rect 240192 462952 240198 462964
rect 362494 462952 362500 462964
rect 362552 462952 362558 463004
rect 54846 462884 54852 462936
rect 54904 462924 54910 462936
rect 85574 462924 85580 462936
rect 54904 462896 85580 462924
rect 54904 462884 54910 462896
rect 85574 462884 85580 462896
rect 85632 462884 85638 462936
rect 189074 462884 189080 462936
rect 189132 462924 189138 462936
rect 212258 462924 212264 462936
rect 189132 462896 212264 462924
rect 189132 462884 189138 462896
rect 212258 462884 212264 462896
rect 212316 462884 212322 462936
rect 284294 462884 284300 462936
rect 284352 462924 284358 462936
rect 357802 462924 357808 462936
rect 284352 462896 357808 462924
rect 284352 462884 284358 462896
rect 357802 462884 357808 462896
rect 357860 462884 357866 462936
rect 47578 462816 47584 462868
rect 47636 462856 47642 462868
rect 64874 462856 64880 462868
rect 47636 462828 64880 462856
rect 47636 462816 47642 462828
rect 64874 462816 64880 462828
rect 64932 462816 64938 462868
rect 182358 462816 182364 462868
rect 182416 462856 182422 462868
rect 202322 462856 202328 462868
rect 182416 462828 202328 462856
rect 182416 462816 182422 462828
rect 202322 462816 202328 462828
rect 202380 462816 202386 462868
rect 47670 462748 47676 462800
rect 47728 462788 47734 462800
rect 63678 462788 63684 462800
rect 47728 462760 63684 462788
rect 47728 462748 47734 462760
rect 63678 462748 63684 462760
rect 63736 462748 63742 462800
rect 193306 462748 193312 462800
rect 193364 462788 193370 462800
rect 213086 462788 213092 462800
rect 193364 462760 213092 462788
rect 193364 462748 193370 462760
rect 213086 462748 213092 462760
rect 213144 462748 213150 462800
rect 133138 462272 133144 462324
rect 133196 462312 133202 462324
rect 178310 462312 178316 462324
rect 133196 462284 178316 462312
rect 133196 462272 133202 462284
rect 178310 462272 178316 462284
rect 178368 462272 178374 462324
rect 185578 462136 185584 462188
rect 185636 462176 185642 462188
rect 203242 462176 203248 462188
rect 185636 462148 203248 462176
rect 185636 462136 185642 462148
rect 203242 462136 203248 462148
rect 203300 462136 203306 462188
rect 190546 462068 190552 462120
rect 190604 462108 190610 462120
rect 208946 462108 208952 462120
rect 190604 462080 208952 462108
rect 190604 462068 190610 462080
rect 208946 462068 208952 462080
rect 209004 462068 209010 462120
rect 282914 462068 282920 462120
rect 282972 462108 282978 462120
rect 358078 462108 358084 462120
rect 282972 462080 358084 462108
rect 282972 462068 282978 462080
rect 358078 462068 358084 462080
rect 358136 462068 358142 462120
rect 176746 462000 176752 462052
rect 176804 462040 176810 462052
rect 202230 462040 202236 462052
rect 176804 462012 202236 462040
rect 176804 462000 176810 462012
rect 202230 462000 202236 462012
rect 202288 462000 202294 462052
rect 296714 462000 296720 462052
rect 296772 462040 296778 462052
rect 373994 462040 374000 462052
rect 296772 462012 374000 462040
rect 296772 462000 296778 462012
rect 373994 462000 374000 462012
rect 374052 462000 374058 462052
rect 184934 461932 184940 461984
rect 184992 461972 184998 461984
rect 213270 461972 213276 461984
rect 184992 461944 213276 461972
rect 184992 461932 184998 461944
rect 213270 461932 213276 461944
rect 213328 461932 213334 461984
rect 278866 461932 278872 461984
rect 278924 461972 278930 461984
rect 357986 461972 357992 461984
rect 278924 461944 357992 461972
rect 278924 461932 278930 461944
rect 357986 461932 357992 461944
rect 358044 461932 358050 461984
rect 182266 461864 182272 461916
rect 182324 461904 182330 461916
rect 212166 461904 212172 461916
rect 182324 461876 212172 461904
rect 182324 461864 182330 461876
rect 212166 461864 212172 461876
rect 212224 461864 212230 461916
rect 277394 461864 277400 461916
rect 277452 461904 277458 461916
rect 366174 461904 366180 461916
rect 277452 461876 366180 461904
rect 277452 461864 277458 461876
rect 366174 461864 366180 461876
rect 366232 461864 366238 461916
rect 180886 461796 180892 461848
rect 180944 461836 180950 461848
rect 213362 461836 213368 461848
rect 180944 461808 213368 461836
rect 180944 461796 180950 461808
rect 213362 461796 213368 461808
rect 213420 461796 213426 461848
rect 253934 461796 253940 461848
rect 253992 461836 253998 461848
rect 363966 461836 363972 461848
rect 253992 461808 363972 461836
rect 253992 461796 253998 461808
rect 363966 461796 363972 461808
rect 364024 461796 364030 461848
rect 179506 461728 179512 461780
rect 179564 461768 179570 461780
rect 212902 461768 212908 461780
rect 179564 461740 212908 461768
rect 179564 461728 179570 461740
rect 212902 461728 212908 461740
rect 212960 461728 212966 461780
rect 260834 461728 260840 461780
rect 260892 461768 260898 461780
rect 376386 461768 376392 461780
rect 260892 461740 376392 461768
rect 260892 461728 260898 461740
rect 376386 461728 376392 461740
rect 376444 461728 376450 461780
rect 57698 461660 57704 461712
rect 57756 461700 57762 461712
rect 111886 461700 111892 461712
rect 57756 461672 111892 461700
rect 57756 461660 57762 461672
rect 111886 461660 111892 461672
rect 111944 461660 111950 461712
rect 158714 461660 158720 461712
rect 158772 461700 158778 461712
rect 206462 461700 206468 461712
rect 158772 461672 206468 461700
rect 158772 461660 158778 461672
rect 206462 461660 206468 461672
rect 206520 461660 206526 461712
rect 252554 461660 252560 461712
rect 252612 461700 252618 461712
rect 373626 461700 373632 461712
rect 252612 461672 373632 461700
rect 252612 461660 252618 461672
rect 373626 461660 373632 461672
rect 373684 461660 373690 461712
rect 52178 461592 52184 461644
rect 52236 461632 52242 461644
rect 71038 461632 71044 461644
rect 52236 461604 71044 461632
rect 52236 461592 52242 461604
rect 71038 461592 71044 461604
rect 71096 461592 71102 461644
rect 107654 461592 107660 461644
rect 107712 461632 107718 461644
rect 198274 461632 198280 461644
rect 107712 461604 198280 461632
rect 107712 461592 107718 461604
rect 198274 461592 198280 461604
rect 198332 461592 198338 461644
rect 252646 461592 252652 461644
rect 252704 461632 252710 461644
rect 376202 461632 376208 461644
rect 252704 461604 376208 461632
rect 252704 461592 252710 461604
rect 376202 461592 376208 461604
rect 376260 461592 376266 461644
rect 498194 461116 498200 461168
rect 498252 461156 498258 461168
rect 517698 461156 517704 461168
rect 498252 461128 517704 461156
rect 498252 461116 498258 461128
rect 517698 461116 517704 461128
rect 517756 461116 517762 461168
rect 339770 461048 339776 461100
rect 339828 461088 339834 461100
rect 356974 461088 356980 461100
rect 339828 461060 356980 461088
rect 339828 461048 339834 461060
rect 356974 461048 356980 461060
rect 357032 461088 357038 461100
rect 357032 461060 489914 461088
rect 357032 461048 357038 461060
rect 178310 460980 178316 461032
rect 178368 461020 178374 461032
rect 201954 461020 201960 461032
rect 178368 460992 201960 461020
rect 178368 460980 178374 460992
rect 201954 460980 201960 460992
rect 202012 461020 202018 461032
rect 338298 461020 338304 461032
rect 202012 460992 338304 461020
rect 202012 460980 202018 460992
rect 338298 460980 338304 460992
rect 338356 461020 338362 461032
rect 362954 461020 362960 461032
rect 338356 460992 362960 461020
rect 338356 460980 338362 460992
rect 362954 460980 362960 460992
rect 363012 461020 363018 461032
rect 489886 461020 489914 461060
rect 499850 461020 499856 461032
rect 363012 460992 364334 461020
rect 489886 460992 499856 461020
rect 363012 460980 363018 460992
rect 190914 460912 190920 460964
rect 190972 460952 190978 460964
rect 207014 460952 207020 460964
rect 190972 460924 207020 460952
rect 190972 460912 190978 460924
rect 207014 460912 207020 460924
rect 207072 460912 207078 460964
rect 212902 460912 212908 460964
rect 212960 460952 212966 460964
rect 339770 460952 339776 460964
rect 212960 460924 339776 460952
rect 212960 460912 212966 460924
rect 339770 460912 339776 460924
rect 339828 460912 339834 460964
rect 350994 460912 351000 460964
rect 351052 460952 351058 460964
rect 360194 460952 360200 460964
rect 351052 460924 360200 460952
rect 351052 460912 351058 460924
rect 360194 460912 360200 460924
rect 360252 460912 360258 460964
rect 364306 460952 364334 460992
rect 499850 460980 499856 460992
rect 499908 461020 499914 461032
rect 517606 461020 517612 461032
rect 499908 460992 517612 461020
rect 499908 460980 499914 460992
rect 517606 460980 517612 460992
rect 517664 460980 517670 461032
rect 498194 460952 498200 460964
rect 364306 460924 498200 460952
rect 498194 460912 498200 460924
rect 498252 460912 498258 460964
rect 510890 460912 510896 460964
rect 510948 460952 510954 460964
rect 517514 460952 517520 460964
rect 510948 460924 517520 460952
rect 510948 460912 510954 460924
rect 517514 460912 517520 460924
rect 517572 460912 517578 460964
rect 50706 460844 50712 460896
rect 50764 460884 50770 460896
rect 80054 460884 80060 460896
rect 50764 460856 80060 460884
rect 50764 460844 50770 460856
rect 80054 460844 80060 460856
rect 80112 460844 80118 460896
rect 287054 460844 287060 460896
rect 287112 460884 287118 460896
rect 367646 460884 367652 460896
rect 287112 460856 367652 460884
rect 287112 460844 287118 460856
rect 367646 460844 367652 460856
rect 367704 460844 367710 460896
rect 53742 460776 53748 460828
rect 53800 460816 53806 460828
rect 78766 460816 78772 460828
rect 53800 460788 78772 460816
rect 53800 460776 53806 460788
rect 78766 460776 78772 460788
rect 78824 460776 78830 460828
rect 179414 460776 179420 460828
rect 179472 460816 179478 460828
rect 218974 460816 218980 460828
rect 179472 460788 218980 460816
rect 179472 460776 179478 460788
rect 218974 460776 218980 460788
rect 219032 460776 219038 460828
rect 262214 460776 262220 460828
rect 262272 460816 262278 460828
rect 361114 460816 361120 460828
rect 262272 460788 361120 460816
rect 262272 460776 262278 460788
rect 361114 460776 361120 460788
rect 361172 460776 361178 460828
rect 53650 460708 53656 460760
rect 53708 460748 53714 460760
rect 66346 460748 66352 460760
rect 53708 460720 66352 460748
rect 53708 460708 53714 460720
rect 66346 460708 66352 460720
rect 66404 460708 66410 460760
rect 258166 460708 258172 460760
rect 258224 460748 258230 460760
rect 363874 460748 363880 460760
rect 258224 460720 363880 460748
rect 258224 460708 258230 460720
rect 363874 460708 363880 460720
rect 363932 460708 363938 460760
rect 43254 460640 43260 460692
rect 43312 460680 43318 460692
rect 60734 460680 60740 460692
rect 43312 460652 60740 460680
rect 43312 460640 43318 460652
rect 60734 460640 60740 460652
rect 60792 460640 60798 460692
rect 183554 460640 183560 460692
rect 183612 460680 183618 460692
rect 203794 460680 203800 460692
rect 183612 460652 203800 460680
rect 183612 460640 183618 460652
rect 203794 460640 203800 460652
rect 203852 460640 203858 460692
rect 267734 460640 267740 460692
rect 267792 460680 267798 460692
rect 373718 460680 373724 460692
rect 267792 460652 373724 460680
rect 267792 460640 267798 460652
rect 373718 460640 373724 460652
rect 373776 460640 373782 460692
rect 43346 460572 43352 460624
rect 43404 460612 43410 460624
rect 62114 460612 62120 460624
rect 43404 460584 62120 460612
rect 43404 460572 43410 460584
rect 62114 460572 62120 460584
rect 62172 460572 62178 460624
rect 187786 460572 187792 460624
rect 187844 460612 187850 460624
rect 209406 460612 209412 460624
rect 187844 460584 209412 460612
rect 187844 460572 187850 460584
rect 209406 460572 209412 460584
rect 209464 460572 209470 460624
rect 248598 460572 248604 460624
rect 248656 460612 248662 460624
rect 367922 460612 367928 460624
rect 248656 460584 367928 460612
rect 248656 460572 248662 460584
rect 367922 460572 367928 460584
rect 367980 460572 367986 460624
rect 49510 460504 49516 460556
rect 49568 460544 49574 460556
rect 70394 460544 70400 460556
rect 49568 460516 70400 460544
rect 49568 460504 49574 460516
rect 70394 460504 70400 460516
rect 70452 460504 70458 460556
rect 180794 460504 180800 460556
rect 180852 460544 180858 460556
rect 205266 460544 205272 460556
rect 180852 460516 205272 460544
rect 180852 460504 180858 460516
rect 205266 460504 205272 460516
rect 205324 460504 205330 460556
rect 248414 460504 248420 460556
rect 248472 460544 248478 460556
rect 370774 460544 370780 460556
rect 248472 460516 370780 460544
rect 248472 460504 248478 460516
rect 370774 460504 370780 460516
rect 370832 460504 370838 460556
rect 39942 460436 39948 460488
rect 40000 460476 40006 460488
rect 66254 460476 66260 460488
rect 40000 460448 66260 460476
rect 40000 460436 40006 460448
rect 66254 460436 66260 460448
rect 66312 460436 66318 460488
rect 193214 460436 193220 460488
rect 193272 460476 193278 460488
rect 219158 460476 219164 460488
rect 193272 460448 219164 460476
rect 193272 460436 193278 460448
rect 219158 460436 219164 460448
rect 219216 460436 219222 460488
rect 248506 460436 248512 460488
rect 248564 460476 248570 460488
rect 373534 460476 373540 460488
rect 248564 460448 373540 460476
rect 248564 460436 248570 460448
rect 373534 460436 373540 460448
rect 373592 460436 373598 460488
rect 44910 460368 44916 460420
rect 44968 460408 44974 460420
rect 73798 460408 73804 460420
rect 44968 460380 73804 460408
rect 44968 460368 44974 460380
rect 73798 460368 73804 460380
rect 73856 460368 73862 460420
rect 168466 460368 168472 460420
rect 168524 460408 168530 460420
rect 206370 460408 206376 460420
rect 168524 460380 206376 460408
rect 168524 460368 168530 460380
rect 206370 460368 206376 460380
rect 206428 460368 206434 460420
rect 244274 460368 244280 460420
rect 244332 460408 244338 460420
rect 369394 460408 369400 460420
rect 244332 460380 369400 460408
rect 244332 460368 244338 460380
rect 369394 460368 369400 460380
rect 369452 460368 369458 460420
rect 49602 460300 49608 460352
rect 49660 460340 49666 460352
rect 78858 460340 78864 460352
rect 49660 460312 78864 460340
rect 49660 460300 49666 460312
rect 78858 460300 78864 460312
rect 78916 460300 78922 460352
rect 165614 460300 165620 460352
rect 165672 460340 165678 460352
rect 203610 460340 203616 460352
rect 165672 460312 203616 460340
rect 165672 460300 165678 460312
rect 203610 460300 203616 460312
rect 203668 460300 203674 460352
rect 247218 460300 247224 460352
rect 247276 460340 247282 460352
rect 376110 460340 376116 460352
rect 247276 460312 376116 460340
rect 247276 460300 247282 460312
rect 376110 460300 376116 460312
rect 376168 460300 376174 460352
rect 50522 460232 50528 460284
rect 50580 460272 50586 460284
rect 92566 460272 92572 460284
rect 50580 460244 92572 460272
rect 50580 460232 50586 460244
rect 92566 460232 92572 460244
rect 92624 460232 92630 460284
rect 247126 460232 247132 460284
rect 247184 460272 247190 460284
rect 376294 460272 376300 460284
rect 247184 460244 376300 460272
rect 247184 460232 247190 460244
rect 376294 460232 376300 460244
rect 376352 460232 376358 460284
rect 44082 460164 44088 460216
rect 44140 460204 44146 460216
rect 71774 460204 71780 460216
rect 44140 460176 71780 460204
rect 44140 460164 44146 460176
rect 71774 460164 71780 460176
rect 71832 460164 71838 460216
rect 72418 460164 72424 460216
rect 72476 460204 72482 460216
rect 199010 460204 199016 460216
rect 72476 460176 199016 460204
rect 72476 460164 72482 460176
rect 199010 460164 199016 460176
rect 199068 460164 199074 460216
rect 237374 460164 237380 460216
rect 237432 460204 237438 460216
rect 374730 460204 374736 460216
rect 237432 460176 374736 460204
rect 237432 460164 237438 460176
rect 374730 460164 374736 460176
rect 374788 460164 374794 460216
rect 59262 460096 59268 460148
rect 59320 460136 59326 460148
rect 67726 460136 67732 460148
rect 59320 460108 67732 460136
rect 59320 460096 59326 460108
rect 67726 460096 67732 460108
rect 67784 460096 67790 460148
rect 59906 460028 59912 460080
rect 59964 460068 59970 460080
rect 68278 460068 68284 460080
rect 59964 460040 68284 460068
rect 59964 460028 59970 460040
rect 68278 460028 68284 460040
rect 68336 460028 68342 460080
rect 194594 459620 194600 459672
rect 194652 459660 194658 459672
rect 199470 459660 199476 459672
rect 194652 459632 199476 459660
rect 194652 459620 194658 459632
rect 199470 459620 199476 459632
rect 199528 459620 199534 459672
rect 215754 459620 215760 459672
rect 215812 459660 215818 459672
rect 220906 459660 220912 459672
rect 215812 459632 220912 459660
rect 215812 459620 215818 459632
rect 220906 459620 220912 459632
rect 220964 459620 220970 459672
rect 218606 459552 218612 459604
rect 218664 459592 218670 459604
rect 220998 459592 221004 459604
rect 218664 459564 221004 459592
rect 218664 459552 218670 459564
rect 220998 459552 221004 459564
rect 221056 459552 221062 459604
rect 187694 459484 187700 459536
rect 187752 459524 187758 459536
rect 200942 459524 200948 459536
rect 187752 459496 200948 459524
rect 187752 459484 187758 459496
rect 200942 459484 200948 459496
rect 201000 459484 201006 459536
rect 191834 459416 191840 459468
rect 191892 459456 191898 459468
rect 205358 459456 205364 459468
rect 191892 459428 205364 459456
rect 191892 459416 191898 459428
rect 205358 459416 205364 459428
rect 205416 459416 205422 459468
rect 295334 459416 295340 459468
rect 295392 459456 295398 459468
rect 357894 459456 357900 459468
rect 295392 459428 357900 459456
rect 295392 459416 295398 459428
rect 357894 459416 357900 459428
rect 357952 459416 357958 459468
rect 190454 459348 190460 459400
rect 190512 459388 190518 459400
rect 208026 459388 208032 459400
rect 190512 459360 208032 459388
rect 190512 459348 190518 459360
rect 208026 459348 208032 459360
rect 208084 459348 208090 459400
rect 298094 459348 298100 459400
rect 298152 459388 298158 459400
rect 364242 459388 364248 459400
rect 298152 459360 364248 459388
rect 298152 459348 298158 459360
rect 364242 459348 364248 459360
rect 364300 459348 364306 459400
rect 58894 459280 58900 459332
rect 58952 459320 58958 459332
rect 92474 459320 92480 459332
rect 58952 459292 92480 459320
rect 58952 459280 58958 459292
rect 92474 459280 92480 459292
rect 92532 459280 92538 459332
rect 182174 459280 182180 459332
rect 182232 459320 182238 459332
rect 207934 459320 207940 459332
rect 182232 459292 207940 459320
rect 182232 459280 182238 459292
rect 207934 459280 207940 459292
rect 207992 459280 207998 459332
rect 281534 459280 281540 459332
rect 281592 459320 281598 459332
rect 359734 459320 359740 459332
rect 281592 459292 359740 459320
rect 281592 459280 281598 459292
rect 359734 459280 359740 459292
rect 359792 459280 359798 459332
rect 55950 459212 55956 459264
rect 56008 459252 56014 459264
rect 89898 459252 89904 459264
rect 56008 459224 89904 459252
rect 56008 459212 56014 459224
rect 89898 459212 89904 459224
rect 89956 459212 89962 459264
rect 173986 459212 173992 459264
rect 174044 459252 174050 459264
rect 206738 459252 206744 459264
rect 174044 459224 206744 459252
rect 174044 459212 174050 459224
rect 206738 459212 206744 459224
rect 206796 459212 206802 459264
rect 280154 459212 280160 459264
rect 280212 459252 280218 459264
rect 362126 459252 362132 459264
rect 280212 459224 362132 459252
rect 280212 459212 280218 459224
rect 362126 459212 362132 459224
rect 362184 459212 362190 459264
rect 57514 459144 57520 459196
rect 57572 459184 57578 459196
rect 111978 459184 111984 459196
rect 57572 459156 111984 459184
rect 57572 459144 57578 459156
rect 111978 459144 111984 459156
rect 112036 459144 112042 459196
rect 176654 459144 176660 459196
rect 176712 459184 176718 459196
rect 210878 459184 210884 459196
rect 176712 459156 210884 459184
rect 176712 459144 176718 459156
rect 210878 459144 210884 459156
rect 210936 459144 210942 459196
rect 276014 459144 276020 459196
rect 276072 459184 276078 459196
rect 367554 459184 367560 459196
rect 276072 459156 367560 459184
rect 276072 459144 276078 459156
rect 367554 459144 367560 459156
rect 367612 459144 367618 459196
rect 54662 459076 54668 459128
rect 54720 459116 54726 459128
rect 117498 459116 117504 459128
rect 54720 459088 117504 459116
rect 54720 459076 54726 459088
rect 117498 459076 117504 459088
rect 117556 459076 117562 459128
rect 173894 459076 173900 459128
rect 173952 459116 173958 459128
rect 216214 459116 216220 459128
rect 173952 459088 216220 459116
rect 173952 459076 173958 459088
rect 216214 459076 216220 459088
rect 216272 459076 216278 459128
rect 271874 459076 271880 459128
rect 271932 459116 271938 459128
rect 364794 459116 364800 459128
rect 271932 459088 364800 459116
rect 271932 459076 271938 459088
rect 364794 459076 364800 459088
rect 364852 459076 364858 459128
rect 51718 459008 51724 459060
rect 51776 459048 51782 459060
rect 121454 459048 121460 459060
rect 51776 459020 121460 459048
rect 51776 459008 51782 459020
rect 121454 459008 121460 459020
rect 121512 459008 121518 459060
rect 125594 459008 125600 459060
rect 125652 459048 125658 459060
rect 197538 459048 197544 459060
rect 125652 459020 197544 459048
rect 125652 459008 125658 459020
rect 197538 459008 197544 459020
rect 197596 459008 197602 459060
rect 263594 459008 263600 459060
rect 263652 459048 263658 459060
rect 366910 459048 366916 459060
rect 263652 459020 366916 459048
rect 263652 459008 263658 459020
rect 366910 459008 366916 459020
rect 366968 459008 366974 459060
rect 55766 458940 55772 458992
rect 55824 458980 55830 458992
rect 130010 458980 130016 458992
rect 55824 458952 130016 458980
rect 55824 458940 55830 458952
rect 130010 458940 130016 458952
rect 130068 458940 130074 458992
rect 136634 458940 136640 458992
rect 136692 458980 136698 458992
rect 199102 458980 199108 458992
rect 136692 458952 199108 458980
rect 136692 458940 136698 458952
rect 199102 458940 199108 458952
rect 199160 458940 199166 458992
rect 258074 458940 258080 458992
rect 258132 458980 258138 458992
rect 372338 458980 372344 458992
rect 258132 458952 372344 458980
rect 258132 458940 258138 458952
rect 372338 458940 372344 458952
rect 372396 458940 372402 458992
rect 54478 458872 54484 458924
rect 54536 458912 54542 458924
rect 134058 458912 134064 458924
rect 54536 458884 134064 458912
rect 54536 458872 54542 458884
rect 134058 458872 134064 458884
rect 134116 458872 134122 458924
rect 142154 458872 142160 458924
rect 142212 458912 142218 458924
rect 211338 458912 211344 458924
rect 142212 458884 211344 458912
rect 142212 458872 142218 458884
rect 211338 458872 211344 458884
rect 211396 458872 211402 458924
rect 242894 458872 242900 458924
rect 242952 458912 242958 458924
rect 374822 458912 374828 458924
rect 242952 458884 374828 458912
rect 242952 458872 242958 458884
rect 374822 458872 374828 458884
rect 374880 458872 374886 458924
rect 52914 458804 52920 458856
rect 52972 458844 52978 458856
rect 99558 458844 99564 458856
rect 52972 458816 99564 458844
rect 52972 458804 52978 458816
rect 99558 458804 99564 458816
rect 99616 458804 99622 458856
rect 109310 458804 109316 458856
rect 109368 458844 109374 458856
rect 197630 458844 197636 458856
rect 109368 458816 197636 458844
rect 109368 458804 109374 458816
rect 197630 458804 197636 458816
rect 197688 458804 197694 458856
rect 247034 458804 247040 458856
rect 247092 458844 247098 458856
rect 379054 458844 379060 458856
rect 247092 458816 379060 458844
rect 247092 458804 247098 458816
rect 379054 458804 379060 458816
rect 379112 458804 379118 458856
rect 191926 458736 191932 458788
rect 191984 458776 191990 458788
rect 202414 458776 202420 458788
rect 191984 458748 202420 458776
rect 191984 458736 191990 458748
rect 202414 458736 202420 458748
rect 202472 458736 202478 458788
rect 199010 458328 199016 458380
rect 199068 458368 199074 458380
rect 199068 458340 354674 458368
rect 199068 458328 199074 458340
rect 46014 458260 46020 458312
rect 46072 458300 46078 458312
rect 354646 458300 354674 458340
rect 358814 458300 358820 458312
rect 46072 458272 200114 458300
rect 354646 458272 358820 458300
rect 46072 458260 46078 458272
rect 200086 458232 200114 458272
rect 358814 458260 358820 458272
rect 358872 458300 358878 458312
rect 516594 458300 516600 458312
rect 358872 458272 516600 458300
rect 358872 458260 358878 458272
rect 516594 458260 516600 458272
rect 516652 458260 516658 458312
rect 207382 458232 207388 458244
rect 200086 458204 207388 458232
rect 207382 458192 207388 458204
rect 207440 458232 207446 458244
rect 208118 458232 208124 458244
rect 207440 458204 208124 458232
rect 207440 458192 207446 458204
rect 208118 458192 208124 458204
rect 208176 458192 208182 458244
rect 204346 457444 204352 457496
rect 204404 457484 204410 457496
rect 217870 457484 217876 457496
rect 204404 457456 217876 457484
rect 204404 457444 204410 457456
rect 217870 457444 217876 457456
rect 217928 457444 217934 457496
rect 50706 456084 50712 456136
rect 50764 456124 50770 456136
rect 50982 456124 50988 456136
rect 50764 456096 50988 456124
rect 50764 456084 50770 456096
rect 50982 456084 50988 456096
rect 51040 456084 51046 456136
rect 356606 456084 356612 456136
rect 356664 456124 356670 456136
rect 356974 456124 356980 456136
rect 356664 456096 356980 456124
rect 356664 456084 356670 456096
rect 356974 456084 356980 456096
rect 357032 456084 357038 456136
rect 519538 454656 519544 454708
rect 519596 454696 519602 454708
rect 580258 454696 580264 454708
rect 519596 454668 580264 454696
rect 519596 454656 519602 454668
rect 580258 454656 580264 454668
rect 580316 454656 580322 454708
rect 54386 414196 54392 414248
rect 54444 414236 54450 414248
rect 55582 414236 55588 414248
rect 54444 414208 55588 414236
rect 54444 414196 54450 414208
rect 55582 414196 55588 414208
rect 55640 414196 55646 414248
rect 205818 413924 205824 413976
rect 205876 413964 205882 413976
rect 207290 413964 207296 413976
rect 205876 413936 207296 413964
rect 205876 413924 205882 413936
rect 207290 413924 207296 413936
rect 207348 413924 207354 413976
rect 208118 413244 208124 413296
rect 208176 413284 208182 413296
rect 216950 413284 216956 413296
rect 208176 413256 216956 413284
rect 208176 413244 208182 413256
rect 216950 413244 216956 413256
rect 217008 413244 217014 413296
rect 46014 412564 46020 412616
rect 46072 412604 46078 412616
rect 56962 412604 56968 412616
rect 46072 412576 56968 412604
rect 46072 412564 46078 412576
rect 56962 412564 56968 412576
rect 57020 412564 57026 412616
rect 54386 411884 54392 411936
rect 54444 411924 54450 411936
rect 58434 411924 58440 411936
rect 54444 411896 58440 411924
rect 54444 411884 54450 411896
rect 58434 411884 58440 411896
rect 58492 411884 58498 411936
rect 199654 411884 199660 411936
rect 199712 411924 199718 411936
rect 205818 411924 205824 411936
rect 199712 411896 205824 411924
rect 199712 411884 199718 411896
rect 205818 411884 205824 411896
rect 205876 411884 205882 411936
rect 363506 411884 363512 411936
rect 363564 411924 363570 411936
rect 377030 411924 377036 411936
rect 363564 411896 377036 411924
rect 363564 411884 363570 411896
rect 377030 411884 377036 411896
rect 377088 411884 377094 411936
rect 2958 411204 2964 411256
rect 3016 411244 3022 411256
rect 14458 411244 14464 411256
rect 3016 411216 14464 411244
rect 3016 411204 3022 411216
rect 14458 411204 14464 411216
rect 14516 411204 14522 411256
rect 57054 410796 57060 410848
rect 57112 410836 57118 410848
rect 58434 410836 58440 410848
rect 57112 410808 58440 410836
rect 57112 410796 57118 410808
rect 58434 410796 58440 410808
rect 58492 410796 58498 410848
rect 198090 410524 198096 410576
rect 198148 410564 198154 410576
rect 199286 410564 199292 410576
rect 198148 410536 199292 410564
rect 198148 410524 198154 410536
rect 199286 410524 199292 410536
rect 199344 410524 199350 410576
rect 362034 410524 362040 410576
rect 362092 410564 362098 410576
rect 377214 410564 377220 410576
rect 362092 410536 377220 410564
rect 362092 410524 362098 410536
rect 377214 410524 377220 410536
rect 377272 410524 377278 410576
rect 44634 409844 44640 409896
rect 44692 409884 44698 409896
rect 57054 409884 57060 409896
rect 44692 409856 57060 409884
rect 44692 409844 44698 409856
rect 57054 409844 57060 409856
rect 57112 409844 57118 409896
rect 53558 409776 53564 409828
rect 53616 409816 53622 409828
rect 56870 409816 56876 409828
rect 53616 409788 56876 409816
rect 53616 409776 53622 409788
rect 56870 409776 56876 409788
rect 56928 409776 56934 409828
rect 205726 409096 205732 409148
rect 205784 409136 205790 409148
rect 216674 409136 216680 409148
rect 205784 409108 216680 409136
rect 205784 409096 205790 409108
rect 216674 409096 216680 409108
rect 216732 409096 216738 409148
rect 360010 409096 360016 409148
rect 360068 409136 360074 409148
rect 377214 409136 377220 409148
rect 360068 409108 377220 409136
rect 360068 409096 360074 409108
rect 377214 409096 377220 409108
rect 377272 409096 377278 409148
rect 47486 408484 47492 408536
rect 47544 408524 47550 408536
rect 57054 408524 57060 408536
rect 47544 408496 57060 408524
rect 47544 408484 47550 408496
rect 57054 408484 57060 408496
rect 57112 408484 57118 408536
rect 373902 407804 373908 407856
rect 373960 407844 373966 407856
rect 376846 407844 376852 407856
rect 373960 407816 376852 407844
rect 373960 407804 373966 407816
rect 376846 407804 376852 407816
rect 376904 407804 376910 407856
rect 207290 407736 207296 407788
rect 207348 407776 207354 407788
rect 216674 407776 216680 407788
rect 207348 407748 216680 407776
rect 207348 407736 207354 407748
rect 216674 407736 216680 407748
rect 216732 407736 216738 407788
rect 357802 407736 357808 407788
rect 357860 407776 357866 407788
rect 377122 407776 377128 407788
rect 357860 407748 377128 407776
rect 357860 407736 357866 407748
rect 377122 407736 377128 407748
rect 377180 407736 377186 407788
rect 47394 407124 47400 407176
rect 47452 407164 47458 407176
rect 56962 407164 56968 407176
rect 47452 407136 56968 407164
rect 47452 407124 47458 407136
rect 56962 407124 56968 407136
rect 57020 407124 57026 407176
rect 359918 406376 359924 406428
rect 359976 406416 359982 406428
rect 377214 406416 377220 406428
rect 359976 406388 377220 406416
rect 359976 406376 359982 406388
rect 377214 406376 377220 406388
rect 377272 406376 377278 406428
rect 53558 405696 53564 405748
rect 53616 405736 53622 405748
rect 57054 405736 57060 405748
rect 53616 405708 57060 405736
rect 53616 405696 53622 405708
rect 57054 405696 57060 405708
rect 57112 405696 57118 405748
rect 375926 405628 375932 405680
rect 375984 405668 375990 405680
rect 376754 405668 376760 405680
rect 375984 405640 376760 405668
rect 375984 405628 375990 405640
rect 376754 405628 376760 405640
rect 376812 405628 376818 405680
rect 377674 405628 377680 405680
rect 377732 405668 377738 405680
rect 378594 405668 378600 405680
rect 377732 405640 378600 405668
rect 377732 405628 377738 405640
rect 378594 405628 378600 405640
rect 378652 405628 378658 405680
rect 358078 404948 358084 405000
rect 358136 404988 358142 405000
rect 377582 404988 377588 405000
rect 358136 404960 377588 404988
rect 358136 404948 358142 404960
rect 377582 404948 377588 404960
rect 377640 404948 377646 405000
rect 51626 404336 51632 404388
rect 51684 404376 51690 404388
rect 57054 404376 57060 404388
rect 51684 404348 57060 404376
rect 51684 404336 51690 404348
rect 57054 404336 57060 404348
rect 57112 404336 57118 404388
rect 51718 404268 51724 404320
rect 51776 404308 51782 404320
rect 53834 404308 53840 404320
rect 51776 404280 53840 404308
rect 51776 404268 51782 404280
rect 53834 404268 53840 404280
rect 53892 404268 53898 404320
rect 359826 403588 359832 403640
rect 359884 403628 359890 403640
rect 377674 403628 377680 403640
rect 359884 403600 377680 403628
rect 359884 403588 359890 403600
rect 377674 403588 377680 403600
rect 377732 403588 377738 403640
rect 52362 402976 52368 403028
rect 52420 403016 52426 403028
rect 56962 403016 56968 403028
rect 52420 402988 56968 403016
rect 52420 402976 52426 402988
rect 56962 402976 56968 402988
rect 57020 402976 57026 403028
rect 199654 393932 199660 393984
rect 199712 393972 199718 393984
rect 214190 393972 214196 393984
rect 199712 393944 214196 393972
rect 199712 393932 199718 393944
rect 214190 393932 214196 393944
rect 214248 393932 214254 393984
rect 198182 393388 198188 393440
rect 198240 393428 198246 393440
rect 198240 393400 200712 393428
rect 198240 393388 198246 393400
rect 198366 393320 198372 393372
rect 198424 393360 198430 393372
rect 200574 393360 200580 393372
rect 198424 393332 200580 393360
rect 198424 393320 198430 393332
rect 200574 393320 200580 393332
rect 200632 393320 200638 393372
rect 200574 393184 200580 393236
rect 200632 393224 200638 393236
rect 200684 393224 200712 393400
rect 200632 393196 200712 393224
rect 200632 393184 200638 393196
rect 199562 391212 199568 391264
rect 199620 391252 199626 391264
rect 211522 391252 211528 391264
rect 199620 391224 211528 391252
rect 199620 391212 199626 391224
rect 211522 391212 211528 391224
rect 211580 391212 211586 391264
rect 377398 388696 377404 388748
rect 377456 388736 377462 388748
rect 377766 388736 377772 388748
rect 377456 388708 377772 388736
rect 377456 388696 377462 388708
rect 377766 388696 377772 388708
rect 377824 388696 377830 388748
rect 216766 388560 216772 388612
rect 216824 388600 216830 388612
rect 216950 388600 216956 388612
rect 216824 388572 216956 388600
rect 216824 388560 216830 388572
rect 216950 388560 216956 388572
rect 217008 388560 217014 388612
rect 520918 388424 520924 388476
rect 520976 388464 520982 388476
rect 580350 388464 580356 388476
rect 520976 388436 580356 388464
rect 520976 388424 520982 388436
rect 580350 388424 580356 388436
rect 580408 388424 580414 388476
rect 46106 384956 46112 385008
rect 46164 384996 46170 385008
rect 56962 384996 56968 385008
rect 46164 384968 56968 384996
rect 46164 384956 46170 384968
rect 56962 384956 56968 384968
rect 57020 384956 57026 385008
rect 209498 384956 209504 385008
rect 209556 384996 209562 385008
rect 216674 384996 216680 385008
rect 209556 384968 216680 384996
rect 209556 384956 209562 384968
rect 216674 384956 216680 384968
rect 216732 384956 216738 385008
rect 359734 384956 359740 385008
rect 359792 384996 359798 385008
rect 376938 384996 376944 385008
rect 359792 384968 376944 384996
rect 359792 384956 359798 384968
rect 376938 384956 376944 384968
rect 376996 384956 377002 385008
rect 56962 383596 56968 383648
rect 57020 383636 57026 383648
rect 57146 383636 57152 383648
rect 57020 383608 57152 383636
rect 57020 383596 57026 383608
rect 57146 383596 57152 383608
rect 57204 383596 57210 383648
rect 57238 383596 57244 383648
rect 57296 383596 57302 383648
rect 57330 383596 57336 383648
rect 57388 383596 57394 383648
rect 207014 383596 207020 383648
rect 207072 383636 207078 383648
rect 216674 383636 216680 383648
rect 207072 383608 216680 383636
rect 207072 383596 207078 383608
rect 216674 383596 216680 383608
rect 216732 383596 216738 383648
rect 360194 383596 360200 383648
rect 360252 383636 360258 383648
rect 376938 383636 376944 383648
rect 360252 383608 376944 383636
rect 360252 383596 360258 383608
rect 376938 383596 376944 383608
rect 376996 383596 377002 383648
rect 57256 383568 57284 383596
rect 57164 383540 57284 383568
rect 57164 383512 57192 383540
rect 57146 383460 57152 383512
rect 57204 383460 57210 383512
rect 57238 383460 57244 383512
rect 57296 383500 57302 383512
rect 57348 383500 57376 383596
rect 359642 383528 359648 383580
rect 359700 383568 359706 383580
rect 376846 383568 376852 383580
rect 359700 383540 376852 383568
rect 359700 383528 359706 383540
rect 376846 383528 376852 383540
rect 376904 383528 376910 383580
rect 57296 383472 57376 383500
rect 57296 383460 57302 383472
rect 216858 383460 216864 383512
rect 216916 383500 216922 383512
rect 217318 383500 217324 383512
rect 216916 383472 217324 383500
rect 216916 383460 216922 383472
rect 217318 383460 217324 383472
rect 217376 383460 217382 383512
rect 212258 383324 212264 383376
rect 212316 383364 212322 383376
rect 216858 383364 216864 383376
rect 212316 383336 216864 383364
rect 212316 383324 212322 383336
rect 216858 383324 216864 383336
rect 216916 383324 216922 383376
rect 358078 382236 358084 382288
rect 358136 382276 358142 382288
rect 360194 382276 360200 382288
rect 358136 382248 360200 382276
rect 358136 382236 358142 382248
rect 360194 382236 360200 382248
rect 360252 382236 360258 382288
rect 42702 382168 42708 382220
rect 42760 382208 42766 382220
rect 56870 382208 56876 382220
rect 42760 382180 56876 382208
rect 42760 382168 42766 382180
rect 56870 382168 56876 382180
rect 56928 382208 56934 382220
rect 57238 382208 57244 382220
rect 56928 382180 57244 382208
rect 56928 382168 56934 382180
rect 57238 382168 57244 382180
rect 57296 382168 57302 382220
rect 212626 379788 212632 379840
rect 212684 379828 212690 379840
rect 213454 379828 213460 379840
rect 212684 379800 213460 379828
rect 212684 379788 212690 379800
rect 213454 379788 213460 379800
rect 213512 379788 213518 379840
rect 51718 379516 51724 379568
rect 51776 379556 51782 379568
rect 53834 379556 53840 379568
rect 51776 379528 53840 379556
rect 51776 379516 51782 379528
rect 53834 379516 53840 379528
rect 53892 379516 53898 379568
rect 218054 378768 218060 378820
rect 218112 378808 218118 378820
rect 218330 378808 218336 378820
rect 218112 378780 218336 378808
rect 218112 378768 218118 378780
rect 218330 378768 218336 378780
rect 218388 378768 218394 378820
rect 57146 378564 57152 378616
rect 57204 378604 57210 378616
rect 57330 378604 57336 378616
rect 57204 378576 57336 378604
rect 57204 378564 57210 378576
rect 57330 378564 57336 378576
rect 57388 378564 57394 378616
rect 53558 375368 53564 375420
rect 53616 375368 53622 375420
rect 53576 375340 53604 375368
rect 53742 375340 53748 375352
rect 53576 375312 53748 375340
rect 53742 375300 53748 375312
rect 53800 375300 53806 375352
rect 197170 375300 197176 375352
rect 197228 375340 197234 375352
rect 198182 375340 198188 375352
rect 197228 375312 198188 375340
rect 197228 375300 197234 375312
rect 198182 375300 198188 375312
rect 198240 375300 198246 375352
rect 217226 375300 217232 375352
rect 217284 375340 217290 375352
rect 217778 375340 217784 375352
rect 217284 375312 217784 375340
rect 217284 375300 217290 375312
rect 217778 375300 217784 375312
rect 217836 375300 217842 375352
rect 51626 375028 51632 375080
rect 51684 375068 51690 375080
rect 217226 375068 217232 375080
rect 51684 375040 217232 375068
rect 51684 375028 51690 375040
rect 217226 375028 217232 375040
rect 217284 375028 217290 375080
rect 53742 374960 53748 375012
rect 53800 375000 53806 375012
rect 217318 375000 217324 375012
rect 53800 374972 217324 375000
rect 53800 374960 53806 374972
rect 217318 374960 217324 374972
rect 217376 374960 217382 375012
rect 375190 374960 375196 375012
rect 375248 375000 375254 375012
rect 380894 375000 380900 375012
rect 375248 374972 380900 375000
rect 375248 374960 375254 374972
rect 380894 374960 380900 374972
rect 380952 374960 380958 375012
rect 56502 374892 56508 374944
rect 56560 374932 56566 374944
rect 60734 374932 60740 374944
rect 56560 374904 60740 374932
rect 56560 374892 56566 374904
rect 60734 374892 60740 374904
rect 60792 374892 60798 374944
rect 200206 374756 200212 374808
rect 200264 374796 200270 374808
rect 304258 374796 304264 374808
rect 200264 374768 304264 374796
rect 200264 374756 200270 374768
rect 304258 374756 304264 374768
rect 304316 374756 304322 374808
rect 200666 374688 200672 374740
rect 200724 374728 200730 374740
rect 304994 374728 305000 374740
rect 200724 374700 305000 374728
rect 200724 374688 200730 374700
rect 304994 374688 305000 374700
rect 305052 374688 305058 374740
rect 375374 374688 375380 374740
rect 375432 374728 375438 374740
rect 375432 374700 379514 374728
rect 375432 374688 375438 374700
rect 201678 374620 201684 374672
rect 201736 374660 201742 374672
rect 311802 374660 311808 374672
rect 201736 374632 311808 374660
rect 201736 374620 201742 374632
rect 311802 374620 311808 374632
rect 311860 374620 311866 374672
rect 377398 374620 377404 374672
rect 377456 374660 377462 374672
rect 377766 374660 377772 374672
rect 377456 374632 377772 374660
rect 377456 374620 377462 374632
rect 377766 374620 377772 374632
rect 377824 374620 377830 374672
rect 379486 374660 379514 374700
rect 404170 374660 404176 374672
rect 379486 374632 404176 374660
rect 404170 374620 404176 374632
rect 404228 374620 404234 374672
rect 165982 374552 165988 374604
rect 166040 374592 166046 374604
rect 200482 374592 200488 374604
rect 166040 374564 200488 374592
rect 166040 374552 166046 374564
rect 200482 374552 200488 374564
rect 200540 374552 200546 374604
rect 201770 374552 201776 374604
rect 201828 374592 201834 374604
rect 320910 374592 320916 374604
rect 201828 374564 320916 374592
rect 201828 374552 201834 374564
rect 320910 374552 320916 374564
rect 320968 374552 320974 374604
rect 371050 374552 371056 374604
rect 371108 374592 371114 374604
rect 407758 374592 407764 374604
rect 371108 374564 407764 374592
rect 371108 374552 371114 374564
rect 407758 374552 407764 374564
rect 407816 374552 407822 374604
rect 158530 374484 158536 374536
rect 158588 374524 158594 374536
rect 204438 374524 204444 374536
rect 158588 374496 204444 374524
rect 158588 374484 158594 374496
rect 204438 374484 204444 374496
rect 204496 374484 204502 374536
rect 215938 374484 215944 374536
rect 215996 374524 216002 374536
rect 220906 374524 220912 374536
rect 215996 374496 220912 374524
rect 215996 374484 216002 374496
rect 220906 374484 220912 374496
rect 220964 374484 220970 374536
rect 373718 374484 373724 374536
rect 373776 374524 373782 374536
rect 410702 374524 410708 374536
rect 373776 374496 410708 374524
rect 373776 374484 373782 374496
rect 410702 374484 410708 374496
rect 410760 374484 410766 374536
rect 156506 374416 156512 374468
rect 156564 374456 156570 374468
rect 203150 374456 203156 374468
rect 156564 374428 203156 374456
rect 156564 374416 156570 374428
rect 203150 374416 203156 374428
rect 203208 374416 203214 374468
rect 208486 374416 208492 374468
rect 208544 374456 208550 374468
rect 210234 374456 210240 374468
rect 208544 374428 210240 374456
rect 208544 374416 208550 374428
rect 210234 374416 210240 374428
rect 210292 374456 210298 374468
rect 221550 374456 221556 374468
rect 210292 374428 221556 374456
rect 210292 374416 210298 374428
rect 221550 374416 221556 374428
rect 221608 374416 221614 374468
rect 380894 374416 380900 374468
rect 380952 374456 380958 374468
rect 425054 374456 425060 374468
rect 380952 374428 425060 374456
rect 380952 374416 380958 374428
rect 425054 374416 425060 374428
rect 425112 374416 425118 374468
rect 163406 374348 163412 374400
rect 163464 374388 163470 374400
rect 211338 374388 211344 374400
rect 163464 374360 211344 374388
rect 163464 374348 163470 374360
rect 211338 374348 211344 374360
rect 211396 374348 211402 374400
rect 240686 374348 240692 374400
rect 240744 374388 240750 374400
rect 244274 374388 244280 374400
rect 240744 374360 244280 374388
rect 240744 374348 240750 374360
rect 244274 374348 244280 374360
rect 244332 374348 244338 374400
rect 378042 374348 378048 374400
rect 378100 374388 378106 374400
rect 443086 374388 443092 374400
rect 378100 374360 443092 374388
rect 378100 374348 378106 374360
rect 443086 374348 443092 374360
rect 443144 374348 443150 374400
rect 160922 374280 160928 374332
rect 160980 374320 160986 374332
rect 208578 374320 208584 374332
rect 160980 374292 208584 374320
rect 160980 374280 160986 374292
rect 208578 374280 208584 374292
rect 208636 374280 208642 374332
rect 211706 374280 211712 374332
rect 211764 374320 211770 374332
rect 221642 374320 221648 374332
rect 211764 374292 221648 374320
rect 211764 374280 211770 374292
rect 221642 374280 221648 374292
rect 221700 374280 221706 374332
rect 240778 374280 240784 374332
rect 240836 374320 240842 374332
rect 247586 374320 247592 374332
rect 240836 374292 247592 374320
rect 240836 374280 240842 374292
rect 247586 374280 247592 374292
rect 247644 374280 247650 374332
rect 367002 374280 367008 374332
rect 367060 374320 367066 374332
rect 436002 374320 436008 374332
rect 367060 374292 436008 374320
rect 367060 374280 367066 374292
rect 436002 374280 436008 374292
rect 436060 374280 436066 374332
rect 146202 374212 146208 374264
rect 146260 374252 146266 374264
rect 207474 374252 207480 374264
rect 146260 374224 207480 374252
rect 146260 374212 146266 374224
rect 207474 374212 207480 374224
rect 207532 374212 207538 374264
rect 208394 374212 208400 374264
rect 208452 374252 208458 374264
rect 218054 374252 218060 374264
rect 208452 374224 218060 374252
rect 208452 374212 208458 374224
rect 218054 374212 218060 374224
rect 218112 374212 218118 374264
rect 219342 374212 219348 374264
rect 219400 374252 219406 374264
rect 265250 374252 265256 374264
rect 219400 374224 265256 374252
rect 219400 374212 219406 374224
rect 265250 374212 265256 374224
rect 265308 374212 265314 374264
rect 369670 374212 369676 374264
rect 369728 374252 369734 374264
rect 438486 374252 438492 374264
rect 369728 374224 438492 374252
rect 369728 374212 369734 374224
rect 438486 374212 438492 374224
rect 438544 374212 438550 374264
rect 143534 374144 143540 374196
rect 143592 374184 143598 374196
rect 205910 374184 205916 374196
rect 143592 374156 205916 374184
rect 143592 374144 143598 374156
rect 205910 374144 205916 374156
rect 205968 374144 205974 374196
rect 217594 374144 217600 374196
rect 217652 374184 217658 374196
rect 270494 374184 270500 374196
rect 217652 374156 270500 374184
rect 217652 374144 217658 374156
rect 270494 374144 270500 374156
rect 270552 374144 270558 374196
rect 372430 374144 372436 374196
rect 372488 374184 372494 374196
rect 440326 374184 440332 374196
rect 372488 374156 440332 374184
rect 372488 374144 372494 374156
rect 440326 374144 440332 374156
rect 440384 374144 440390 374196
rect 56962 374076 56968 374128
rect 57020 374116 57026 374128
rect 105446 374116 105452 374128
rect 57020 374088 105452 374116
rect 57020 374076 57026 374088
rect 105446 374076 105452 374088
rect 105504 374076 105510 374128
rect 148962 374076 148968 374128
rect 149020 374116 149026 374128
rect 197078 374116 197084 374128
rect 149020 374088 197084 374116
rect 149020 374076 149026 374088
rect 197078 374076 197084 374088
rect 197136 374076 197142 374128
rect 199470 374076 199476 374128
rect 199528 374116 199534 374128
rect 283006 374116 283012 374128
rect 199528 374088 283012 374116
rect 199528 374076 199534 374088
rect 283006 374076 283012 374088
rect 283064 374076 283070 374128
rect 364794 374076 364800 374128
rect 364852 374116 364858 374128
rect 433610 374116 433616 374128
rect 364852 374088 433616 374116
rect 364852 374076 364858 374088
rect 433610 374076 433616 374088
rect 433668 374076 433674 374128
rect 54478 374008 54484 374060
rect 54536 374048 54542 374060
rect 116026 374048 116032 374060
rect 54536 374020 116032 374048
rect 54536 374008 54542 374020
rect 116026 374008 116032 374020
rect 116084 374008 116090 374060
rect 140958 374008 140964 374060
rect 141016 374048 141022 374060
rect 203242 374048 203248 374060
rect 141016 374020 203248 374048
rect 141016 374008 141022 374020
rect 203242 374008 203248 374020
rect 203300 374008 203306 374060
rect 209958 374008 209964 374060
rect 210016 374048 210022 374060
rect 211706 374048 211712 374060
rect 210016 374020 211712 374048
rect 210016 374008 210022 374020
rect 211706 374008 211712 374020
rect 211764 374008 211770 374060
rect 218054 374008 218060 374060
rect 218112 374048 218118 374060
rect 219066 374048 219072 374060
rect 218112 374020 219072 374048
rect 218112 374008 218118 374020
rect 219066 374008 219072 374020
rect 219124 374048 219130 374060
rect 240686 374048 240692 374060
rect 219124 374020 240692 374048
rect 219124 374008 219130 374020
rect 240686 374008 240692 374020
rect 240744 374008 240750 374060
rect 240870 374008 240876 374060
rect 240928 374048 240934 374060
rect 244734 374048 244740 374060
rect 240928 374020 244740 374048
rect 240928 374008 240934 374020
rect 244734 374008 244740 374020
rect 244792 374008 244798 374060
rect 250622 374008 250628 374060
rect 250680 374048 250686 374060
rect 253474 374048 253480 374060
rect 250680 374020 253480 374048
rect 250680 374008 250686 374020
rect 253474 374008 253480 374020
rect 253532 374008 253538 374060
rect 364150 374008 364156 374060
rect 364208 374048 364214 374060
rect 450998 374048 451004 374060
rect 364208 374020 451004 374048
rect 364208 374008 364214 374020
rect 450998 374008 451004 374020
rect 451056 374008 451062 374060
rect 44634 373940 44640 373992
rect 44692 373980 44698 373992
rect 217042 373980 217048 373992
rect 44692 373952 217048 373980
rect 44692 373940 44698 373952
rect 217042 373940 217048 373952
rect 217100 373940 217106 373992
rect 377950 373940 377956 373992
rect 378008 373980 378014 373992
rect 421006 373980 421012 373992
rect 378008 373952 421012 373980
rect 378008 373940 378014 373952
rect 421006 373940 421012 373952
rect 421064 373940 421070 373992
rect 47394 373872 47400 373924
rect 47452 373912 47458 373924
rect 216858 373912 216864 373924
rect 47452 373884 216864 373912
rect 47452 373872 47458 373884
rect 216858 373872 216864 373884
rect 216916 373872 216922 373924
rect 376478 373872 376484 373924
rect 376536 373912 376542 373924
rect 423030 373912 423036 373924
rect 376536 373884 423036 373912
rect 376536 373872 376542 373884
rect 423030 373872 423036 373884
rect 423088 373872 423094 373924
rect 47762 373804 47768 373856
rect 47820 373844 47826 373856
rect 96062 373844 96068 373856
rect 47820 373816 96068 373844
rect 47820 373804 47826 373816
rect 96062 373804 96068 373816
rect 96120 373804 96126 373856
rect 139210 373804 139216 373856
rect 139268 373844 139274 373856
rect 200390 373844 200396 373856
rect 139268 373816 200396 373844
rect 139268 373804 139274 373816
rect 200390 373804 200396 373816
rect 200448 373804 200454 373856
rect 215386 373804 215392 373856
rect 215444 373844 215450 373856
rect 219342 373844 219348 373856
rect 215444 373816 219348 373844
rect 215444 373804 215450 373816
rect 219342 373804 219348 373816
rect 219400 373804 219406 373856
rect 372614 373804 372620 373856
rect 372672 373844 372678 373856
rect 373718 373844 373724 373856
rect 372672 373816 373724 373844
rect 372672 373804 372678 373816
rect 373718 373804 373724 373816
rect 373776 373844 373782 373856
rect 426894 373844 426900 373856
rect 373776 373816 426900 373844
rect 373776 373804 373782 373816
rect 426894 373804 426900 373816
rect 426952 373804 426958 373856
rect 57330 373736 57336 373788
rect 57388 373776 57394 373788
rect 118326 373776 118332 373788
rect 57388 373748 118332 373776
rect 57388 373736 57394 373748
rect 118326 373736 118332 373748
rect 118384 373736 118390 373788
rect 136450 373736 136456 373788
rect 136508 373776 136514 373788
rect 200298 373776 200304 373788
rect 136508 373748 200304 373776
rect 136508 373736 136514 373748
rect 200298 373736 200304 373748
rect 200356 373736 200362 373788
rect 361390 373736 361396 373788
rect 361448 373776 361454 373788
rect 416038 373776 416044 373788
rect 361448 373748 416044 373776
rect 361448 373736 361454 373748
rect 416038 373736 416044 373748
rect 416096 373736 416102 373788
rect 43438 373668 43444 373720
rect 43496 373708 43502 373720
rect 103514 373708 103520 373720
rect 43496 373680 103520 373708
rect 43496 373668 43502 373680
rect 103514 373668 103520 373680
rect 103572 373668 103578 373720
rect 133690 373668 133696 373720
rect 133748 373708 133754 373720
rect 199286 373708 199292 373720
rect 133748 373680 199292 373708
rect 133748 373668 133754 373680
rect 199286 373668 199292 373680
rect 199344 373668 199350 373720
rect 371786 373668 371792 373720
rect 371844 373708 371850 373720
rect 430574 373708 430580 373720
rect 371844 373680 430580 373708
rect 371844 373668 371850 373680
rect 430574 373668 430580 373680
rect 430632 373668 430638 373720
rect 51534 373600 51540 373652
rect 51592 373640 51598 373652
rect 113542 373640 113548 373652
rect 51592 373612 113548 373640
rect 51592 373600 51598 373612
rect 113542 373600 113548 373612
rect 113600 373600 113606 373652
rect 131022 373600 131028 373652
rect 131080 373640 131086 373652
rect 199102 373640 199108 373652
rect 131080 373612 199108 373640
rect 131080 373600 131086 373612
rect 199102 373600 199108 373612
rect 199160 373600 199166 373652
rect 204254 373600 204260 373652
rect 204312 373640 204318 373652
rect 219250 373640 219256 373652
rect 204312 373612 219256 373640
rect 204312 373600 204318 373612
rect 219250 373600 219256 373612
rect 219308 373600 219314 373652
rect 377306 373600 377312 373652
rect 377364 373640 377370 373652
rect 455414 373640 455420 373652
rect 377364 373612 455420 373640
rect 377364 373600 377370 373612
rect 455414 373600 455420 373612
rect 455472 373600 455478 373652
rect 46198 373532 46204 373584
rect 46256 373572 46262 373584
rect 107838 373572 107844 373584
rect 46256 373544 107844 373572
rect 46256 373532 46262 373544
rect 107838 373532 107844 373544
rect 107896 373532 107902 373584
rect 124122 373532 124128 373584
rect 124180 373572 124186 373584
rect 197814 373572 197820 373584
rect 124180 373544 197820 373572
rect 124180 373532 124186 373544
rect 197814 373532 197820 373544
rect 197872 373532 197878 373584
rect 362862 373532 362868 373584
rect 362920 373572 362926 373584
rect 445846 373572 445852 373584
rect 362920 373544 445852 373572
rect 362920 373532 362926 373544
rect 445846 373532 445852 373544
rect 445904 373532 445910 373584
rect 58434 373464 58440 373516
rect 58492 373504 58498 373516
rect 125686 373504 125692 373516
rect 58492 373476 125692 373504
rect 58492 373464 58498 373476
rect 125686 373464 125692 373476
rect 125744 373464 125750 373516
rect 128906 373464 128912 373516
rect 128964 373504 128970 373516
rect 205818 373504 205824 373516
rect 128964 373476 205824 373504
rect 128964 373464 128970 373476
rect 205818 373464 205824 373476
rect 205876 373464 205882 373516
rect 209682 373464 209688 373516
rect 209740 373504 209746 373516
rect 214190 373504 214196 373516
rect 209740 373476 214196 373504
rect 209740 373464 209746 373476
rect 214190 373464 214196 373476
rect 214248 373464 214254 373516
rect 215294 373464 215300 373516
rect 215352 373504 215358 373516
rect 263686 373504 263692 373516
rect 215352 373476 263692 373504
rect 215352 373464 215358 373476
rect 263686 373464 263692 373476
rect 263744 373464 263750 373516
rect 358722 373464 358728 373516
rect 358780 373504 358786 373516
rect 447686 373504 447692 373516
rect 358780 373476 447692 373504
rect 358780 373464 358786 373476
rect 447686 373464 447692 373476
rect 447744 373464 447750 373516
rect 48774 373396 48780 373448
rect 48832 373436 48838 373448
rect 110414 373436 110420 373448
rect 48832 373408 110420 373436
rect 48832 373396 48838 373408
rect 110414 373396 110420 373408
rect 110472 373396 110478 373448
rect 121362 373396 121368 373448
rect 121420 373436 121426 373448
rect 200574 373436 200580 373448
rect 121420 373408 200580 373436
rect 121420 373396 121426 373408
rect 200574 373396 200580 373408
rect 200632 373396 200638 373448
rect 367554 373396 367560 373448
rect 367612 373436 367618 373448
rect 458174 373436 458180 373448
rect 367612 373408 458180 373436
rect 367612 373396 367618 373408
rect 458174 373396 458180 373408
rect 458232 373396 458238 373448
rect 50154 373328 50160 373380
rect 50212 373368 50218 373380
rect 98270 373368 98276 373380
rect 50212 373340 98276 373368
rect 50212 373328 50218 373340
rect 98270 373328 98276 373340
rect 98328 373328 98334 373380
rect 99374 373328 99380 373380
rect 99432 373368 99438 373380
rect 204254 373368 204260 373380
rect 99432 373340 204260 373368
rect 99432 373328 99438 373340
rect 204254 373328 204260 373340
rect 204312 373328 204318 373380
rect 262766 373328 262772 373380
rect 262824 373368 262830 373380
rect 269206 373368 269212 373380
rect 262824 373340 269212 373368
rect 262824 373328 262830 373340
rect 269206 373328 269212 373340
rect 269264 373328 269270 373380
rect 359458 373328 359464 373380
rect 359516 373368 359522 373380
rect 452838 373368 452844 373380
rect 359516 373340 452844 373368
rect 359516 373328 359522 373340
rect 452838 373328 452844 373340
rect 452896 373328 452902 373380
rect 46290 373260 46296 373312
rect 46348 373300 46354 373312
rect 93670 373300 93676 373312
rect 46348 373272 93676 373300
rect 46348 373260 46354 373272
rect 93670 373260 93676 373272
rect 93728 373260 93734 373312
rect 95050 373260 95056 373312
rect 95108 373300 95114 373312
rect 213454 373300 213460 373312
rect 95108 373272 213460 373300
rect 95108 373260 95114 373272
rect 213454 373260 213460 373272
rect 213512 373300 213518 373312
rect 219802 373300 219808 373312
rect 213512 373272 219808 373300
rect 213512 373260 213518 373272
rect 219802 373260 219808 373272
rect 219860 373300 219866 373312
rect 220722 373300 220728 373312
rect 219860 373272 220728 373300
rect 219860 373260 219866 373272
rect 220722 373260 220728 373272
rect 220780 373260 220786 373312
rect 364058 373260 364064 373312
rect 364116 373300 364122 373312
rect 485774 373300 485780 373312
rect 364116 373272 485780 373300
rect 364116 373260 364122 373272
rect 485774 373260 485780 373272
rect 485832 373260 485838 373312
rect 57054 373192 57060 373244
rect 57112 373232 57118 373244
rect 100846 373232 100852 373244
rect 57112 373204 100852 373232
rect 57112 373192 57118 373204
rect 100846 373192 100852 373204
rect 100904 373192 100910 373244
rect 151722 373192 151728 373244
rect 151780 373232 151786 373244
rect 197722 373232 197728 373244
rect 151780 373204 197728 373232
rect 151780 373192 151786 373204
rect 197722 373192 197728 373204
rect 197780 373192 197786 373244
rect 213914 373192 213920 373244
rect 213972 373232 213978 373244
rect 261294 373232 261300 373244
rect 213972 373204 261300 373232
rect 213972 373192 213978 373204
rect 261294 373192 261300 373204
rect 261352 373192 261358 373244
rect 367646 373192 367652 373244
rect 367704 373232 367710 373244
rect 376754 373232 376760 373244
rect 367704 373204 376760 373232
rect 367704 373192 367710 373204
rect 376754 373192 376760 373204
rect 376812 373192 376818 373244
rect 48866 373124 48872 373176
rect 48924 373164 48930 373176
rect 88334 373164 88340 373176
rect 48924 373136 88340 373164
rect 48924 373124 48930 373136
rect 88334 373124 88340 373136
rect 88392 373124 88398 373176
rect 154114 373124 154120 373176
rect 154172 373164 154178 373176
rect 198366 373164 198372 373176
rect 154172 373136 198372 373164
rect 154172 373124 154178 373136
rect 198366 373124 198372 373136
rect 198424 373124 198430 373176
rect 207198 373124 207204 373176
rect 207256 373164 207262 373176
rect 213546 373164 213552 373176
rect 207256 373136 213552 373164
rect 207256 373124 207262 373136
rect 213546 373124 213552 373136
rect 213604 373164 213610 373176
rect 242894 373164 242900 373176
rect 213604 373136 242900 373164
rect 213604 373124 213610 373136
rect 242894 373124 242900 373136
rect 242952 373124 242958 373176
rect 55766 373056 55772 373108
rect 55824 373096 55830 373108
rect 90174 373096 90180 373108
rect 55824 373068 90180 373096
rect 55824 373056 55830 373068
rect 90174 373056 90180 373068
rect 90232 373056 90238 373108
rect 214098 373056 214104 373108
rect 214156 373096 214162 373108
rect 217778 373096 217784 373108
rect 214156 373068 217784 373096
rect 214156 373056 214162 373068
rect 217778 373056 217784 373068
rect 217836 373056 217842 373108
rect 220722 373056 220728 373108
rect 220780 373096 220786 373108
rect 253934 373096 253940 373108
rect 220780 373068 253940 373096
rect 220780 373056 220786 373068
rect 253934 373056 253940 373068
rect 253992 373056 253998 373108
rect 212902 372988 212908 373040
rect 212960 373028 212966 373040
rect 255406 373028 255412 373040
rect 212960 373000 255412 373028
rect 212960 372988 212966 373000
rect 255406 372988 255412 373000
rect 255464 372988 255470 373040
rect 212626 372920 212632 372972
rect 212684 372960 212690 372972
rect 256694 372960 256700 372972
rect 212684 372932 256700 372960
rect 212684 372920 212690 372932
rect 256694 372920 256700 372932
rect 256752 372920 256758 372972
rect 214006 372852 214012 372904
rect 214064 372892 214070 372904
rect 214064 372864 224264 372892
rect 214064 372852 214070 372864
rect 217042 372784 217048 372836
rect 217100 372824 217106 372836
rect 217686 372824 217692 372836
rect 217100 372796 217692 372824
rect 217100 372784 217106 372796
rect 217686 372784 217692 372796
rect 217744 372784 217750 372836
rect 217778 372784 217784 372836
rect 217836 372824 217842 372836
rect 224126 372824 224132 372836
rect 217836 372796 224132 372824
rect 217836 372784 217842 372796
rect 224126 372784 224132 372796
rect 224184 372784 224190 372836
rect 224236 372824 224264 372864
rect 224310 372852 224316 372904
rect 224368 372892 224374 372904
rect 259638 372892 259644 372904
rect 224368 372864 259644 372892
rect 224368 372852 224374 372864
rect 259638 372852 259644 372864
rect 259696 372852 259702 372904
rect 259454 372824 259460 372836
rect 224236 372796 259460 372824
rect 259454 372784 259460 372796
rect 259512 372784 259518 372836
rect 210142 372716 210148 372768
rect 210200 372756 210206 372768
rect 210326 372756 210332 372768
rect 210200 372728 210332 372756
rect 210200 372716 210206 372728
rect 210326 372716 210332 372728
rect 210384 372716 210390 372768
rect 212534 372716 212540 372768
rect 212592 372756 212598 372768
rect 258074 372756 258080 372768
rect 212592 372728 258080 372756
rect 212592 372716 212598 372728
rect 258074 372716 258080 372728
rect 258132 372716 258138 372768
rect 203058 372648 203064 372700
rect 203116 372688 203122 372700
rect 216306 372688 216312 372700
rect 203116 372660 216312 372688
rect 203116 372648 203122 372660
rect 216306 372648 216312 372660
rect 216364 372688 216370 372700
rect 216364 372660 218560 372688
rect 216364 372648 216370 372660
rect 51626 372580 51632 372632
rect 51684 372620 51690 372632
rect 54386 372620 54392 372632
rect 51684 372592 54392 372620
rect 51684 372580 51690 372592
rect 54386 372580 54392 372592
rect 54444 372580 54450 372632
rect 56962 372580 56968 372632
rect 57020 372620 57026 372632
rect 58526 372620 58532 372632
rect 57020 372592 58532 372620
rect 57020 372580 57026 372592
rect 58526 372580 58532 372592
rect 58584 372580 58590 372632
rect 95970 372580 95976 372632
rect 96028 372620 96034 372632
rect 212902 372620 212908 372632
rect 96028 372592 212908 372620
rect 96028 372580 96034 372592
rect 212902 372580 212908 372592
rect 212960 372580 212966 372632
rect 215294 372580 215300 372632
rect 215352 372620 215358 372632
rect 215662 372620 215668 372632
rect 215352 372592 215668 372620
rect 215352 372580 215358 372592
rect 215662 372580 215668 372592
rect 215720 372580 215726 372632
rect 218532 372620 218560 372660
rect 219250 372648 219256 372700
rect 219308 372688 219314 372700
rect 236086 372688 236092 372700
rect 219308 372660 236092 372688
rect 219308 372648 219314 372660
rect 236086 372648 236092 372660
rect 236144 372648 236150 372700
rect 369670 372648 369676 372700
rect 369728 372688 369734 372700
rect 373718 372688 373724 372700
rect 369728 372660 373724 372688
rect 369728 372648 369734 372660
rect 373718 372648 373724 372660
rect 373776 372648 373782 372700
rect 376754 372648 376760 372700
rect 376812 372688 376818 372700
rect 378042 372688 378048 372700
rect 376812 372660 378048 372688
rect 376812 372648 376818 372660
rect 378042 372648 378048 372660
rect 378100 372688 378106 372700
rect 408494 372688 408500 372700
rect 378100 372660 408500 372688
rect 378100 372648 378106 372660
rect 408494 372648 408500 372660
rect 408552 372648 408558 372700
rect 235994 372620 236000 372632
rect 218532 372592 236000 372620
rect 235994 372580 236000 372592
rect 236052 372580 236058 372632
rect 372522 372580 372528 372632
rect 372580 372620 372586 372632
rect 373994 372620 374000 372632
rect 372580 372592 374000 372620
rect 372580 372580 372586 372592
rect 373994 372580 374000 372592
rect 374052 372620 374058 372632
rect 375190 372620 375196 372632
rect 374052 372592 375196 372620
rect 374052 372580 374058 372592
rect 375190 372580 375196 372592
rect 375248 372580 375254 372632
rect 379146 372580 379152 372632
rect 379204 372620 379210 372632
rect 379330 372620 379336 372632
rect 379204 372592 379336 372620
rect 379204 372580 379210 372592
rect 379330 372580 379336 372592
rect 379388 372620 379394 372632
rect 426434 372620 426440 372632
rect 379388 372592 426440 372620
rect 379388 372580 379394 372592
rect 426434 372580 426440 372592
rect 426492 372580 426498 372632
rect 89346 372512 89352 372564
rect 89404 372552 89410 372564
rect 209866 372552 209872 372564
rect 89404 372524 209872 372552
rect 89404 372512 89410 372524
rect 209866 372512 209872 372524
rect 209924 372552 209930 372564
rect 210326 372552 210332 372564
rect 209924 372524 210332 372552
rect 209924 372512 209930 372524
rect 210326 372512 210332 372524
rect 210384 372512 210390 372564
rect 211706 372512 211712 372564
rect 211764 372552 211770 372564
rect 213730 372552 213736 372564
rect 211764 372524 213736 372552
rect 211764 372512 211770 372524
rect 213730 372512 213736 372524
rect 213788 372512 213794 372564
rect 214466 372512 214472 372564
rect 214524 372552 214530 372564
rect 219526 372552 219532 372564
rect 214524 372524 219532 372552
rect 214524 372512 214530 372524
rect 219526 372512 219532 372524
rect 219584 372552 219590 372564
rect 273254 372552 273260 372564
rect 219584 372524 273260 372552
rect 219584 372512 219590 372524
rect 273254 372512 273260 372524
rect 273312 372512 273318 372564
rect 304994 372512 305000 372564
rect 305052 372552 305058 372564
rect 313274 372552 313280 372564
rect 305052 372524 313280 372552
rect 305052 372512 305058 372524
rect 313274 372512 313280 372524
rect 313332 372512 313338 372564
rect 369854 372512 369860 372564
rect 369912 372552 369918 372564
rect 437474 372552 437480 372564
rect 369912 372524 437480 372552
rect 369912 372512 369918 372524
rect 437474 372512 437480 372524
rect 437532 372512 437538 372564
rect 92382 372444 92388 372496
rect 92440 372484 92446 372496
rect 92440 372456 209774 372484
rect 92440 372444 92446 372456
rect 90082 372376 90088 372428
rect 90140 372416 90146 372428
rect 90140 372388 200114 372416
rect 90140 372376 90146 372388
rect 77202 372308 77208 372360
rect 77260 372348 77266 372360
rect 99374 372348 99380 372360
rect 77260 372320 99380 372348
rect 77260 372308 77266 372320
rect 99374 372308 99380 372320
rect 99432 372308 99438 372360
rect 200086 372280 200114 372388
rect 209746 372348 209774 372456
rect 304258 372444 304264 372496
rect 304316 372484 304322 372496
rect 310514 372484 310520 372496
rect 304316 372456 310520 372484
rect 304316 372444 304322 372456
rect 310514 372444 310520 372456
rect 310572 372444 310578 372496
rect 375190 372444 375196 372496
rect 375248 372484 375254 372496
rect 433334 372484 433340 372496
rect 375248 372456 433340 372484
rect 375248 372444 375254 372456
rect 433334 372444 433340 372456
rect 433392 372444 433398 372496
rect 220722 372376 220728 372428
rect 220780 372416 220786 372428
rect 248414 372416 248420 372428
rect 220780 372388 248420 372416
rect 220780 372376 220786 372388
rect 248414 372376 248420 372388
rect 248472 372376 248478 372428
rect 211154 372348 211160 372360
rect 209746 372320 211160 372348
rect 211154 372308 211160 372320
rect 211212 372348 211218 372360
rect 220998 372348 221004 372360
rect 211212 372320 221004 372348
rect 211212 372308 211218 372320
rect 220998 372308 221004 372320
rect 221056 372348 221062 372360
rect 221918 372348 221924 372360
rect 221056 372320 221924 372348
rect 221056 372308 221062 372320
rect 221918 372308 221924 372320
rect 221976 372308 221982 372360
rect 209774 372280 209780 372292
rect 200086 372252 209780 372280
rect 209774 372240 209780 372252
rect 209832 372280 209838 372292
rect 220078 372280 220084 372292
rect 209832 372252 220084 372280
rect 209832 372240 209838 372252
rect 220078 372240 220084 372252
rect 220136 372240 220142 372292
rect 221550 372172 221556 372224
rect 221608 372212 221614 372224
rect 240870 372212 240876 372224
rect 221608 372184 240876 372212
rect 221608 372172 221614 372184
rect 240870 372172 240876 372184
rect 240928 372172 240934 372224
rect 86586 372104 86592 372156
rect 86644 372144 86650 372156
rect 210142 372144 210148 372156
rect 86644 372116 210148 372144
rect 86644 372104 86650 372116
rect 210142 372104 210148 372116
rect 210200 372144 210206 372156
rect 215754 372144 215760 372156
rect 210200 372116 215760 372144
rect 210200 372104 210206 372116
rect 215754 372104 215760 372116
rect 215812 372144 215818 372156
rect 245654 372144 245660 372156
rect 215812 372116 245660 372144
rect 215812 372104 215818 372116
rect 245654 372104 245660 372116
rect 245712 372104 245718 372156
rect 210326 372036 210332 372088
rect 210384 372076 210390 372088
rect 219526 372076 219532 372088
rect 210384 372048 219532 372076
rect 210384 372036 210390 372048
rect 219526 372036 219532 372048
rect 219584 372076 219590 372088
rect 220722 372076 220728 372088
rect 219584 372048 220728 372076
rect 219584 372036 219590 372048
rect 220722 372036 220728 372048
rect 220780 372036 220786 372088
rect 251174 372076 251180 372088
rect 221568 372048 251180 372076
rect 47670 371968 47676 372020
rect 47728 372008 47734 372020
rect 78490 372008 78496 372020
rect 47728 371980 78496 372008
rect 47728 371968 47734 371980
rect 78490 371968 78496 371980
rect 78548 371968 78554 372020
rect 213454 371968 213460 372020
rect 213512 372008 213518 372020
rect 219618 372008 219624 372020
rect 213512 371980 219624 372008
rect 213512 371968 213518 371980
rect 219618 371968 219624 371980
rect 219676 372008 219682 372020
rect 221568 372008 221596 372048
rect 251174 372036 251180 372048
rect 251232 372036 251238 372088
rect 368382 372036 368388 372088
rect 368440 372076 368446 372088
rect 376754 372076 376760 372088
rect 368440 372048 376760 372076
rect 368440 372036 368446 372048
rect 376754 372036 376760 372048
rect 376812 372036 376818 372088
rect 219676 371980 221596 372008
rect 219676 371968 219682 371980
rect 221642 371968 221648 372020
rect 221700 372008 221706 372020
rect 240778 372008 240784 372020
rect 221700 371980 240784 372008
rect 221700 371968 221706 371980
rect 240778 371968 240784 371980
rect 240836 371968 240842 372020
rect 357250 371968 357256 372020
rect 357308 372008 357314 372020
rect 379514 372008 379520 372020
rect 357308 371980 379520 372008
rect 357308 371968 357314 371980
rect 379514 371968 379520 371980
rect 379572 371968 379578 372020
rect 379974 371968 379980 372020
rect 380032 372008 380038 372020
rect 396074 372008 396080 372020
rect 380032 371980 396080 372008
rect 380032 371968 380038 371980
rect 396074 371968 396080 371980
rect 396132 371968 396138 372020
rect 44726 371900 44732 371952
rect 44784 371940 44790 371952
rect 48866 371940 48872 371952
rect 44784 371912 48872 371940
rect 44784 371900 44790 371912
rect 48866 371900 48872 371912
rect 48924 371900 48930 371952
rect 108850 371900 108856 371952
rect 108908 371940 108914 371952
rect 204162 371940 204168 371952
rect 108908 371912 204168 371940
rect 108908 371900 108914 371912
rect 204162 371900 204168 371912
rect 204220 371940 204226 371952
rect 217042 371940 217048 371952
rect 204220 371912 217048 371940
rect 204220 371900 204226 371912
rect 217042 371900 217048 371912
rect 217100 371940 217106 371952
rect 262858 371940 262864 371952
rect 217100 371912 262864 371940
rect 217100 371900 217106 371912
rect 262858 371900 262864 371912
rect 262916 371900 262922 371952
rect 360746 371900 360752 371952
rect 360804 371940 360810 371952
rect 376478 371940 376484 371952
rect 360804 371912 376484 371940
rect 360804 371900 360810 371912
rect 376478 371900 376484 371912
rect 376536 371900 376542 371952
rect 379422 371900 379428 371952
rect 379480 371940 379486 371952
rect 404354 371940 404360 371952
rect 379480 371912 404360 371940
rect 379480 371900 379486 371912
rect 404354 371900 404360 371912
rect 404412 371900 404418 371952
rect 47578 371832 47584 371884
rect 47636 371872 47642 371884
rect 79962 371872 79968 371884
rect 47636 371844 79968 371872
rect 47636 371832 47642 371844
rect 79962 371832 79968 371844
rect 80020 371832 80026 371884
rect 85482 371832 85488 371884
rect 85540 371872 85546 371884
rect 106182 371872 106188 371884
rect 85540 371844 106188 371872
rect 85540 371832 85546 371844
rect 106182 371832 106188 371844
rect 106240 371832 106246 371884
rect 114002 371832 114008 371884
rect 114060 371872 114066 371884
rect 214466 371872 214472 371884
rect 114060 371844 214472 371872
rect 114060 371832 114066 371844
rect 214466 371832 214472 371844
rect 214524 371872 214530 371884
rect 215018 371872 215024 371884
rect 214524 371844 215024 371872
rect 214524 371832 214530 371844
rect 215018 371832 215024 371844
rect 215076 371832 215082 371884
rect 220906 371872 220912 371884
rect 219406 371844 220912 371872
rect 88058 371764 88064 371816
rect 88116 371804 88122 371816
rect 211706 371804 211712 371816
rect 88116 371776 211712 371804
rect 88116 371764 88122 371776
rect 211706 371764 211712 371776
rect 211764 371764 211770 371816
rect 93578 371696 93584 371748
rect 93636 371736 93642 371748
rect 219406 371736 219434 371844
rect 220906 371832 220912 371844
rect 220964 371872 220970 371884
rect 250622 371872 250628 371884
rect 220964 371844 250628 371872
rect 220964 371832 220970 371844
rect 250622 371832 250628 371844
rect 250680 371832 250686 371884
rect 275370 371832 275376 371884
rect 275428 371872 275434 371884
rect 356974 371872 356980 371884
rect 275428 371844 356980 371872
rect 275428 371832 275434 371844
rect 356974 371832 356980 371844
rect 357032 371832 357038 371884
rect 375190 371832 375196 371884
rect 375248 371872 375254 371884
rect 400214 371872 400220 371884
rect 375248 371844 400220 371872
rect 375248 371832 375254 371844
rect 400214 371832 400220 371844
rect 400272 371832 400278 371884
rect 517882 371832 517888 371884
rect 517940 371872 517946 371884
rect 580442 371872 580448 371884
rect 517940 371844 580448 371872
rect 517940 371832 517946 371844
rect 580442 371832 580448 371844
rect 580500 371832 580506 371884
rect 222102 371764 222108 371816
rect 222160 371804 222166 371816
rect 241514 371804 241520 371816
rect 222160 371776 241520 371804
rect 222160 371764 222166 371776
rect 241514 371764 241520 371776
rect 241572 371804 241578 371816
rect 241572 371776 248414 371804
rect 241572 371764 241578 371776
rect 93636 371708 219434 371736
rect 93636 371696 93642 371708
rect 92198 371628 92204 371680
rect 92256 371668 92262 371680
rect 211246 371668 211252 371680
rect 92256 371640 211252 371668
rect 92256 371628 92262 371640
rect 211246 371628 211252 371640
rect 211304 371668 211310 371680
rect 213454 371668 213460 371680
rect 211304 371640 213460 371668
rect 211304 371628 211310 371640
rect 213454 371628 213460 371640
rect 213512 371628 213518 371680
rect 215294 371560 215300 371612
rect 215352 371600 215358 371612
rect 215570 371600 215576 371612
rect 215352 371572 215576 371600
rect 215352 371560 215358 371572
rect 215570 371560 215576 371572
rect 215628 371600 215634 371612
rect 240410 371600 240416 371612
rect 215628 371572 240416 371600
rect 215628 371560 215634 371572
rect 240410 371560 240416 371572
rect 240468 371600 240474 371612
rect 241422 371600 241428 371612
rect 240468 371572 241428 371600
rect 240468 371560 240474 371572
rect 241422 371560 241428 371572
rect 241480 371560 241486 371612
rect 248386 371600 248414 371776
rect 276290 371764 276296 371816
rect 276348 371804 276354 371816
rect 357250 371804 357256 371816
rect 276348 371776 357256 371804
rect 276348 371764 276354 371776
rect 357250 371764 357256 371776
rect 357308 371764 357314 371816
rect 372982 371764 372988 371816
rect 373040 371804 373046 371816
rect 398834 371804 398840 371816
rect 373040 371776 398840 371804
rect 373040 371764 373046 371776
rect 398834 371764 398840 371776
rect 398892 371764 398898 371816
rect 273254 371696 273260 371748
rect 273312 371736 273318 371748
rect 304994 371736 305000 371748
rect 273312 371708 305000 371736
rect 273312 371696 273318 371708
rect 304994 371696 305000 371708
rect 305052 371696 305058 371748
rect 371050 371696 371056 371748
rect 371108 371736 371114 371748
rect 397454 371736 397460 371748
rect 371108 371708 397460 371736
rect 371108 371696 371114 371708
rect 397454 371696 397460 371708
rect 397512 371696 397518 371748
rect 278682 371628 278688 371680
rect 278740 371668 278746 371680
rect 357434 371668 357440 371680
rect 278740 371640 357440 371668
rect 278740 371628 278746 371640
rect 357434 371628 357440 371640
rect 357492 371628 357498 371680
rect 379514 371628 379520 371680
rect 379572 371668 379578 371680
rect 379882 371668 379888 371680
rect 379572 371640 379888 371668
rect 379572 371628 379578 371640
rect 379882 371628 379888 371640
rect 379940 371668 379946 371680
rect 409874 371668 409880 371680
rect 379940 371640 409880 371668
rect 379940 371628 379946 371640
rect 409874 371628 409880 371640
rect 409932 371628 409938 371680
rect 371142 371600 371148 371612
rect 248386 371572 371148 371600
rect 371142 371560 371148 371572
rect 371200 371600 371206 371612
rect 371200 371572 373488 371600
rect 371200 371560 371206 371572
rect 48866 371492 48872 371544
rect 48924 371532 48930 371544
rect 81894 371532 81900 371544
rect 48924 371504 81900 371532
rect 48924 371492 48930 371504
rect 81894 371492 81900 371504
rect 81952 371532 81958 371544
rect 82446 371532 82452 371544
rect 81952 371504 82452 371532
rect 81952 371492 81958 371504
rect 82446 371492 82452 371504
rect 82504 371492 82510 371544
rect 85114 371492 85120 371544
rect 85172 371532 85178 371544
rect 210234 371532 210240 371544
rect 85172 371504 210240 371532
rect 85172 371492 85178 371504
rect 210234 371492 210240 371504
rect 210292 371532 210298 371544
rect 215110 371532 215116 371544
rect 210292 371504 215116 371532
rect 210292 371492 210298 371504
rect 215110 371492 215116 371504
rect 215168 371492 215174 371544
rect 221918 371492 221924 371544
rect 221976 371532 221982 371544
rect 223114 371532 223120 371544
rect 221976 371504 223120 371532
rect 221976 371492 221982 371504
rect 223114 371492 223120 371504
rect 223172 371492 223178 371544
rect 237374 371492 237380 371544
rect 237432 371532 237438 371544
rect 238110 371532 238116 371544
rect 237432 371504 238116 371532
rect 237432 371492 237438 371504
rect 238110 371492 238116 371504
rect 238168 371532 238174 371544
rect 371050 371532 371056 371544
rect 238168 371504 371056 371532
rect 238168 371492 238174 371504
rect 371050 371492 371056 371504
rect 371108 371492 371114 371544
rect 373460 371532 373488 371572
rect 376570 371560 376576 371612
rect 376628 371600 376634 371612
rect 380986 371600 380992 371612
rect 376628 371572 380992 371600
rect 376628 371560 376634 371572
rect 380986 371560 380992 371572
rect 381044 371600 381050 371612
rect 411254 371600 411260 371612
rect 381044 371572 411260 371600
rect 381044 371560 381050 371572
rect 411254 371560 411260 371572
rect 411312 371560 411318 371612
rect 401594 371532 401600 371544
rect 373460 371504 401600 371532
rect 401594 371492 401600 371504
rect 401652 371492 401658 371544
rect 79962 371424 79968 371476
rect 80020 371464 80026 371476
rect 209590 371464 209596 371476
rect 80020 371436 209596 371464
rect 80020 371424 80026 371436
rect 209590 371424 209596 371436
rect 209648 371464 209654 371476
rect 239306 371464 239312 371476
rect 209648 371436 239312 371464
rect 209648 371424 209654 371436
rect 239306 371424 239312 371436
rect 239364 371464 239370 371476
rect 372982 371464 372988 371476
rect 239364 371436 372988 371464
rect 239364 371424 239370 371436
rect 372982 371424 372988 371436
rect 373040 371424 373046 371476
rect 376478 371424 376484 371476
rect 376536 371464 376542 371476
rect 407114 371464 407120 371476
rect 376536 371436 407120 371464
rect 376536 371424 376542 371436
rect 407114 371424 407120 371436
rect 407172 371424 407178 371476
rect 78490 371356 78496 371408
rect 78548 371396 78554 371408
rect 208210 371396 208216 371408
rect 78548 371368 208216 371396
rect 78548 371356 78554 371368
rect 208210 371356 208216 371368
rect 208268 371396 208274 371408
rect 237374 371396 237380 371408
rect 208268 371368 237380 371396
rect 208268 371356 208274 371368
rect 237374 371356 237380 371368
rect 237432 371356 237438 371408
rect 241422 371356 241428 371408
rect 241480 371396 241486 371408
rect 375190 371396 375196 371408
rect 241480 371368 375196 371396
rect 241480 371356 241486 371368
rect 375190 371356 375196 371368
rect 375248 371356 375254 371408
rect 376754 371356 376760 371408
rect 376812 371396 376818 371408
rect 377950 371396 377956 371408
rect 376812 371368 377956 371396
rect 376812 371356 376818 371368
rect 377950 371356 377956 371368
rect 378008 371396 378014 371408
rect 411254 371396 411260 371408
rect 378008 371368 411260 371396
rect 378008 371356 378014 371368
rect 411254 371356 411260 371368
rect 411312 371356 411318 371408
rect 439866 371356 439872 371408
rect 439924 371396 439930 371408
rect 516594 371396 516600 371408
rect 439924 371368 516600 371396
rect 439924 371356 439930 371368
rect 516594 371356 516600 371368
rect 516652 371356 516658 371408
rect 80514 371328 80520 371340
rect 64846 371300 80520 371328
rect 44818 371220 44824 371272
rect 44876 371260 44882 371272
rect 46290 371260 46296 371272
rect 44876 371232 46296 371260
rect 44876 371220 44882 371232
rect 46290 371220 46296 371232
rect 46348 371260 46354 371272
rect 64846 371260 64874 371300
rect 80514 371288 80520 371300
rect 80572 371328 80578 371340
rect 215294 371328 215300 371340
rect 80572 371300 215300 371328
rect 80572 371288 80578 371300
rect 215294 371288 215300 371300
rect 215352 371288 215358 371340
rect 219894 371288 219900 371340
rect 219952 371328 219958 371340
rect 220078 371328 220084 371340
rect 219952 371300 220084 371328
rect 219952 371288 219958 371300
rect 220078 371288 220084 371300
rect 220136 371328 220142 371340
rect 249794 371328 249800 371340
rect 220136 371300 249800 371328
rect 220136 371288 220142 371300
rect 249794 371288 249800 371300
rect 249852 371288 249858 371340
rect 342898 371288 342904 371340
rect 342956 371328 342962 371340
rect 343450 371328 343456 371340
rect 342956 371300 343456 371328
rect 342956 371288 342962 371300
rect 343450 371288 343456 371300
rect 343508 371328 343514 371340
rect 363046 371328 363052 371340
rect 343508 371300 363052 371328
rect 343508 371288 343514 371300
rect 363046 371288 363052 371300
rect 363104 371328 363110 371340
rect 503530 371328 503536 371340
rect 363104 371300 503536 371328
rect 363104 371288 363110 371300
rect 503530 371288 503536 371300
rect 503588 371328 503594 371340
rect 517882 371328 517888 371340
rect 503588 371300 517888 371328
rect 503588 371288 503594 371300
rect 517882 371288 517888 371300
rect 517940 371288 517946 371340
rect 46348 371232 64874 371260
rect 46348 371220 46354 371232
rect 82446 371220 82452 371272
rect 82504 371260 82510 371272
rect 220814 371260 220820 371272
rect 82504 371232 220820 371260
rect 82504 371220 82510 371232
rect 220814 371220 220820 371232
rect 220872 371260 220878 371272
rect 222102 371260 222108 371272
rect 220872 371232 222108 371260
rect 220872 371220 220878 371232
rect 222102 371220 222108 371232
rect 222160 371220 222166 371272
rect 223114 371220 223120 371272
rect 223172 371260 223178 371272
rect 251174 371260 251180 371272
rect 223172 371232 251180 371260
rect 223172 371220 223178 371232
rect 251174 371220 251180 371232
rect 251232 371220 251238 371272
rect 343082 371220 343088 371272
rect 343140 371260 343146 371272
rect 360194 371260 360200 371272
rect 343140 371232 360200 371260
rect 343140 371220 343146 371232
rect 360194 371220 360200 371232
rect 360252 371260 360258 371272
rect 503162 371260 503168 371272
rect 360252 371232 503168 371260
rect 360252 371220 360258 371232
rect 503162 371220 503168 371232
rect 503220 371260 503226 371272
rect 517790 371260 517796 371272
rect 503220 371232 517796 371260
rect 503220 371220 503226 371232
rect 517790 371220 517796 371232
rect 517848 371260 517854 371272
rect 580258 371260 580264 371272
rect 517848 371232 580264 371260
rect 517848 371220 517854 371232
rect 580258 371220 580264 371232
rect 580316 371220 580322 371272
rect 43346 371152 43352 371204
rect 43404 371192 43410 371204
rect 183186 371192 183192 371204
rect 43404 371164 183192 371192
rect 43404 371152 43410 371164
rect 183186 371152 183192 371164
rect 183244 371192 183250 371204
rect 201034 371192 201040 371204
rect 183244 371164 201040 371192
rect 183244 371152 183250 371164
rect 201034 371152 201040 371164
rect 201092 371152 201098 371204
rect 201494 371152 201500 371204
rect 201552 371192 201558 371204
rect 317414 371192 317420 371204
rect 201552 371164 317420 371192
rect 201552 371152 201558 371164
rect 317414 371152 317420 371164
rect 317472 371152 317478 371204
rect 375098 371152 375104 371204
rect 375156 371192 375162 371204
rect 376570 371192 376576 371204
rect 375156 371164 376576 371192
rect 375156 371152 375162 371164
rect 376570 371152 376576 371164
rect 376628 371152 376634 371204
rect 376754 371152 376760 371204
rect 376812 371192 376818 371204
rect 402974 371192 402980 371204
rect 376812 371164 402980 371192
rect 376812 371152 376818 371164
rect 402974 371152 402980 371164
rect 403032 371152 403038 371204
rect 54570 371084 54576 371136
rect 54628 371124 54634 371136
rect 182818 371124 182824 371136
rect 54628 371096 182824 371124
rect 54628 371084 54634 371096
rect 182818 371084 182824 371096
rect 182876 371084 182882 371136
rect 198826 371084 198832 371136
rect 198884 371124 198890 371136
rect 302234 371124 302240 371136
rect 198884 371096 302240 371124
rect 198884 371084 198890 371096
rect 302234 371084 302240 371096
rect 302292 371084 302298 371136
rect 357986 371084 357992 371136
rect 358044 371124 358050 371136
rect 473354 371124 473360 371136
rect 358044 371096 473360 371124
rect 358044 371084 358050 371096
rect 473354 371084 473360 371096
rect 473412 371084 473418 371136
rect 197354 371016 197360 371068
rect 197412 371056 197418 371068
rect 295334 371056 295340 371068
rect 197412 371028 295340 371056
rect 197412 371016 197418 371028
rect 295334 371016 295340 371028
rect 295392 371016 295398 371068
rect 357158 371016 357164 371068
rect 357216 371056 357222 371068
rect 465074 371056 465080 371068
rect 357216 371028 465080 371056
rect 357216 371016 357222 371028
rect 465074 371016 465080 371028
rect 465132 371016 465138 371068
rect 102778 370948 102784 371000
rect 102836 370988 102842 371000
rect 215478 370988 215484 371000
rect 102836 370960 215484 370988
rect 102836 370948 102842 370960
rect 215478 370948 215484 370960
rect 215536 370948 215542 371000
rect 217502 370948 217508 371000
rect 217560 370988 217566 371000
rect 307754 370988 307760 371000
rect 217560 370960 307760 370988
rect 217560 370948 217566 370960
rect 307754 370948 307760 370960
rect 307812 370948 307818 371000
rect 366174 370948 366180 371000
rect 366232 370988 366238 371000
rect 467834 370988 467840 371000
rect 366232 370960 467840 370988
rect 366232 370948 366238 370960
rect 467834 370948 467840 370960
rect 467892 370948 467898 371000
rect 198918 370880 198924 370932
rect 198976 370920 198982 370932
rect 300854 370920 300860 370932
rect 198976 370892 300860 370920
rect 198976 370880 198982 370892
rect 300854 370880 300860 370892
rect 300912 370880 300918 370932
rect 368934 370880 368940 370932
rect 368992 370920 368998 370932
rect 470594 370920 470600 370932
rect 368992 370892 470600 370920
rect 368992 370880 368998 370892
rect 470594 370880 470600 370892
rect 470652 370880 470658 370932
rect 197446 370812 197452 370864
rect 197504 370852 197510 370864
rect 292574 370852 292580 370864
rect 197504 370824 292580 370852
rect 197504 370812 197510 370824
rect 292574 370812 292580 370824
rect 292632 370812 292638 370864
rect 361482 370812 361488 370864
rect 361540 370852 361546 370864
rect 462314 370852 462320 370864
rect 361540 370824 462320 370852
rect 361540 370812 361546 370824
rect 462314 370812 462320 370824
rect 462372 370812 462378 370864
rect 196710 370744 196716 370796
rect 196768 370784 196774 370796
rect 289814 370784 289820 370796
rect 196768 370756 289820 370784
rect 196768 370744 196774 370756
rect 289814 370744 289820 370756
rect 289872 370744 289878 370796
rect 364886 370744 364892 370796
rect 364944 370784 364950 370796
rect 460934 370784 460940 370796
rect 364944 370756 460940 370784
rect 364944 370744 364950 370756
rect 460934 370744 460940 370756
rect 460992 370744 460998 370796
rect 196802 370676 196808 370728
rect 196860 370716 196866 370728
rect 287238 370716 287244 370728
rect 196860 370688 287244 370716
rect 196860 370676 196866 370688
rect 287238 370676 287244 370688
rect 287296 370676 287302 370728
rect 359550 370676 359556 370728
rect 359608 370716 359614 370728
rect 413186 370716 413192 370728
rect 359608 370688 413192 370716
rect 359608 370676 359614 370688
rect 413186 370676 413192 370688
rect 413244 370676 413250 370728
rect 196618 370608 196624 370660
rect 196676 370648 196682 370660
rect 285674 370648 285680 370660
rect 196676 370620 285680 370648
rect 196676 370608 196682 370620
rect 285674 370608 285680 370620
rect 285732 370608 285738 370660
rect 373810 370608 373816 370660
rect 373868 370648 373874 370660
rect 375926 370648 375932 370660
rect 373868 370620 375932 370648
rect 373868 370608 373874 370620
rect 375926 370608 375932 370620
rect 375984 370648 375990 370660
rect 376754 370648 376760 370660
rect 375984 370620 376760 370648
rect 375984 370608 375990 370620
rect 376754 370608 376760 370620
rect 376812 370608 376818 370660
rect 379238 370608 379244 370660
rect 379296 370648 379302 370660
rect 415394 370648 415400 370660
rect 379296 370620 415400 370648
rect 379296 370608 379302 370620
rect 415394 370608 415400 370620
rect 415452 370608 415458 370660
rect 199378 370540 199384 370592
rect 199436 370580 199442 370592
rect 280154 370580 280160 370592
rect 199436 370552 280160 370580
rect 199436 370540 199442 370552
rect 280154 370540 280160 370552
rect 280212 370540 280218 370592
rect 369026 370540 369032 370592
rect 369084 370580 369090 370592
rect 373994 370580 374000 370592
rect 369084 370552 374000 370580
rect 369084 370540 369090 370552
rect 373994 370540 374000 370552
rect 374052 370580 374058 370592
rect 422294 370580 422300 370592
rect 374052 370552 422300 370580
rect 374052 370540 374058 370552
rect 422294 370540 422300 370552
rect 422352 370540 422358 370592
rect 102042 370472 102048 370524
rect 102100 370512 102106 370524
rect 209498 370512 209504 370524
rect 102100 370484 209504 370512
rect 102100 370472 102106 370484
rect 209498 370472 209504 370484
rect 209556 370512 209562 370524
rect 213914 370512 213920 370524
rect 209556 370484 213920 370512
rect 209556 370472 209562 370484
rect 213914 370472 213920 370484
rect 213972 370472 213978 370524
rect 217410 370472 217416 370524
rect 217468 370512 217474 370524
rect 298094 370512 298100 370524
rect 217468 370484 298100 370512
rect 217468 370472 217474 370484
rect 298094 370472 298100 370484
rect 298152 370472 298158 370524
rect 360010 370472 360016 370524
rect 360068 370512 360074 370524
rect 518986 370512 518992 370524
rect 360068 370484 518992 370512
rect 360068 370472 360074 370484
rect 518986 370472 518992 370484
rect 519044 370472 519050 370524
rect 196986 370404 196992 370456
rect 197044 370444 197050 370456
rect 277762 370444 277768 370456
rect 197044 370416 277768 370444
rect 197044 370404 197050 370416
rect 277762 370404 277768 370416
rect 277820 370404 277826 370456
rect 376662 370404 376668 370456
rect 376720 370444 376726 370456
rect 379790 370444 379796 370456
rect 376720 370416 379796 370444
rect 376720 370404 376726 370416
rect 379790 370404 379796 370416
rect 379848 370444 379854 370456
rect 414014 370444 414020 370456
rect 379848 370416 414020 370444
rect 379848 370404 379854 370416
rect 414014 370404 414020 370416
rect 414072 370404 414078 370456
rect 198734 370336 198740 370388
rect 198792 370376 198798 370388
rect 273254 370376 273260 370388
rect 198792 370348 273260 370376
rect 198792 370336 198798 370348
rect 273254 370336 273260 370348
rect 273312 370336 273318 370388
rect 376570 370336 376576 370388
rect 376628 370376 376634 370388
rect 396074 370376 396080 370388
rect 376628 370348 396080 370376
rect 376628 370336 376634 370348
rect 396074 370336 396080 370348
rect 396132 370336 396138 370388
rect 77018 370268 77024 370320
rect 77076 370308 77082 370320
rect 203058 370308 203064 370320
rect 77076 370280 203064 370308
rect 77076 370268 77082 370280
rect 203058 370268 203064 370280
rect 203116 370268 203122 370320
rect 212902 370268 212908 370320
rect 212960 370308 212966 370320
rect 213454 370308 213460 370320
rect 212960 370280 213460 370308
rect 212960 370268 212966 370280
rect 213454 370268 213460 370280
rect 213512 370268 213518 370320
rect 215662 370268 215668 370320
rect 215720 370308 215726 370320
rect 217134 370308 217140 370320
rect 215720 370280 217140 370308
rect 215720 370268 215726 370280
rect 217134 370268 217140 370280
rect 217192 370268 217198 370320
rect 362126 370268 362132 370320
rect 362184 370308 362190 370320
rect 483014 370308 483020 370320
rect 362184 370280 483020 370308
rect 362184 370268 362190 370280
rect 483014 370268 483020 370280
rect 483072 370268 483078 370320
rect 359458 369860 359464 369912
rect 359516 369900 359522 369912
rect 360010 369900 360016 369912
rect 359516 369872 360016 369900
rect 359516 369860 359522 369872
rect 360010 369860 360016 369872
rect 360068 369860 360074 369912
rect 83826 369792 83832 369844
rect 83884 369832 83890 369844
rect 207198 369832 207204 369844
rect 83884 369804 207204 369832
rect 83884 369792 83890 369804
rect 207198 369792 207204 369804
rect 207256 369792 207262 369844
rect 216398 369792 216404 369844
rect 216456 369832 216462 369844
rect 247034 369832 247040 369844
rect 216456 369804 247040 369832
rect 216456 369792 216462 369804
rect 247034 369792 247040 369804
rect 247092 369792 247098 369844
rect 373902 369792 373908 369844
rect 373960 369832 373966 369844
rect 376938 369832 376944 369844
rect 373960 369804 376944 369832
rect 373960 369792 373966 369804
rect 376938 369792 376944 369804
rect 376996 369832 377002 369844
rect 378042 369832 378048 369844
rect 376996 369804 378048 369832
rect 376996 369792 377002 369804
rect 378042 369792 378048 369804
rect 378100 369792 378106 369844
rect 202874 369724 202880 369776
rect 202932 369764 202938 369776
rect 325878 369764 325884 369776
rect 202932 369736 325884 369764
rect 202932 369724 202938 369736
rect 325878 369724 325884 369736
rect 325936 369724 325942 369776
rect 374454 369724 374460 369776
rect 374512 369764 374518 369776
rect 477494 369764 477500 369776
rect 374512 369736 477500 369764
rect 374512 369724 374518 369736
rect 477494 369724 477500 369736
rect 477552 369724 477558 369776
rect 202966 369656 202972 369708
rect 203024 369696 203030 369708
rect 322934 369696 322940 369708
rect 203024 369668 322940 369696
rect 203024 369656 203030 369668
rect 322934 369656 322940 369668
rect 322992 369656 322998 369708
rect 356882 369656 356888 369708
rect 356940 369696 356946 369708
rect 418154 369696 418160 369708
rect 356940 369668 418160 369696
rect 356940 369656 356946 369668
rect 418154 369656 418160 369668
rect 418212 369656 418218 369708
rect 205358 369588 205364 369640
rect 205416 369628 205422 369640
rect 264974 369628 264980 369640
rect 205416 369600 264980 369628
rect 205416 369588 205422 369600
rect 264974 369588 264980 369600
rect 265032 369588 265038 369640
rect 373166 369588 373172 369640
rect 373224 369628 373230 369640
rect 427814 369628 427820 369640
rect 373224 369600 427820 369628
rect 373224 369588 373230 369600
rect 427814 369588 427820 369600
rect 427872 369588 427878 369640
rect 54570 369520 54576 369572
rect 54628 369560 54634 369572
rect 56502 369560 56508 369572
rect 54628 369532 56508 369560
rect 54628 369520 54634 369532
rect 56502 369520 56508 369532
rect 56560 369520 56566 369572
rect 211522 369520 211528 369572
rect 211580 369560 211586 369572
rect 267734 369560 267740 369572
rect 211580 369532 267740 369560
rect 211580 369520 211586 369532
rect 267734 369520 267740 369532
rect 267792 369520 267798 369572
rect 370406 369520 370412 369572
rect 370464 369560 370470 369572
rect 370464 369532 373994 369560
rect 370464 369520 370470 369532
rect 202414 369452 202420 369504
rect 202472 369492 202478 369504
rect 263594 369492 263600 369504
rect 202472 369464 263600 369492
rect 202472 369452 202478 369464
rect 263594 369452 263600 369464
rect 263652 369452 263658 369504
rect 201126 369384 201132 369436
rect 201184 369424 201190 369436
rect 260834 369424 260840 369436
rect 201184 369396 260840 369424
rect 201184 369384 201190 369396
rect 260834 369384 260840 369396
rect 260892 369384 260898 369436
rect 373966 369424 373994 369532
rect 378594 369520 378600 369572
rect 378652 369560 378658 369572
rect 425054 369560 425060 369572
rect 378652 369532 425060 369560
rect 378652 369520 378658 369532
rect 425054 369520 425060 369532
rect 425112 369520 425118 369572
rect 378042 369452 378048 369504
rect 378100 369492 378106 369504
rect 423674 369492 423680 369504
rect 378100 369464 423680 369492
rect 378100 369452 378106 369464
rect 423674 369452 423680 369464
rect 423732 369452 423738 369504
rect 374546 369424 374552 369436
rect 373966 369396 374552 369424
rect 374546 369384 374552 369396
rect 374604 369424 374610 369436
rect 416774 369424 416780 369436
rect 374604 369396 416780 369424
rect 374604 369384 374610 369396
rect 416774 369384 416780 369396
rect 416832 369384 416838 369436
rect 203886 369316 203892 369368
rect 203944 369356 203950 369368
rect 258166 369356 258172 369368
rect 203944 369328 258172 369356
rect 203944 369316 203950 369328
rect 258166 369316 258172 369328
rect 258224 369316 258230 369368
rect 371694 369316 371700 369368
rect 371752 369356 371758 369368
rect 375926 369356 375932 369368
rect 371752 369328 375932 369356
rect 371752 369316 371758 369328
rect 375926 369316 375932 369328
rect 375984 369356 375990 369368
rect 418246 369356 418252 369368
rect 375984 369328 418252 369356
rect 375984 369316 375990 369328
rect 418246 369316 418252 369328
rect 418304 369316 418310 369368
rect 100110 369248 100116 369300
rect 100168 369288 100174 369300
rect 214006 369288 214012 369300
rect 100168 369260 214012 369288
rect 100168 369248 100174 369260
rect 214006 369248 214012 369260
rect 214064 369288 214070 369300
rect 214374 369288 214380 369300
rect 214064 369260 214380 369288
rect 214064 369248 214070 369260
rect 214374 369248 214380 369260
rect 214432 369248 214438 369300
rect 219158 369248 219164 369300
rect 219216 369288 219222 369300
rect 273346 369288 273352 369300
rect 219216 369260 273352 369288
rect 219216 369248 219222 369260
rect 273346 369248 273352 369260
rect 273404 369248 273410 369300
rect 365622 369248 365628 369300
rect 365680 369288 365686 369300
rect 377122 369288 377128 369300
rect 365680 369260 377128 369288
rect 365680 369248 365686 369260
rect 377122 369248 377128 369260
rect 377180 369288 377186 369300
rect 419534 369288 419540 369300
rect 377180 369260 419540 369288
rect 377180 369248 377186 369260
rect 419534 369248 419540 369260
rect 419592 369248 419598 369300
rect 99282 369180 99288 369232
rect 99340 369220 99346 369232
rect 211614 369220 211620 369232
rect 99340 369192 211620 369220
rect 99340 369180 99346 369192
rect 211614 369180 211620 369192
rect 211672 369220 211678 369232
rect 212534 369220 212540 369232
rect 211672 369192 212540 369220
rect 211672 369180 211678 369192
rect 212534 369180 212540 369192
rect 212592 369180 212598 369232
rect 366266 369180 366272 369232
rect 366324 369220 366330 369232
rect 371786 369220 371792 369232
rect 366324 369192 371792 369220
rect 366324 369180 366330 369192
rect 371786 369180 371792 369192
rect 371844 369220 371850 369232
rect 420914 369220 420920 369232
rect 371844 369192 420920 369220
rect 371844 369180 371850 369192
rect 420914 369180 420920 369192
rect 420972 369180 420978 369232
rect 97718 369112 97724 369164
rect 97776 369152 97782 369164
rect 210234 369152 210240 369164
rect 97776 369124 210240 369152
rect 97776 369112 97782 369124
rect 210234 369112 210240 369124
rect 210292 369152 210298 369164
rect 212626 369152 212632 369164
rect 210292 369124 212632 369152
rect 210292 369112 210298 369124
rect 212626 369112 212632 369124
rect 212684 369112 212690 369164
rect 359550 369112 359556 369164
rect 359608 369152 359614 369164
rect 360102 369152 360108 369164
rect 359608 369124 360108 369152
rect 359608 369112 359614 369124
rect 360102 369112 360108 369124
rect 360160 369152 360166 369164
rect 519078 369152 519084 369164
rect 360160 369124 519084 369152
rect 360160 369112 360166 369124
rect 519078 369112 519084 369124
rect 519136 369112 519142 369164
rect 206278 369044 206284 369096
rect 206336 369084 206342 369096
rect 249886 369084 249892 369096
rect 206336 369056 249892 369084
rect 206336 369044 206342 369056
rect 249886 369044 249892 369056
rect 249944 369044 249950 369096
rect 368290 369044 368296 369096
rect 368348 369084 368354 369096
rect 376662 369084 376668 369096
rect 368348 369056 376668 369084
rect 368348 369044 368354 369056
rect 376662 369044 376668 369056
rect 376720 369084 376726 369096
rect 418338 369084 418344 369096
rect 376720 369056 418344 369084
rect 376720 369044 376726 369056
rect 418338 369044 418344 369056
rect 418396 369044 418402 369096
rect 106182 368976 106188 369028
rect 106240 369016 106246 369028
rect 208394 369016 208400 369028
rect 106240 368988 208400 369016
rect 106240 368976 106246 368988
rect 208394 368976 208400 368988
rect 208452 368976 208458 369028
rect 213086 368976 213092 369028
rect 213144 369016 213150 369028
rect 276014 369016 276020 369028
rect 213144 368988 276020 369016
rect 213144 368976 213150 368988
rect 276014 368976 276020 368988
rect 276072 368976 276078 369028
rect 361298 368976 361304 369028
rect 361356 369016 361362 369028
rect 378686 369016 378692 369028
rect 361356 368988 378692 369016
rect 361356 368976 361362 368988
rect 378686 368976 378692 368988
rect 378744 369016 378750 369028
rect 405734 369016 405740 369028
rect 378744 368988 405740 369016
rect 378744 368976 378750 368988
rect 405734 368976 405740 368988
rect 405792 368976 405798 369028
rect 208026 368908 208032 368960
rect 208084 368948 208090 368960
rect 252554 368948 252560 368960
rect 208084 368920 252560 368948
rect 208084 368908 208090 368920
rect 252554 368908 252560 368920
rect 252612 368908 252618 368960
rect 370314 368908 370320 368960
rect 370372 368948 370378 368960
rect 480254 368948 480260 368960
rect 370372 368920 480260 368948
rect 370372 368908 370378 368920
rect 480254 368908 480260 368920
rect 480312 368908 480318 368960
rect 208854 368840 208860 368892
rect 208912 368880 208918 368892
rect 255314 368880 255320 368892
rect 208912 368852 255320 368880
rect 208912 368840 208918 368852
rect 255314 368840 255320 368852
rect 255372 368840 255378 368892
rect 101030 368772 101036 368824
rect 101088 368812 101094 368824
rect 214098 368812 214104 368824
rect 101088 368784 214104 368812
rect 101088 368772 101094 368784
rect 214098 368772 214104 368784
rect 214156 368812 214162 368824
rect 214466 368812 214472 368824
rect 214156 368784 214472 368812
rect 214156 368772 214162 368784
rect 214466 368772 214472 368784
rect 214524 368772 214530 368824
rect 54478 368636 54484 368688
rect 54536 368676 54542 368688
rect 55858 368676 55864 368688
rect 54536 368648 55864 368676
rect 54536 368636 54542 368648
rect 55858 368636 55864 368648
rect 55916 368636 55922 368688
rect 215294 368432 215300 368484
rect 215352 368472 215358 368484
rect 216582 368472 216588 368484
rect 215352 368444 216588 368472
rect 215352 368432 215358 368444
rect 216582 368432 216588 368444
rect 216640 368472 216646 368484
rect 219710 368472 219716 368484
rect 216640 368444 219716 368472
rect 216640 368432 216646 368444
rect 219710 368432 219716 368444
rect 219768 368472 219774 368484
rect 266354 368472 266360 368484
rect 219768 368444 266360 368472
rect 219768 368432 219774 368444
rect 266354 368432 266360 368444
rect 266412 368432 266418 368484
rect 365530 368092 365536 368144
rect 365588 368132 365594 368144
rect 379330 368132 379336 368144
rect 365588 368104 379336 368132
rect 365588 368092 365594 368104
rect 379330 368092 379336 368104
rect 379388 368132 379394 368144
rect 412634 368132 412640 368144
rect 379388 368104 412640 368132
rect 379388 368092 379394 368104
rect 412634 368092 412640 368104
rect 412692 368092 412698 368144
rect 357894 368024 357900 368076
rect 357952 368064 357958 368076
rect 368382 368064 368388 368076
rect 357952 368036 368388 368064
rect 357952 368024 357958 368036
rect 368382 368024 368388 368036
rect 368440 368064 368446 368076
rect 427906 368064 427912 368076
rect 368440 368036 427912 368064
rect 368440 368024 368446 368036
rect 427906 368024 427912 368036
rect 427964 368024 427970 368076
rect 357066 367956 357072 368008
rect 357124 367996 357130 368008
rect 375098 367996 375104 368008
rect 357124 367968 375104 367996
rect 357124 367956 357130 367968
rect 375098 367956 375104 367968
rect 375156 367996 375162 368008
rect 436094 367996 436100 368008
rect 375156 367968 436100 367996
rect 375156 367956 375162 367968
rect 436094 367956 436100 367968
rect 436152 367956 436158 368008
rect 362770 367888 362776 367940
rect 362828 367928 362834 367940
rect 370406 367928 370412 367940
rect 362828 367900 370412 367928
rect 362828 367888 362834 367900
rect 370406 367888 370412 367900
rect 370464 367928 370470 367940
rect 431954 367928 431960 367940
rect 370464 367900 431960 367928
rect 370464 367888 370470 367900
rect 431954 367888 431960 367900
rect 432012 367888 432018 367940
rect 364242 367820 364248 367872
rect 364300 367860 364306 367872
rect 368290 367860 368296 367872
rect 364300 367832 368296 367860
rect 364300 367820 364306 367832
rect 368290 367820 368296 367832
rect 368348 367860 368354 367872
rect 434714 367860 434720 367872
rect 368348 367832 434720 367860
rect 368348 367820 368354 367832
rect 434714 367820 434720 367832
rect 434772 367820 434778 367872
rect 107562 367752 107568 367804
rect 107620 367792 107626 367804
rect 215294 367792 215300 367804
rect 107620 367764 215300 367792
rect 107620 367752 107626 367764
rect 215294 367752 215300 367764
rect 215352 367752 215358 367804
rect 358998 367752 359004 367804
rect 359056 367792 359062 367804
rect 359918 367792 359924 367804
rect 359056 367764 359924 367792
rect 359056 367752 359062 367764
rect 359918 367752 359924 367764
rect 359976 367792 359982 367804
rect 519170 367792 519176 367804
rect 359976 367764 519176 367792
rect 359976 367752 359982 367764
rect 519170 367752 519176 367764
rect 519228 367752 519234 367804
rect 199378 366324 199384 366376
rect 199436 366364 199442 366376
rect 199746 366364 199752 366376
rect 199436 366336 199752 366364
rect 199436 366324 199442 366336
rect 199746 366324 199752 366336
rect 199804 366364 199810 366376
rect 358998 366364 359004 366376
rect 199804 366336 359004 366364
rect 199804 366324 199810 366336
rect 358998 366324 359004 366336
rect 359056 366324 359062 366376
rect 201034 364284 201040 364336
rect 201092 364324 201098 364336
rect 343082 364324 343088 364336
rect 201092 364296 343088 364324
rect 201092 364284 201098 364296
rect 343082 364284 343088 364296
rect 343140 364284 343146 364336
rect 199470 362176 199476 362228
rect 199528 362216 199534 362228
rect 359090 362216 359096 362228
rect 199528 362188 359096 362216
rect 199528 362176 199534 362188
rect 359090 362176 359096 362188
rect 359148 362216 359154 362228
rect 359458 362216 359464 362228
rect 359148 362188 359464 362216
rect 359148 362176 359154 362188
rect 359458 362176 359464 362188
rect 359516 362176 359522 362228
rect 208394 360136 208400 360188
rect 208452 360176 208458 360188
rect 209682 360176 209688 360188
rect 208452 360148 209688 360176
rect 208452 360136 208458 360148
rect 209682 360136 209688 360148
rect 209740 360176 209746 360188
rect 359182 360176 359188 360188
rect 209740 360148 359188 360176
rect 209740 360136 209746 360148
rect 359182 360136 359188 360148
rect 359240 360136 359246 360188
rect 199746 359456 199752 359508
rect 199804 359496 199810 359508
rect 208394 359496 208400 359508
rect 199804 359468 208400 359496
rect 199804 359456 199810 359468
rect 208394 359456 208400 359468
rect 208452 359456 208458 359508
rect 359274 359456 359280 359508
rect 359332 359496 359338 359508
rect 359826 359496 359832 359508
rect 359332 359468 359832 359496
rect 359332 359456 359338 359468
rect 359826 359456 359832 359468
rect 359884 359496 359890 359508
rect 519262 359496 519268 359508
rect 359884 359468 519268 359496
rect 359884 359456 359890 359468
rect 519262 359456 519268 359468
rect 519320 359456 519326 359508
rect 3326 358708 3332 358760
rect 3384 358748 3390 358760
rect 18598 358748 18604 358760
rect 3384 358720 18604 358748
rect 3384 358708 3390 358720
rect 18598 358708 18604 358720
rect 18656 358708 18662 358760
rect 359458 358096 359464 358148
rect 359516 358136 359522 358148
rect 519354 358136 519360 358148
rect 359516 358108 519360 358136
rect 359516 358096 359522 358108
rect 519354 358096 519360 358108
rect 519412 358096 519418 358148
rect 199562 358028 199568 358080
rect 199620 358068 199626 358080
rect 359274 358068 359280 358080
rect 199620 358040 359280 358068
rect 199620 358028 199626 358040
rect 359274 358028 359280 358040
rect 359332 358028 359338 358080
rect 182818 356668 182824 356720
rect 182876 356708 182882 356720
rect 202874 356708 202880 356720
rect 182876 356680 202880 356708
rect 182876 356668 182882 356680
rect 202874 356668 202880 356680
rect 202932 356708 202938 356720
rect 342898 356708 342904 356720
rect 202932 356680 342904 356708
rect 202932 356668 202938 356680
rect 342898 356668 342904 356680
rect 342956 356668 342962 356720
rect 206922 356096 206928 356108
rect 205652 356068 206928 356096
rect 191374 355988 191380 356040
rect 191432 356028 191438 356040
rect 205652 356028 205680 356068
rect 206922 356056 206928 356068
rect 206980 356096 206986 356108
rect 215938 356096 215944 356108
rect 206980 356068 215944 356096
rect 206980 356056 206986 356068
rect 215938 356056 215944 356068
rect 215996 356056 216002 356108
rect 191432 356000 205680 356028
rect 191432 355988 191438 356000
rect 357342 355988 357348 356040
rect 357400 356028 357406 356040
rect 362954 356028 362960 356040
rect 357400 356000 362960 356028
rect 357400 355988 357406 356000
rect 362954 355988 362960 356000
rect 363012 355988 363018 356040
rect 179782 355920 179788 355972
rect 179840 355960 179846 355972
rect 195882 355960 195888 355972
rect 179840 355932 195888 355960
rect 179840 355920 179846 355932
rect 195882 355920 195888 355932
rect 195940 355920 195946 355972
rect 500862 355444 500868 355496
rect 500920 355484 500926 355496
rect 517606 355484 517612 355496
rect 500920 355456 517612 355484
rect 500920 355444 500926 355456
rect 517606 355444 517612 355456
rect 517664 355444 517670 355496
rect 340046 355376 340052 355428
rect 340104 355416 340110 355428
rect 356606 355416 356612 355428
rect 340104 355388 356612 355416
rect 340104 355376 340110 355388
rect 356606 355376 356612 355388
rect 356664 355376 356670 355428
rect 498838 355376 498844 355428
rect 498896 355416 498902 355428
rect 517698 355416 517704 355428
rect 498896 355388 517704 355416
rect 498896 355376 498902 355388
rect 517698 355376 517704 355388
rect 517756 355376 517762 355428
rect 351730 355308 351736 355360
rect 351788 355348 351794 355360
rect 358078 355348 358084 355360
rect 351788 355320 358084 355348
rect 351788 355308 351794 355320
rect 358078 355308 358084 355320
rect 358136 355308 358142 355360
rect 195882 355172 195888 355224
rect 195940 355212 195946 355224
rect 197354 355212 197360 355224
rect 195940 355184 197360 355212
rect 195940 355172 195946 355184
rect 197354 355172 197360 355184
rect 197412 355172 197418 355224
rect 356606 354968 356612 355020
rect 356664 355008 356670 355020
rect 356882 355008 356888 355020
rect 356664 354980 356888 355008
rect 356664 354968 356670 354980
rect 356882 354968 356888 354980
rect 356940 354968 356946 355020
rect 338114 354764 338120 354816
rect 338172 354804 338178 354816
rect 357342 354804 357348 354816
rect 338172 354776 357348 354804
rect 338172 354764 338178 354776
rect 357342 354764 357348 354776
rect 357400 354764 357406 354816
rect 510890 354764 510896 354816
rect 510948 354804 510954 354816
rect 517514 354804 517520 354816
rect 510948 354776 517520 354804
rect 510948 354764 510954 354776
rect 517514 354764 517520 354776
rect 517572 354764 517578 354816
rect 178586 354696 178592 354748
rect 178644 354736 178650 354748
rect 197722 354736 197728 354748
rect 178644 354708 197728 354736
rect 178644 354696 178650 354708
rect 197722 354696 197728 354708
rect 197780 354736 197786 354748
rect 201954 354736 201960 354748
rect 197780 354708 201960 354736
rect 197780 354696 197786 354708
rect 201954 354696 201960 354708
rect 202012 354696 202018 354748
rect 199654 353948 199660 354000
rect 199712 353988 199718 354000
rect 359550 353988 359556 354000
rect 199712 353960 359556 353988
rect 199712 353948 199718 353960
rect 359550 353948 359556 353960
rect 359608 353948 359614 354000
rect 373166 353948 373172 354000
rect 373224 353988 373230 354000
rect 381078 353988 381084 354000
rect 373224 353960 381084 353988
rect 373224 353948 373230 353960
rect 381078 353948 381084 353960
rect 381136 353948 381142 354000
rect 217870 353404 217876 353456
rect 217928 353444 217934 353456
rect 220814 353444 220820 353456
rect 217928 353416 220820 353444
rect 217928 353404 217934 353416
rect 220814 353404 220820 353416
rect 220872 353404 220878 353456
rect 55858 353336 55864 353388
rect 55916 353376 55922 353388
rect 60734 353376 60740 353388
rect 55916 353348 60740 353376
rect 55916 353336 55922 353348
rect 60734 353336 60740 353348
rect 60792 353336 60798 353388
rect 218606 353336 218612 353388
rect 218664 353376 218670 353388
rect 220906 353376 220912 353388
rect 218664 353348 220912 353376
rect 218664 353336 218670 353348
rect 220906 353336 220912 353348
rect 220964 353336 220970 353388
rect 378594 353336 378600 353388
rect 378652 353376 378658 353388
rect 380894 353376 380900 353388
rect 378652 353348 380900 353376
rect 378652 353336 378658 353348
rect 380894 353336 380900 353348
rect 380952 353336 380958 353388
rect 58618 353268 58624 353320
rect 58676 353308 58682 353320
rect 62114 353308 62120 353320
rect 58676 353280 62120 353308
rect 58676 353268 58682 353280
rect 62114 353268 62120 353280
rect 62172 353268 62178 353320
rect 219158 353268 219164 353320
rect 219216 353308 219222 353320
rect 220998 353308 221004 353320
rect 219216 353280 221004 353308
rect 219216 353268 219222 353280
rect 220998 353268 221004 353280
rect 221056 353268 221062 353320
rect 359182 353268 359188 353320
rect 359240 353308 359246 353320
rect 359550 353308 359556 353320
rect 359240 353280 359556 353308
rect 359240 353268 359246 353280
rect 359550 353268 359556 353280
rect 359608 353268 359614 353320
rect 379238 353268 379244 353320
rect 379296 353308 379302 353320
rect 380986 353308 380992 353320
rect 379296 353280 380992 353308
rect 379296 353268 379302 353280
rect 380986 353268 380992 353280
rect 381044 353268 381050 353320
rect 54386 352520 54392 352572
rect 54444 352560 54450 352572
rect 59446 352560 59452 352572
rect 54444 352532 59452 352560
rect 54444 352520 54450 352532
rect 59446 352520 59452 352532
rect 59504 352520 59510 352572
rect 56870 351908 56876 351960
rect 56928 351948 56934 351960
rect 59354 351948 59360 351960
rect 56928 351920 59360 351948
rect 56928 351908 56934 351920
rect 59354 351908 59360 351920
rect 59412 351908 59418 351960
rect 58526 350548 58532 350600
rect 58584 350588 58590 350600
rect 59722 350588 59728 350600
rect 58584 350560 59728 350588
rect 58584 350548 58590 350560
rect 59722 350548 59728 350560
rect 59780 350548 59786 350600
rect 47854 298052 47860 298104
rect 47912 298092 47918 298104
rect 57514 298092 57520 298104
rect 47912 298064 57520 298092
rect 47912 298052 47918 298064
rect 57514 298052 57520 298064
rect 57572 298052 57578 298104
rect 520182 284316 520188 284368
rect 520240 284356 520246 284368
rect 580258 284356 580264 284368
rect 520240 284328 580264 284356
rect 520240 284316 520246 284328
rect 580258 284316 580264 284328
rect 580316 284316 580322 284368
rect 519078 282888 519084 282940
rect 519136 282928 519142 282940
rect 580350 282928 580356 282940
rect 519136 282900 580356 282928
rect 519136 282888 519142 282900
rect 580350 282888 580356 282900
rect 580408 282888 580414 282940
rect 200942 280100 200948 280152
rect 201000 280140 201006 280152
rect 216674 280140 216680 280152
rect 201000 280112 216680 280140
rect 201000 280100 201006 280112
rect 216674 280100 216680 280112
rect 216732 280100 216738 280152
rect 55674 278672 55680 278724
rect 55732 278712 55738 278724
rect 58710 278712 58716 278724
rect 55732 278684 58716 278712
rect 55732 278672 55738 278684
rect 58710 278672 58716 278684
rect 58768 278672 58774 278724
rect 206738 278672 206744 278724
rect 206796 278712 206802 278724
rect 216674 278712 216680 278724
rect 206796 278684 216680 278712
rect 206796 278672 206802 278684
rect 216674 278672 216680 278684
rect 216732 278672 216738 278724
rect 361206 278672 361212 278724
rect 361264 278712 361270 278724
rect 376754 278712 376760 278724
rect 361264 278684 376760 278712
rect 361264 278672 361270 278684
rect 376754 278672 376760 278684
rect 376812 278672 376818 278724
rect 215938 278264 215944 278316
rect 215996 278304 216002 278316
rect 216950 278304 216956 278316
rect 215996 278276 216956 278304
rect 215996 278264 216002 278276
rect 216950 278264 216956 278276
rect 217008 278264 217014 278316
rect 358078 277992 358084 278044
rect 358136 278032 358142 278044
rect 376846 278032 376852 278044
rect 358136 278004 376852 278032
rect 358136 277992 358142 278004
rect 376846 277992 376852 278004
rect 376904 277992 376910 278044
rect 378594 270444 378600 270496
rect 378652 270484 378658 270496
rect 379606 270484 379612 270496
rect 378652 270456 379612 270484
rect 378652 270444 378658 270456
rect 379606 270444 379612 270456
rect 379664 270444 379670 270496
rect 51442 269764 51448 269816
rect 51500 269804 51506 269816
rect 54478 269804 54484 269816
rect 51500 269776 54484 269804
rect 51500 269764 51506 269776
rect 54478 269764 54484 269776
rect 54536 269804 54542 269816
rect 55214 269804 55220 269816
rect 54536 269776 55220 269804
rect 54536 269764 54542 269776
rect 55214 269764 55220 269776
rect 55272 269764 55278 269816
rect 373166 269764 373172 269816
rect 373224 269804 373230 269816
rect 374454 269804 374460 269816
rect 373224 269776 374460 269804
rect 373224 269764 373230 269776
rect 374454 269764 374460 269776
rect 374512 269764 374518 269816
rect 45186 269696 45192 269748
rect 45244 269736 45250 269748
rect 148502 269736 148508 269748
rect 45244 269708 148508 269736
rect 45244 269696 45250 269708
rect 148502 269696 148508 269708
rect 148560 269696 148566 269748
rect 46198 269628 46204 269680
rect 46256 269668 46262 269680
rect 59814 269668 59820 269680
rect 46256 269640 59820 269668
rect 46256 269628 46262 269640
rect 59814 269628 59820 269640
rect 59872 269668 59878 269680
rect 60090 269668 60096 269680
rect 59872 269640 60096 269668
rect 59872 269628 59878 269640
rect 60090 269628 60096 269640
rect 60148 269628 60154 269680
rect 51534 269560 51540 269612
rect 51592 269600 51598 269612
rect 51718 269600 51724 269612
rect 51592 269572 51724 269600
rect 51592 269560 51598 269572
rect 51718 269560 51724 269572
rect 51776 269560 51782 269612
rect 52914 269560 52920 269612
rect 52972 269600 52978 269612
rect 110966 269600 110972 269612
rect 52972 269572 110972 269600
rect 52972 269560 52978 269572
rect 110966 269560 110972 269572
rect 111024 269560 111030 269612
rect 43530 269492 43536 269544
rect 43588 269532 43594 269544
rect 133414 269532 133420 269544
rect 43588 269504 133420 269532
rect 43588 269492 43594 269504
rect 133414 269492 133420 269504
rect 133472 269492 133478 269544
rect 379606 269492 379612 269544
rect 379664 269532 379670 269544
rect 425238 269532 425244 269544
rect 379664 269504 425244 269532
rect 379664 269492 379670 269504
rect 425238 269492 425244 269504
rect 425296 269492 425302 269544
rect 44910 269424 44916 269476
rect 44968 269464 44974 269476
rect 135898 269464 135904 269476
rect 44968 269436 135904 269464
rect 44968 269424 44974 269436
rect 135898 269424 135904 269436
rect 135956 269424 135962 269476
rect 363966 269424 363972 269476
rect 364024 269464 364030 269476
rect 416038 269464 416044 269476
rect 364024 269436 416044 269464
rect 364024 269424 364030 269436
rect 416038 269424 416044 269436
rect 416096 269424 416102 269476
rect 45002 269356 45008 269408
rect 45060 269396 45066 269408
rect 138474 269396 138480 269408
rect 45060 269368 138480 269396
rect 45060 269356 45066 269368
rect 138474 269356 138480 269368
rect 138532 269356 138538 269408
rect 374454 269356 374460 269408
rect 374512 269396 374518 269408
rect 433334 269396 433340 269408
rect 374512 269368 433340 269396
rect 374512 269356 374518 269368
rect 433334 269356 433340 269368
rect 433392 269356 433398 269408
rect 45094 269288 45100 269340
rect 45152 269328 45158 269340
rect 140866 269328 140872 269340
rect 45152 269300 140872 269328
rect 45152 269288 45158 269300
rect 140866 269288 140872 269300
rect 140924 269288 140930 269340
rect 210786 269288 210792 269340
rect 210844 269328 210850 269340
rect 250714 269328 250720 269340
rect 210844 269300 250720 269328
rect 210844 269288 210850 269300
rect 250714 269288 250720 269300
rect 250772 269288 250778 269340
rect 371694 269288 371700 269340
rect 371752 269328 371758 269340
rect 372522 269328 372528 269340
rect 371752 269300 372528 269328
rect 371752 269288 371758 269300
rect 372522 269288 372528 269300
rect 372580 269328 372586 269340
rect 434346 269328 434352 269340
rect 372580 269300 434352 269328
rect 372580 269288 372586 269300
rect 434346 269288 434352 269300
rect 434404 269288 434410 269340
rect 45370 269220 45376 269272
rect 45428 269260 45434 269272
rect 143534 269260 143540 269272
rect 45428 269232 143540 269260
rect 45428 269220 45434 269232
rect 143534 269220 143540 269232
rect 143592 269220 143598 269272
rect 205266 269220 205272 269272
rect 205324 269260 205330 269272
rect 283466 269260 283472 269272
rect 205324 269232 283472 269260
rect 205324 269220 205330 269232
rect 283466 269220 283472 269232
rect 283524 269220 283530 269272
rect 370958 269220 370964 269272
rect 371016 269260 371022 269272
rect 436002 269260 436008 269272
rect 371016 269232 436008 269260
rect 371016 269220 371022 269232
rect 436002 269220 436008 269232
rect 436060 269220 436066 269272
rect 45278 269152 45284 269204
rect 45336 269192 45342 269204
rect 145926 269192 145932 269204
rect 45336 269164 145932 269192
rect 45336 269152 45342 269164
rect 145926 269152 145932 269164
rect 145984 269152 145990 269204
rect 206646 269152 206652 269204
rect 206704 269192 206710 269204
rect 288250 269192 288256 269204
rect 206704 269164 288256 269192
rect 206704 269152 206710 269164
rect 288250 269152 288256 269164
rect 288308 269152 288314 269204
rect 372522 269152 372528 269204
rect 372580 269192 372586 269204
rect 373994 269192 374000 269204
rect 372580 269164 374000 269192
rect 372580 269152 372586 269164
rect 373994 269152 374000 269164
rect 374052 269192 374058 269204
rect 374454 269192 374460 269204
rect 374052 269164 374460 269192
rect 374052 269152 374058 269164
rect 374454 269152 374460 269164
rect 374512 269152 374518 269204
rect 375006 269152 375012 269204
rect 375064 269192 375070 269204
rect 468478 269192 468484 269204
rect 375064 269164 468484 269192
rect 375064 269152 375070 269164
rect 468478 269152 468484 269164
rect 468536 269152 468542 269204
rect 91278 269124 91284 269136
rect 62132 269096 91284 269124
rect 45462 269016 45468 269068
rect 45520 269056 45526 269068
rect 45520 269016 45554 269056
rect 50338 269016 50344 269068
rect 50396 269056 50402 269068
rect 51718 269056 51724 269068
rect 50396 269028 51724 269056
rect 50396 269016 50402 269028
rect 51718 269016 51724 269028
rect 51776 269016 51782 269068
rect 45526 268988 45554 269016
rect 62132 269000 62160 269096
rect 91278 269084 91284 269096
rect 91336 269084 91342 269136
rect 207934 269084 207940 269136
rect 207992 269124 207998 269136
rect 291010 269124 291016 269136
rect 207992 269096 291016 269124
rect 207992 269084 207998 269096
rect 291010 269084 291016 269096
rect 291068 269084 291074 269136
rect 365346 269084 365352 269136
rect 365404 269124 365410 269136
rect 470962 269124 470968 269136
rect 365404 269096 470968 269124
rect 365404 269084 365410 269096
rect 470962 269084 470968 269096
rect 471020 269084 471026 269136
rect 196618 269016 196624 269068
rect 196676 269056 196682 269068
rect 197170 269056 197176 269068
rect 196676 269028 197176 269056
rect 196676 269016 196682 269028
rect 197170 269016 197176 269028
rect 197228 269016 197234 269068
rect 213546 269016 213552 269068
rect 213604 269056 213610 269068
rect 215386 269056 215392 269068
rect 213604 269028 215392 269056
rect 213604 269016 213610 269028
rect 215386 269016 215392 269028
rect 215444 269016 215450 269068
rect 373074 269016 373080 269068
rect 373132 269056 373138 269068
rect 373718 269056 373724 269068
rect 373132 269028 373724 269056
rect 373132 269016 373138 269028
rect 373718 269016 373724 269028
rect 373776 269016 373782 269068
rect 379514 269016 379520 269068
rect 379572 269056 379578 269068
rect 379790 269056 379796 269068
rect 379572 269028 379796 269056
rect 379572 269016 379578 269028
rect 379790 269016 379796 269028
rect 379848 269016 379854 269068
rect 62114 268988 62120 269000
rect 45526 268960 62120 268988
rect 62114 268948 62120 268960
rect 62172 268948 62178 269000
rect 211614 268948 211620 269000
rect 211672 268988 211678 269000
rect 216950 268988 216956 269000
rect 211672 268960 216956 268988
rect 211672 268948 211678 268960
rect 216950 268948 216956 268960
rect 217008 268948 217014 269000
rect 46474 268880 46480 268932
rect 46532 268920 46538 268932
rect 54662 268920 54668 268932
rect 46532 268892 54668 268920
rect 46532 268880 46538 268892
rect 54662 268880 54668 268892
rect 54720 268880 54726 268932
rect 213454 268880 213460 268932
rect 213512 268920 213518 268932
rect 235994 268920 236000 268932
rect 213512 268892 236000 268920
rect 213512 268880 213518 268892
rect 235994 268880 236000 268892
rect 236052 268880 236058 268932
rect 212166 268812 212172 268864
rect 212224 268852 212230 268864
rect 298462 268852 298468 268864
rect 212224 268824 298468 268852
rect 212224 268812 212230 268824
rect 298462 268812 298468 268824
rect 298520 268812 298526 268864
rect 374454 268812 374460 268864
rect 374512 268852 374518 268864
rect 422846 268852 422852 268864
rect 374512 268824 422852 268852
rect 374512 268812 374518 268824
rect 422846 268812 422852 268824
rect 422904 268812 422910 268864
rect 209314 268744 209320 268796
rect 209372 268784 209378 268796
rect 295886 268784 295892 268796
rect 209372 268756 295892 268784
rect 209372 268744 209378 268756
rect 295886 268744 295892 268756
rect 295944 268744 295950 268796
rect 368106 268744 368112 268796
rect 368164 268784 368170 268796
rect 430942 268784 430948 268796
rect 368164 268756 430948 268784
rect 368164 268744 368170 268756
rect 430942 268744 430948 268756
rect 431000 268744 431006 268796
rect 60090 268676 60096 268728
rect 60148 268716 60154 268728
rect 94498 268716 94504 268728
rect 60148 268688 94504 268716
rect 60148 268676 60154 268688
rect 94498 268676 94504 268688
rect 94556 268676 94562 268728
rect 202322 268676 202328 268728
rect 202380 268716 202386 268728
rect 293402 268716 293408 268728
rect 202380 268688 293408 268716
rect 202380 268676 202386 268688
rect 293402 268676 293408 268688
rect 293460 268676 293466 268728
rect 361022 268676 361028 268728
rect 361080 268716 361086 268728
rect 425974 268716 425980 268728
rect 361080 268688 425980 268716
rect 361080 268676 361086 268688
rect 425974 268676 425980 268688
rect 426032 268676 426038 268728
rect 58526 268608 58532 268660
rect 58584 268648 58590 268660
rect 93578 268648 93584 268660
rect 58584 268620 93584 268648
rect 58584 268608 58590 268620
rect 93578 268608 93584 268620
rect 93636 268608 93642 268660
rect 203794 268608 203800 268660
rect 203852 268648 203858 268660
rect 300854 268648 300860 268660
rect 203852 268620 300860 268648
rect 203852 268608 203858 268620
rect 300854 268608 300860 268620
rect 300912 268608 300918 268660
rect 356790 268608 356796 268660
rect 356848 268648 356854 268660
rect 421006 268648 421012 268660
rect 356848 268620 421012 268648
rect 356848 268608 356854 268620
rect 421006 268608 421012 268620
rect 421064 268608 421070 268660
rect 48038 268540 48044 268592
rect 48096 268580 48102 268592
rect 90726 268580 90732 268592
rect 48096 268552 90732 268580
rect 48096 268540 48102 268552
rect 90726 268540 90732 268552
rect 90784 268540 90790 268592
rect 205174 268540 205180 268592
rect 205232 268580 205238 268592
rect 305914 268580 305920 268592
rect 205232 268552 305920 268580
rect 205232 268540 205238 268552
rect 305914 268540 305920 268552
rect 305972 268540 305978 268592
rect 366910 268540 366916 268592
rect 366968 268580 366974 268592
rect 475838 268580 475844 268592
rect 366968 268552 475844 268580
rect 366968 268540 366974 268552
rect 475838 268540 475844 268552
rect 475896 268540 475902 268592
rect 51902 268472 51908 268524
rect 51960 268512 51966 268524
rect 98454 268512 98460 268524
rect 51960 268484 98460 268512
rect 51960 268472 51966 268484
rect 98454 268472 98460 268484
rect 98512 268472 98518 268524
rect 200758 268472 200764 268524
rect 200816 268512 200822 268524
rect 303430 268512 303436 268524
rect 200816 268484 303436 268512
rect 200816 268472 200822 268484
rect 303430 268472 303436 268484
rect 303488 268472 303494 268524
rect 369578 268472 369584 268524
rect 369636 268512 369642 268524
rect 478414 268512 478420 268524
rect 369636 268484 478420 268512
rect 369636 268472 369642 268484
rect 478414 268472 478420 268484
rect 478472 268472 478478 268524
rect 49050 268404 49056 268456
rect 49108 268444 49114 268456
rect 96062 268444 96068 268456
rect 49108 268416 96068 268444
rect 49108 268404 49114 268416
rect 96062 268404 96068 268416
rect 96120 268404 96126 268456
rect 209498 268404 209504 268456
rect 209556 268444 209562 268456
rect 214466 268444 214472 268456
rect 209556 268416 214472 268444
rect 209556 268404 209562 268416
rect 214466 268404 214472 268416
rect 214524 268404 214530 268456
rect 214926 268404 214932 268456
rect 214984 268444 214990 268456
rect 323302 268444 323308 268456
rect 214984 268416 323308 268444
rect 214984 268404 214990 268416
rect 323302 268404 323308 268416
rect 323360 268404 323366 268456
rect 372154 268404 372160 268456
rect 372212 268444 372218 268456
rect 480898 268444 480904 268456
rect 372212 268416 480904 268444
rect 372212 268404 372218 268416
rect 480898 268404 480904 268416
rect 480956 268404 480962 268456
rect 51534 268336 51540 268388
rect 51592 268376 51598 268388
rect 53742 268376 53748 268388
rect 51592 268348 53748 268376
rect 51592 268336 51598 268348
rect 53742 268336 53748 268348
rect 53800 268336 53806 268388
rect 55214 268336 55220 268388
rect 55272 268376 55278 268388
rect 100754 268376 100760 268388
rect 55272 268348 100760 268376
rect 55272 268336 55278 268348
rect 100754 268336 100760 268348
rect 100812 268336 100818 268388
rect 197998 268336 198004 268388
rect 198056 268376 198062 268388
rect 318426 268376 318432 268388
rect 198056 268348 318432 268376
rect 198056 268336 198062 268348
rect 318426 268336 318432 268348
rect 318484 268336 318490 268388
rect 362678 268336 362684 268388
rect 362736 268376 362742 268388
rect 483382 268376 483388 268388
rect 362736 268348 483388 268376
rect 362736 268336 362742 268348
rect 483382 268336 483388 268348
rect 483440 268336 483446 268388
rect 48130 268200 48136 268252
rect 48188 268240 48194 268252
rect 77110 268240 77116 268252
rect 48188 268212 77116 268240
rect 48188 268200 48194 268212
rect 77110 268200 77116 268212
rect 77168 268200 77174 268252
rect 373718 268200 373724 268252
rect 373776 268240 373782 268252
rect 429746 268240 429752 268252
rect 373776 268212 429752 268240
rect 373776 268200 373782 268212
rect 429746 268200 429752 268212
rect 429804 268200 429810 268252
rect 54202 268132 54208 268184
rect 54260 268172 54266 268184
rect 54478 268172 54484 268184
rect 54260 268144 54484 268172
rect 54260 268132 54266 268144
rect 54478 268132 54484 268144
rect 54536 268132 54542 268184
rect 66254 268132 66260 268184
rect 66312 268172 66318 268184
rect 95878 268172 95884 268184
rect 66312 268144 95884 268172
rect 66312 268132 66318 268144
rect 95878 268132 95884 268144
rect 95936 268132 95942 268184
rect 373166 268132 373172 268184
rect 373224 268172 373230 268184
rect 432230 268172 432236 268184
rect 373224 268144 432236 268172
rect 373224 268132 373230 268144
rect 432230 268132 432236 268144
rect 432288 268132 432294 268184
rect 46382 268064 46388 268116
rect 46440 268104 46446 268116
rect 76006 268104 76012 268116
rect 46440 268076 76012 268104
rect 46440 268064 46446 268076
rect 76006 268064 76012 268076
rect 76064 268064 76070 268116
rect 79318 268064 79324 268116
rect 79376 268104 79382 268116
rect 106366 268104 106372 268116
rect 79376 268076 106372 268104
rect 79376 268064 79382 268076
rect 106366 268064 106372 268076
rect 106424 268064 106430 268116
rect 396718 268064 396724 268116
rect 396776 268104 396782 268116
rect 415394 268104 415400 268116
rect 396776 268076 415400 268104
rect 396776 268064 396782 268076
rect 415394 268064 415400 268076
rect 415452 268064 415458 268116
rect 48958 267996 48964 268048
rect 49016 268036 49022 268048
rect 83090 268036 83096 268048
rect 49016 268008 83096 268036
rect 49016 267996 49022 268008
rect 83090 267996 83096 268008
rect 83148 267996 83154 268048
rect 395338 267996 395344 268048
rect 395396 268036 395402 268048
rect 416958 268036 416964 268048
rect 395396 268008 416964 268036
rect 395396 267996 395402 268008
rect 416958 267996 416964 268008
rect 417016 267996 417022 268048
rect 54294 267928 54300 267980
rect 54352 267968 54358 267980
rect 54662 267968 54668 267980
rect 54352 267940 54668 267968
rect 54352 267928 54358 267940
rect 54662 267928 54668 267940
rect 54720 267968 54726 267980
rect 96982 267968 96988 267980
rect 54720 267940 96988 267968
rect 54720 267928 54726 267940
rect 96982 267928 96988 267940
rect 97040 267928 97046 267980
rect 235994 267928 236000 267980
rect 236052 267968 236058 267980
rect 247034 267968 247040 267980
rect 236052 267940 247040 267968
rect 236052 267928 236058 267940
rect 247034 267928 247040 267940
rect 247092 267928 247098 267980
rect 373810 267928 373816 267980
rect 373868 267968 373874 267980
rect 374270 267968 374276 267980
rect 373868 267940 374276 267968
rect 373868 267928 373874 267940
rect 374270 267928 374276 267940
rect 374328 267968 374334 267980
rect 402974 267968 402980 267980
rect 374328 267940 402980 267968
rect 374328 267928 374334 267940
rect 402974 267928 402980 267940
rect 403032 267928 403038 267980
rect 58710 267860 58716 267912
rect 58768 267900 58774 267912
rect 59814 267900 59820 267912
rect 58768 267872 59820 267900
rect 58768 267860 58774 267872
rect 59814 267860 59820 267872
rect 59872 267900 59878 267912
rect 102686 267900 102692 267912
rect 59872 267872 102692 267900
rect 59872 267860 59878 267872
rect 102686 267860 102692 267872
rect 102744 267860 102750 267912
rect 106918 267860 106924 267912
rect 106976 267900 106982 267912
rect 119062 267900 119068 267912
rect 106976 267872 119068 267900
rect 106976 267860 106982 267872
rect 119062 267860 119068 267872
rect 119120 267860 119126 267912
rect 215386 267860 215392 267912
rect 215444 267900 215450 267912
rect 243078 267900 243084 267912
rect 215444 267872 243084 267900
rect 215444 267860 215450 267872
rect 243078 267860 243084 267872
rect 243136 267860 243142 267912
rect 379514 267860 379520 267912
rect 379572 267900 379578 267912
rect 414382 267900 414388 267912
rect 379572 267872 414388 267900
rect 379572 267860 379578 267872
rect 414382 267860 414388 267872
rect 414440 267860 414446 267912
rect 54202 267792 54208 267844
rect 54260 267832 54266 267844
rect 99374 267832 99380 267844
rect 54260 267804 99380 267832
rect 54260 267792 54266 267804
rect 99374 267792 99380 267804
rect 99432 267792 99438 267844
rect 112346 267792 112352 267844
rect 112404 267832 112410 267844
rect 197906 267832 197912 267844
rect 112404 267804 197912 267832
rect 112404 267792 112410 267804
rect 197906 267792 197912 267804
rect 197964 267832 197970 267844
rect 201586 267832 201592 267844
rect 197964 267804 201592 267832
rect 197964 267792 197970 267804
rect 201586 267792 201592 267804
rect 201644 267792 201650 267844
rect 217962 267792 217968 267844
rect 218020 267832 218026 267844
rect 258074 267832 258080 267844
rect 218020 267804 258080 267832
rect 218020 267792 218026 267804
rect 258074 267792 258080 267804
rect 258132 267792 258138 267844
rect 427078 267792 427084 267844
rect 427136 267832 427142 267844
rect 434714 267832 434720 267844
rect 427136 267804 434720 267832
rect 427136 267792 427142 267804
rect 434714 267792 434720 267804
rect 434772 267792 434778 267844
rect 51442 267724 51448 267776
rect 51500 267764 51506 267776
rect 51718 267764 51724 267776
rect 51500 267736 51724 267764
rect 51500 267724 51506 267736
rect 51718 267724 51724 267736
rect 51776 267764 51782 267776
rect 97994 267764 98000 267776
rect 51776 267736 98000 267764
rect 51776 267724 51782 267736
rect 97994 267724 98000 267736
rect 98052 267724 98058 267776
rect 111242 267724 111248 267776
rect 111300 267764 111306 267776
rect 196618 267764 196624 267776
rect 111300 267736 196624 267764
rect 111300 267724 111306 267736
rect 196618 267724 196624 267736
rect 196676 267724 196682 267776
rect 214466 267724 214472 267776
rect 214524 267764 214530 267776
rect 261662 267764 261668 267776
rect 214524 267736 261668 267764
rect 214524 267724 214530 267736
rect 261662 267724 261668 267736
rect 261720 267724 261726 267776
rect 425698 267724 425704 267776
rect 425756 267764 425762 267776
rect 428550 267764 428556 267776
rect 425756 267736 428556 267764
rect 425756 267724 425762 267736
rect 428550 267724 428556 267736
rect 428608 267724 428614 267776
rect 43622 267656 43628 267708
rect 43680 267696 43686 267708
rect 128354 267696 128360 267708
rect 43680 267668 128360 267696
rect 43680 267656 43686 267668
rect 128354 267656 128360 267668
rect 128412 267656 128418 267708
rect 158530 267656 158536 267708
rect 158588 267696 158594 267708
rect 205634 267696 205640 267708
rect 158588 267668 205640 267696
rect 158588 267656 158594 267668
rect 205634 267656 205640 267668
rect 205692 267656 205698 267708
rect 247034 267656 247040 267708
rect 247092 267696 247098 267708
rect 255314 267696 255320 267708
rect 247092 267668 255320 267696
rect 247092 267656 247098 267668
rect 255314 267656 255320 267668
rect 255372 267656 255378 267708
rect 372246 267656 372252 267708
rect 372304 267696 372310 267708
rect 460934 267696 460940 267708
rect 372304 267668 460940 267696
rect 372304 267656 372310 267668
rect 460934 267656 460940 267668
rect 460992 267656 460998 267708
rect 42242 267588 42248 267640
rect 42300 267628 42306 267640
rect 125594 267628 125600 267640
rect 42300 267600 125600 267628
rect 42300 267588 42306 267600
rect 125594 267588 125600 267600
rect 125652 267588 125658 267640
rect 150986 267588 150992 267640
rect 151044 267628 151050 267640
rect 198090 267628 198096 267640
rect 151044 267600 198096 267628
rect 151044 267588 151050 267600
rect 198090 267588 198096 267600
rect 198148 267588 198154 267640
rect 209222 267588 209228 267640
rect 209280 267628 209286 267640
rect 280154 267628 280160 267640
rect 209280 267600 280160 267628
rect 209280 267588 209286 267600
rect 280154 267588 280160 267600
rect 280212 267588 280218 267640
rect 369486 267588 369492 267640
rect 369544 267628 369550 267640
rect 452654 267628 452660 267640
rect 369544 267600 452660 267628
rect 369544 267588 369550 267600
rect 452654 267588 452660 267600
rect 452712 267588 452718 267640
rect 43806 267520 43812 267572
rect 43864 267560 43870 267572
rect 120074 267560 120080 267572
rect 43864 267532 120080 267560
rect 43864 267520 43870 267532
rect 120074 267520 120080 267532
rect 120132 267520 120138 267572
rect 203518 267520 203524 267572
rect 203576 267560 203582 267572
rect 267826 267560 267832 267572
rect 203576 267532 267832 267560
rect 203576 267520 203582 267532
rect 267826 267520 267832 267532
rect 267884 267520 267890 267572
rect 370406 267520 370412 267572
rect 370464 267560 370470 267572
rect 373166 267560 373172 267572
rect 370464 267532 373172 267560
rect 370464 267520 370470 267532
rect 373166 267520 373172 267532
rect 373224 267520 373230 267572
rect 376386 267520 376392 267572
rect 376444 267560 376450 267572
rect 458174 267560 458180 267572
rect 376444 267532 458180 267560
rect 376444 267520 376450 267532
rect 458174 267520 458180 267532
rect 458232 267520 458238 267572
rect 42334 267452 42340 267504
rect 42392 267492 42398 267504
rect 50982 267492 50988 267504
rect 42392 267464 50988 267492
rect 42392 267452 42398 267464
rect 50982 267452 50988 267464
rect 51040 267452 51046 267504
rect 55858 267452 55864 267504
rect 55916 267492 55922 267504
rect 129734 267492 129740 267504
rect 55916 267464 129740 267492
rect 55916 267452 55922 267464
rect 129734 267452 129740 267464
rect 129792 267452 129798 267504
rect 163498 267452 163504 267504
rect 163556 267492 163562 267504
rect 197630 267492 197636 267504
rect 163556 267464 197636 267492
rect 163556 267452 163562 267464
rect 197630 267452 197636 267464
rect 197688 267452 197694 267504
rect 200850 267452 200856 267504
rect 200908 267492 200914 267504
rect 264974 267492 264980 267504
rect 200908 267464 264980 267492
rect 200908 267452 200914 267464
rect 264974 267452 264980 267464
rect 265032 267452 265038 267504
rect 368198 267452 368204 267504
rect 368256 267492 368262 267504
rect 449894 267492 449900 267504
rect 368256 267464 449900 267492
rect 368256 267452 368262 267464
rect 449894 267452 449900 267464
rect 449952 267452 449958 267504
rect 53098 267384 53104 267436
rect 53156 267424 53162 267436
rect 117314 267424 117320 267436
rect 53156 267396 117320 267424
rect 53156 267384 53162 267396
rect 117314 267384 117320 267396
rect 117372 267384 117378 267436
rect 155954 267384 155960 267436
rect 156012 267424 156018 267436
rect 201862 267424 201868 267436
rect 156012 267396 201868 267424
rect 156012 267384 156018 267396
rect 201862 267384 201868 267396
rect 201920 267384 201926 267436
rect 202230 267384 202236 267436
rect 202288 267424 202294 267436
rect 263594 267424 263600 267436
rect 202288 267396 263600 267424
rect 202288 267384 202294 267396
rect 263594 267384 263600 267396
rect 263652 267384 263658 267436
rect 374914 267384 374920 267436
rect 374972 267424 374978 267436
rect 455782 267424 455788 267436
rect 374972 267396 455788 267424
rect 374972 267384 374978 267396
rect 455782 267384 455788 267396
rect 455840 267384 455846 267436
rect 53190 267316 53196 267368
rect 53248 267356 53254 267368
rect 115934 267356 115940 267368
rect 53248 267328 115940 267356
rect 53248 267316 53254 267328
rect 115934 267316 115940 267328
rect 115992 267316 115998 267368
rect 160922 267316 160928 267368
rect 160980 267356 160986 267368
rect 207106 267356 207112 267368
rect 160980 267328 207112 267356
rect 160980 267316 160986 267328
rect 207106 267316 207112 267328
rect 207164 267316 207170 267368
rect 214834 267316 214840 267368
rect 214892 267356 214898 267368
rect 273254 267356 273260 267368
rect 214892 267328 273260 267356
rect 214892 267316 214898 267328
rect 273254 267316 273260 267328
rect 273312 267316 273318 267368
rect 360194 267356 360200 267368
rect 354646 267328 360200 267356
rect 49142 267248 49148 267300
rect 49200 267288 49206 267300
rect 52914 267288 52920 267300
rect 49200 267260 52920 267288
rect 49200 267248 49206 267260
rect 52914 267248 52920 267260
rect 52972 267248 52978 267300
rect 53006 267248 53012 267300
rect 53064 267288 53070 267300
rect 113542 267288 113548 267300
rect 53064 267260 113548 267288
rect 53064 267248 53070 267260
rect 113542 267248 113548 267260
rect 113600 267248 113606 267300
rect 218974 267248 218980 267300
rect 219032 267288 219038 267300
rect 276014 267288 276020 267300
rect 219032 267260 276020 267288
rect 219032 267248 219038 267260
rect 276014 267248 276020 267260
rect 276072 267248 276078 267300
rect 343450 267248 343456 267300
rect 343508 267288 343514 267300
rect 354646 267288 354674 267328
rect 360194 267316 360200 267328
rect 360252 267316 360258 267368
rect 363874 267316 363880 267368
rect 363932 267356 363938 267368
rect 442994 267356 443000 267368
rect 363932 267328 443000 267356
rect 363932 267316 363938 267328
rect 442994 267316 443000 267328
rect 443052 267316 443058 267368
rect 357710 267288 357716 267300
rect 343508 267260 354674 267288
rect 356532 267260 357716 267288
rect 343508 267248 343514 267260
rect 51994 267180 52000 267232
rect 52052 267220 52058 267232
rect 107654 267220 107660 267232
rect 52052 267192 107660 267220
rect 52052 267180 52058 267192
rect 107654 267180 107660 267192
rect 107712 267180 107718 267232
rect 216122 267180 216128 267232
rect 216180 267220 216186 267232
rect 270494 267220 270500 267232
rect 216180 267192 270500 267220
rect 216180 267180 216186 267192
rect 270494 267180 270500 267192
rect 270552 267180 270558 267232
rect 278130 267180 278136 267232
rect 278188 267220 278194 267232
rect 356532 267220 356560 267260
rect 357710 267248 357716 267260
rect 357768 267248 357774 267300
rect 362586 267248 362592 267300
rect 362644 267288 362650 267300
rect 440234 267288 440240 267300
rect 362644 267260 440240 267288
rect 362644 267248 362650 267260
rect 440234 267248 440240 267260
rect 440292 267248 440298 267300
rect 278188 267192 356560 267220
rect 278188 267180 278194 267192
rect 356606 267180 356612 267232
rect 356664 267220 356670 267232
rect 357250 267220 357256 267232
rect 356664 267192 357256 267220
rect 356664 267180 356670 267192
rect 357250 267180 357256 267192
rect 357308 267180 357314 267232
rect 370866 267180 370872 267232
rect 370924 267220 370930 267232
rect 447134 267220 447140 267232
rect 370924 267192 447140 267220
rect 370924 267180 370930 267192
rect 447134 267180 447140 267192
rect 447192 267180 447198 267232
rect 503162 267180 503168 267232
rect 503220 267220 503226 267232
rect 517790 267220 517796 267232
rect 503220 267192 517796 267220
rect 503220 267180 503226 267192
rect 517790 267180 517796 267192
rect 517848 267180 517854 267232
rect 51810 267112 51816 267164
rect 51868 267152 51874 267164
rect 104894 267152 104900 267164
rect 51868 267124 104900 267152
rect 51868 267112 51874 267124
rect 104894 267112 104900 267124
rect 104952 267112 104958 267164
rect 205082 267112 205088 267164
rect 205140 267152 205146 267164
rect 258258 267152 258264 267164
rect 205140 267124 258264 267152
rect 205140 267112 205146 267124
rect 258258 267112 258264 267124
rect 258316 267112 258322 267164
rect 279142 267112 279148 267164
rect 279200 267152 279206 267164
rect 358814 267152 358820 267164
rect 279200 267124 358820 267152
rect 279200 267112 279206 267124
rect 358814 267112 358820 267124
rect 358872 267112 358878 267164
rect 372338 267112 372344 267164
rect 372396 267152 372402 267164
rect 445754 267152 445760 267164
rect 372396 267124 445760 267152
rect 372396 267112 372402 267124
rect 445754 267112 445760 267124
rect 445812 267112 445818 267164
rect 52086 267044 52092 267096
rect 52144 267084 52150 267096
rect 103514 267084 103520 267096
rect 52144 267056 103520 267084
rect 52144 267044 52150 267056
rect 103514 267044 103520 267056
rect 103572 267044 103578 267096
rect 198274 267044 198280 267096
rect 198332 267084 198338 267096
rect 202874 267084 202880 267096
rect 198332 267056 202880 267084
rect 198332 267044 198338 267056
rect 202874 267044 202880 267056
rect 202932 267044 202938 267096
rect 210878 267044 210884 267096
rect 210936 267084 210942 267096
rect 260834 267084 260840 267096
rect 210936 267056 260840 267084
rect 210936 267044 210942 267056
rect 260834 267044 260840 267056
rect 260892 267044 260898 267096
rect 277026 267044 277032 267096
rect 277084 267084 277090 267096
rect 356606 267084 356612 267096
rect 277084 267056 356612 267084
rect 277084 267044 277090 267056
rect 356606 267044 356612 267056
rect 356664 267044 356670 267096
rect 366818 267044 366824 267096
rect 366876 267084 366882 267096
rect 437474 267084 437480 267096
rect 366876 267056 437480 267084
rect 366876 267044 366882 267056
rect 437474 267044 437480 267056
rect 437532 267044 437538 267096
rect 503530 267044 503536 267096
rect 503588 267084 503594 267096
rect 517882 267084 517888 267096
rect 503588 267056 517888 267084
rect 503588 267044 503594 267056
rect 517882 267044 517888 267056
rect 517940 267044 517946 267096
rect 50246 266976 50252 267028
rect 50304 267016 50310 267028
rect 100754 267016 100760 267028
rect 50304 266988 100760 267016
rect 50304 266976 50310 266988
rect 100754 266976 100760 266988
rect 100812 266976 100818 267028
rect 183278 266976 183284 267028
rect 183336 267016 183342 267028
rect 200114 267016 200120 267028
rect 183336 266988 200120 267016
rect 183336 266976 183342 266988
rect 200114 266976 200120 266988
rect 200172 267016 200178 267028
rect 201034 267016 201040 267028
rect 200172 266988 201040 267016
rect 200172 266976 200178 266988
rect 201034 266976 201040 266988
rect 201092 266976 201098 267028
rect 215018 266976 215024 267028
rect 215076 267016 215082 267028
rect 273254 267016 273260 267028
rect 215076 266988 273260 267016
rect 215076 266976 215082 266988
rect 273254 266976 273260 266988
rect 273312 266976 273318 267028
rect 275922 266976 275928 267028
rect 275980 267016 275986 267028
rect 356974 267016 356980 267028
rect 275980 266988 356980 267016
rect 275980 266976 275986 266988
rect 356974 266976 356980 266988
rect 357032 266976 357038 267028
rect 365438 266976 365444 267028
rect 365496 267016 365502 267028
rect 433334 267016 433340 267028
rect 365496 266988 433340 267016
rect 365496 266976 365502 266988
rect 433334 266976 433340 266988
rect 433392 266976 433398 267028
rect 440050 266976 440056 267028
rect 440108 267016 440114 267028
rect 516594 267016 516600 267028
rect 440108 266988 516600 267016
rect 440108 266976 440114 266988
rect 516594 266976 516600 266988
rect 516652 266976 516658 267028
rect 54754 266908 54760 266960
rect 54812 266948 54818 266960
rect 88334 266948 88340 266960
rect 54812 266920 88340 266948
rect 54812 266908 54818 266920
rect 88334 266908 88340 266920
rect 88392 266908 88398 266960
rect 206554 266908 206560 266960
rect 206612 266948 206618 266960
rect 255314 266948 255320 266960
rect 206612 266920 255320 266948
rect 206612 266908 206618 266920
rect 255314 266908 255320 266920
rect 255372 266908 255378 266960
rect 358446 266908 358452 266960
rect 358504 266948 358510 266960
rect 418154 266948 418160 266960
rect 358504 266920 418160 266948
rect 358504 266908 358510 266920
rect 418154 266908 418160 266920
rect 418212 266908 418218 266960
rect 48038 266840 48044 266892
rect 48096 266880 48102 266892
rect 78674 266880 78680 266892
rect 48096 266852 78680 266880
rect 48096 266840 48102 266852
rect 78674 266840 78680 266852
rect 78732 266840 78738 266892
rect 207842 266840 207848 266892
rect 207900 266880 207906 266892
rect 252554 266880 252560 266892
rect 207900 266852 252560 266880
rect 207900 266840 207906 266852
rect 252554 266840 252560 266852
rect 252612 266840 252618 266892
rect 376202 266840 376208 266892
rect 376260 266880 376266 266892
rect 412910 266880 412916 266892
rect 376260 266852 412916 266880
rect 376260 266840 376266 266852
rect 412910 266840 412916 266852
rect 412968 266840 412974 266892
rect 47762 266772 47768 266824
rect 47820 266812 47826 266824
rect 77294 266812 77300 266824
rect 47820 266784 77300 266812
rect 47820 266772 47826 266784
rect 77294 266772 77300 266784
rect 77352 266772 77358 266824
rect 216214 266772 216220 266824
rect 216272 266812 216278 266824
rect 247034 266812 247040 266824
rect 216272 266784 247040 266812
rect 216272 266772 216278 266784
rect 247034 266772 247040 266784
rect 247092 266772 247098 266824
rect 373626 266772 373632 266824
rect 373684 266812 373690 266824
rect 409874 266812 409880 266824
rect 373684 266784 409880 266812
rect 373684 266772 373690 266784
rect 409874 266772 409880 266784
rect 409932 266772 409938 266824
rect 213362 266704 213368 266756
rect 213420 266744 213426 266756
rect 285674 266744 285680 266756
rect 213420 266716 285680 266744
rect 213420 266704 213426 266716
rect 285674 266704 285680 266716
rect 285732 266704 285738 266756
rect 47670 266500 47676 266552
rect 47728 266540 47734 266552
rect 48038 266540 48044 266552
rect 47728 266512 48044 266540
rect 47728 266500 47734 266512
rect 48038 266500 48044 266512
rect 48096 266500 48102 266552
rect 357066 266472 357072 266484
rect 354646 266444 357072 266472
rect 50338 266364 50344 266416
rect 50396 266404 50402 266416
rect 50982 266404 50988 266416
rect 50396 266376 50988 266404
rect 50396 266364 50402 266376
rect 50982 266364 50988 266376
rect 51040 266364 51046 266416
rect 80054 266364 80060 266416
rect 80112 266404 80118 266416
rect 104894 266404 104900 266416
rect 80112 266376 104900 266404
rect 80112 266364 80118 266376
rect 104894 266364 104900 266376
rect 104952 266364 104958 266416
rect 183462 266364 183468 266416
rect 183520 266404 183526 266416
rect 197446 266404 197452 266416
rect 183520 266376 197452 266404
rect 183520 266364 183526 266376
rect 197446 266364 197452 266376
rect 197504 266404 197510 266416
rect 198274 266404 198280 266416
rect 197504 266376 198280 266404
rect 197504 266364 197510 266376
rect 198274 266364 198280 266376
rect 198332 266364 198338 266416
rect 343450 266364 343456 266416
rect 343508 266404 343514 266416
rect 354646 266404 354674 266444
rect 357066 266432 357072 266444
rect 357124 266472 357130 266484
rect 363046 266472 363052 266484
rect 357124 266444 363052 266472
rect 357124 266432 357130 266444
rect 363046 266432 363052 266444
rect 363104 266432 363110 266484
rect 343508 266376 354674 266404
rect 343508 266364 343514 266376
rect 356790 266364 356796 266416
rect 356848 266404 356854 266416
rect 356974 266404 356980 266416
rect 356848 266376 356980 266404
rect 356848 266364 356854 266376
rect 356974 266364 356980 266376
rect 357032 266364 357038 266416
rect 421558 266364 421564 266416
rect 421616 266404 421622 266416
rect 437474 266404 437480 266416
rect 421616 266376 437480 266404
rect 421616 266364 421622 266376
rect 437474 266364 437480 266376
rect 437532 266364 437538 266416
rect 517790 266364 517796 266416
rect 517848 266404 517854 266416
rect 517974 266404 517980 266416
rect 517848 266376 517980 266404
rect 517848 266364 517854 266376
rect 517974 266364 517980 266376
rect 518032 266364 518038 266416
rect 55766 266296 55772 266348
rect 55824 266336 55830 266348
rect 56870 266336 56876 266348
rect 55824 266308 56876 266336
rect 55824 266296 55830 266308
rect 56870 266296 56876 266308
rect 56928 266296 56934 266348
rect 57974 266296 57980 266348
rect 58032 266336 58038 266348
rect 58618 266336 58624 266348
rect 58032 266308 58624 266336
rect 58032 266296 58038 266308
rect 58618 266296 58624 266308
rect 58676 266336 58682 266348
rect 92382 266336 92388 266348
rect 58676 266308 92388 266336
rect 58676 266296 58682 266308
rect 92382 266296 92388 266308
rect 92440 266296 92446 266348
rect 109954 266296 109960 266348
rect 110012 266336 110018 266348
rect 196802 266336 196808 266348
rect 110012 266308 196808 266336
rect 110012 266296 110018 266308
rect 196802 266296 196808 266308
rect 196860 266296 196866 266348
rect 216214 266296 216220 266348
rect 216272 266336 216278 266348
rect 262214 266336 262220 266348
rect 216272 266308 262220 266336
rect 216272 266296 216278 266308
rect 262214 266296 262220 266308
rect 262272 266296 262278 266348
rect 379974 266296 379980 266348
rect 380032 266336 380038 266348
rect 396074 266336 396080 266348
rect 380032 266308 396080 266336
rect 380032 266296 380038 266308
rect 396074 266296 396080 266308
rect 396132 266296 396138 266348
rect 54570 266228 54576 266280
rect 54628 266268 54634 266280
rect 55858 266268 55864 266280
rect 54628 266240 55864 266268
rect 54628 266228 54634 266240
rect 55858 266228 55864 266240
rect 55916 266228 55922 266280
rect 56888 266268 56916 266296
rect 117314 266268 117320 266280
rect 56888 266240 117320 266268
rect 117314 266228 117320 266240
rect 117372 266228 117378 266280
rect 213730 266228 213736 266280
rect 213788 266268 213794 266280
rect 247034 266268 247040 266280
rect 213788 266240 247040 266268
rect 213788 266228 213794 266240
rect 247034 266228 247040 266240
rect 247092 266228 247098 266280
rect 379238 266228 379244 266280
rect 379296 266268 379302 266280
rect 411254 266268 411260 266280
rect 379296 266240 411260 266268
rect 379296 266228 379302 266240
rect 411254 266228 411260 266240
rect 411312 266228 411318 266280
rect 51902 266160 51908 266212
rect 51960 266200 51966 266212
rect 57974 266200 57980 266212
rect 51960 266172 57980 266200
rect 51960 266160 51966 266172
rect 57974 266160 57980 266172
rect 58032 266160 58038 266212
rect 216950 266160 216956 266212
rect 217008 266200 217014 266212
rect 219158 266200 219164 266212
rect 217008 266172 219164 266200
rect 217008 266160 217014 266172
rect 219158 266160 219164 266172
rect 219216 266200 219222 266212
rect 251266 266200 251272 266212
rect 219216 266172 251272 266200
rect 219216 266160 219222 266172
rect 251266 266160 251272 266172
rect 251324 266160 251330 266212
rect 373902 266160 373908 266212
rect 373960 266200 373966 266212
rect 376478 266200 376484 266212
rect 373960 266172 376484 266200
rect 373960 266160 373966 266172
rect 376478 266160 376484 266172
rect 376536 266200 376542 266212
rect 407114 266200 407120 266212
rect 376536 266172 407120 266200
rect 376536 266160 376542 266172
rect 407114 266160 407120 266172
rect 407172 266160 407178 266212
rect 62206 266092 62212 266144
rect 62264 266132 62270 266144
rect 92474 266132 92480 266144
rect 62264 266104 92480 266132
rect 62264 266092 62270 266104
rect 92474 266092 92480 266104
rect 92532 266092 92538 266144
rect 219250 266092 219256 266144
rect 219308 266132 219314 266144
rect 219618 266132 219624 266144
rect 219308 266104 219624 266132
rect 219308 266092 219314 266104
rect 219618 266092 219624 266104
rect 219676 266132 219682 266144
rect 251174 266132 251180 266144
rect 219676 266104 251180 266132
rect 219676 266092 219682 266104
rect 251174 266092 251180 266104
rect 251232 266092 251238 266144
rect 378042 266092 378048 266144
rect 378100 266132 378106 266144
rect 408494 266132 408500 266144
rect 378100 266104 408500 266132
rect 378100 266092 378106 266104
rect 408494 266092 408500 266104
rect 408552 266092 408558 266144
rect 54478 266024 54484 266076
rect 54536 266064 54542 266076
rect 84194 266064 84200 266076
rect 54536 266036 84200 266064
rect 54536 266024 54542 266036
rect 84194 266024 84200 266036
rect 84252 266024 84258 266076
rect 215662 266024 215668 266076
rect 215720 266064 215726 266076
rect 245654 266064 245660 266076
rect 215720 266036 245660 266064
rect 215720 266024 215726 266036
rect 245654 266024 245660 266036
rect 245712 266024 245718 266076
rect 379882 266024 379888 266076
rect 379940 266064 379946 266076
rect 409874 266064 409880 266076
rect 379940 266036 409880 266064
rect 379940 266024 379946 266036
rect 409874 266024 409880 266036
rect 409932 266024 409938 266076
rect 57974 265956 57980 266008
rect 58032 265996 58038 266008
rect 89714 265996 89720 266008
rect 58032 265968 89720 265996
rect 58032 265956 58038 265968
rect 89714 265956 89720 265968
rect 89772 265956 89778 266008
rect 196710 265956 196716 266008
rect 196768 265996 196774 266008
rect 197538 265996 197544 266008
rect 196768 265968 197544 265996
rect 196768 265956 196774 265968
rect 197538 265956 197544 265968
rect 197596 265956 197602 266008
rect 215110 265956 215116 266008
rect 215168 265996 215174 266008
rect 216122 265996 216128 266008
rect 215168 265968 216128 265996
rect 215168 265956 215174 265968
rect 216122 265956 216128 265968
rect 216180 265956 216186 266008
rect 217962 265956 217968 266008
rect 218020 265996 218026 266008
rect 219894 265996 219900 266008
rect 218020 265968 219900 265996
rect 218020 265956 218026 265968
rect 219894 265956 219900 265968
rect 219952 265996 219958 266008
rect 249794 265996 249800 266008
rect 219952 265968 249800 265996
rect 219952 265956 219958 265968
rect 249794 265956 249800 265968
rect 249852 265956 249858 266008
rect 375190 265956 375196 266008
rect 375248 265996 375254 266008
rect 400214 265996 400220 266008
rect 375248 265968 400220 265996
rect 375248 265956 375254 265968
rect 400214 265956 400220 265968
rect 400272 265956 400278 266008
rect 54570 265888 54576 265940
rect 54628 265928 54634 265940
rect 85574 265928 85580 265940
rect 54628 265900 85580 265928
rect 54628 265888 54634 265900
rect 85574 265888 85580 265900
rect 85632 265888 85638 265940
rect 219158 265888 219164 265940
rect 219216 265928 219222 265940
rect 219526 265928 219532 265940
rect 219216 265900 219532 265928
rect 219216 265888 219222 265900
rect 219526 265888 219532 265900
rect 219584 265928 219590 265940
rect 248506 265928 248512 265940
rect 219584 265900 248512 265928
rect 219584 265888 219590 265900
rect 248506 265888 248512 265900
rect 248564 265888 248570 265940
rect 370222 265888 370228 265940
rect 370280 265928 370286 265940
rect 372982 265928 372988 265940
rect 370280 265900 372988 265928
rect 370280 265888 370286 265900
rect 372982 265888 372988 265900
rect 373040 265928 373046 265940
rect 398834 265928 398840 265940
rect 373040 265900 398840 265928
rect 373040 265888 373046 265900
rect 398834 265888 398840 265900
rect 398892 265888 398898 265940
rect 51994 265860 52000 265872
rect 51046 265832 52000 265860
rect 50430 265684 50436 265736
rect 50488 265724 50494 265736
rect 51046 265724 51074 265832
rect 51994 265820 52000 265832
rect 52052 265860 52058 265872
rect 85390 265860 85396 265872
rect 52052 265832 85396 265860
rect 52052 265820 52058 265832
rect 85390 265820 85396 265832
rect 85448 265820 85454 265872
rect 218606 265820 218612 265872
rect 218664 265860 218670 265872
rect 219894 265860 219900 265872
rect 218664 265832 219900 265860
rect 218664 265820 218670 265832
rect 219894 265820 219900 265832
rect 219952 265860 219958 265872
rect 252554 265860 252560 265872
rect 219952 265832 252560 265860
rect 219952 265820 219958 265832
rect 252554 265820 252560 265832
rect 252612 265820 252618 265872
rect 379698 265820 379704 265872
rect 379756 265860 379762 265872
rect 404354 265860 404360 265872
rect 379756 265832 404360 265860
rect 379756 265820 379762 265832
rect 404354 265820 404360 265832
rect 404412 265820 404418 265872
rect 55858 265752 55864 265804
rect 55916 265792 55922 265804
rect 88334 265792 88340 265804
rect 55916 265764 88340 265792
rect 55916 265752 55922 265764
rect 88334 265752 88340 265764
rect 88392 265752 88398 265804
rect 217134 265752 217140 265804
rect 217192 265792 217198 265804
rect 218974 265792 218980 265804
rect 217192 265764 218980 265792
rect 217192 265752 217198 265764
rect 218974 265752 218980 265764
rect 219032 265792 219038 265804
rect 263594 265792 263600 265804
rect 219032 265764 263600 265792
rect 219032 265752 219038 265764
rect 263594 265752 263600 265764
rect 263652 265752 263658 265804
rect 371050 265752 371056 265804
rect 371108 265792 371114 265804
rect 372430 265792 372436 265804
rect 371108 265764 372436 265792
rect 371108 265752 371114 265764
rect 372430 265752 372436 265764
rect 372488 265792 372494 265804
rect 398190 265792 398196 265804
rect 372488 265764 398196 265792
rect 372488 265752 372494 265764
rect 398190 265752 398196 265764
rect 398248 265752 398254 265804
rect 50488 265696 51074 265724
rect 50488 265684 50494 265696
rect 53098 265684 53104 265736
rect 53156 265724 53162 265736
rect 86954 265724 86960 265736
rect 53156 265696 86960 265724
rect 53156 265684 53162 265696
rect 86954 265684 86960 265696
rect 87012 265684 87018 265736
rect 88242 265684 88248 265736
rect 88300 265724 88306 265736
rect 113726 265724 113732 265736
rect 88300 265696 113732 265724
rect 88300 265684 88306 265696
rect 113726 265684 113732 265696
rect 113784 265684 113790 265736
rect 215478 265684 215484 265736
rect 215536 265724 215542 265736
rect 216214 265724 216220 265736
rect 215536 265696 216220 265724
rect 215536 265684 215542 265696
rect 216214 265684 216220 265696
rect 216272 265684 216278 265736
rect 219342 265684 219348 265736
rect 219400 265724 219406 265736
rect 219618 265724 219624 265736
rect 219400 265696 219624 265724
rect 219400 265684 219406 265696
rect 219618 265684 219624 265696
rect 219676 265724 219682 265736
rect 265158 265724 265164 265736
rect 219676 265696 265164 265724
rect 219676 265684 219682 265696
rect 265158 265684 265164 265696
rect 265216 265684 265222 265736
rect 376570 265684 376576 265736
rect 376628 265724 376634 265736
rect 403158 265724 403164 265736
rect 376628 265696 403164 265724
rect 376628 265684 376634 265696
rect 403158 265684 403164 265696
rect 403216 265684 403222 265736
rect 59722 265616 59728 265668
rect 59780 265656 59786 265668
rect 107654 265656 107660 265668
rect 59780 265628 107660 265656
rect 59780 265616 59786 265628
rect 107654 265616 107660 265628
rect 107712 265616 107718 265668
rect 114370 265616 114376 265668
rect 114428 265656 114434 265668
rect 196710 265656 196716 265668
rect 114428 265628 196716 265656
rect 114428 265616 114434 265628
rect 196710 265616 196716 265628
rect 196768 265616 196774 265668
rect 216582 265616 216588 265668
rect 216640 265656 216646 265668
rect 218606 265656 218612 265668
rect 216640 265628 218612 265656
rect 216640 265616 216646 265628
rect 218606 265616 218612 265628
rect 218664 265656 218670 265668
rect 266354 265656 266360 265668
rect 218664 265628 266360 265656
rect 218664 265616 218670 265628
rect 266354 265616 266360 265628
rect 266412 265616 266418 265668
rect 371142 265616 371148 265668
rect 371200 265656 371206 265668
rect 372338 265656 372344 265668
rect 371200 265628 372344 265656
rect 371200 265616 371206 265628
rect 372338 265616 372344 265628
rect 372396 265656 372402 265668
rect 401686 265656 401692 265668
rect 372396 265628 401692 265656
rect 372396 265616 372402 265628
rect 401686 265616 401692 265628
rect 401744 265616 401750 265668
rect 216122 265548 216128 265600
rect 216180 265588 216186 265600
rect 244274 265588 244280 265600
rect 216180 265560 244280 265588
rect 216180 265548 216186 265560
rect 244274 265548 244280 265560
rect 244332 265548 244338 265600
rect 377950 265548 377956 265600
rect 378008 265588 378014 265600
rect 411346 265588 411352 265600
rect 378008 265560 411352 265588
rect 378008 265548 378014 265560
rect 411346 265548 411352 265560
rect 411404 265548 411410 265600
rect 375282 265412 375288 265464
rect 375340 265452 375346 265464
rect 376570 265452 376576 265464
rect 375340 265424 376576 265452
rect 375340 265412 375346 265424
rect 376570 265412 376576 265424
rect 376628 265412 376634 265464
rect 376386 265276 376392 265328
rect 376444 265316 376450 265328
rect 376444 265288 383654 265316
rect 376444 265276 376450 265288
rect 374086 265208 374092 265260
rect 374144 265248 374150 265260
rect 379974 265248 379980 265260
rect 374144 265220 379980 265248
rect 374144 265208 374150 265220
rect 379974 265208 379980 265220
rect 380032 265208 380038 265260
rect 375926 265140 375932 265192
rect 375984 265180 375990 265192
rect 375984 265152 380020 265180
rect 375984 265140 375990 265152
rect 213638 265072 213644 265124
rect 213696 265112 213702 265124
rect 215662 265112 215668 265124
rect 213696 265084 215668 265112
rect 213696 265072 213702 265084
rect 215662 265072 215668 265084
rect 215720 265072 215726 265124
rect 214374 265004 214380 265056
rect 214432 265044 214438 265056
rect 230382 265044 230388 265056
rect 214432 265016 230388 265044
rect 214432 265004 214438 265016
rect 230382 265004 230388 265016
rect 230440 265004 230446 265056
rect 378502 265004 378508 265056
rect 378560 265044 378566 265056
rect 379698 265044 379704 265056
rect 378560 265016 379704 265044
rect 378560 265004 378566 265016
rect 379698 265004 379704 265016
rect 379756 265004 379762 265056
rect 47946 264936 47952 264988
rect 48004 264976 48010 264988
rect 48004 264948 51074 264976
rect 48004 264936 48010 264948
rect 51046 264908 51074 264948
rect 214282 264936 214288 264988
rect 214340 264976 214346 264988
rect 215754 264976 215760 264988
rect 214340 264948 215760 264976
rect 214340 264936 214346 264948
rect 215754 264936 215760 264948
rect 215812 264976 215818 264988
rect 233142 264976 233148 264988
rect 215812 264948 233148 264976
rect 215812 264936 215818 264948
rect 233142 264936 233148 264948
rect 233200 264936 233206 264988
rect 376846 264936 376852 264988
rect 376904 264976 376910 264988
rect 378042 264976 378048 264988
rect 376904 264948 378048 264976
rect 376904 264936 376910 264948
rect 378042 264936 378048 264948
rect 378100 264936 378106 264988
rect 378594 264936 378600 264988
rect 378652 264976 378658 264988
rect 379882 264976 379888 264988
rect 378652 264948 379888 264976
rect 378652 264936 378658 264948
rect 379882 264936 379888 264948
rect 379940 264936 379946 264988
rect 379992 264976 380020 265152
rect 383626 265044 383654 265288
rect 390554 265044 390560 265056
rect 383626 265016 390560 265044
rect 390554 265004 390560 265016
rect 390612 265004 390618 265056
rect 391934 264976 391940 264988
rect 379992 264948 391940 264976
rect 391934 264936 391940 264948
rect 391992 264936 391998 264988
rect 51626 264908 51632 264920
rect 51046 264880 51632 264908
rect 51626 264868 51632 264880
rect 51684 264908 51690 264920
rect 88242 264908 88248 264920
rect 51684 264880 88248 264908
rect 51684 264868 51690 264880
rect 88242 264868 88248 264880
rect 88300 264868 88306 264920
rect 212166 264868 212172 264920
rect 212224 264908 212230 264920
rect 273162 264908 273168 264920
rect 212224 264880 273168 264908
rect 212224 264868 212230 264880
rect 273162 264868 273168 264880
rect 273220 264868 273226 264920
rect 388438 264868 388444 264920
rect 388496 264908 388502 264920
rect 420914 264908 420920 264920
rect 388496 264880 420920 264908
rect 388496 264868 388502 264880
rect 420914 264868 420920 264880
rect 420972 264868 420978 264920
rect 43714 264800 43720 264852
rect 43772 264840 43778 264852
rect 59722 264840 59728 264852
rect 43772 264812 59728 264840
rect 43772 264800 43778 264812
rect 59722 264800 59728 264812
rect 59780 264800 59786 264852
rect 211706 264800 211712 264852
rect 211764 264840 211770 264852
rect 270494 264840 270500 264852
rect 211764 264812 270500 264840
rect 211764 264800 211770 264812
rect 270494 264800 270500 264812
rect 270552 264800 270558 264852
rect 389174 264800 389180 264852
rect 389232 264840 389238 264852
rect 419534 264840 419540 264852
rect 389232 264812 419540 264840
rect 389232 264800 389238 264812
rect 419534 264800 419540 264812
rect 419592 264800 419598 264852
rect 49234 264732 49240 264784
rect 49292 264772 49298 264784
rect 62206 264772 62212 264784
rect 49292 264744 62212 264772
rect 49292 264732 49298 264744
rect 62206 264732 62212 264744
rect 62264 264732 62270 264784
rect 219802 264732 219808 264784
rect 219860 264772 219866 264784
rect 253934 264772 253940 264784
rect 219860 264744 253940 264772
rect 219860 264732 219866 264744
rect 253934 264732 253940 264744
rect 253992 264732 253998 264784
rect 378686 264732 378692 264784
rect 378744 264772 378750 264784
rect 405734 264772 405740 264784
rect 378744 264744 405740 264772
rect 378744 264732 378750 264744
rect 405734 264732 405740 264744
rect 405792 264732 405798 264784
rect 48222 264664 48228 264716
rect 48280 264704 48286 264716
rect 57974 264704 57980 264716
rect 48280 264676 57980 264704
rect 48280 264664 48286 264676
rect 57974 264664 57980 264676
rect 58032 264664 58038 264716
rect 230382 264664 230388 264716
rect 230440 264704 230446 264716
rect 259546 264704 259552 264716
rect 230440 264676 259552 264704
rect 230440 264664 230446 264676
rect 259546 264664 259552 264676
rect 259604 264664 259610 264716
rect 390554 264664 390560 264716
rect 390612 264704 390618 264716
rect 418246 264704 418252 264716
rect 390612 264676 418252 264704
rect 390612 264664 390618 264676
rect 418246 264664 418252 264676
rect 418304 264664 418310 264716
rect 46750 264596 46756 264648
rect 46808 264636 46814 264648
rect 54478 264636 54484 264648
rect 46808 264608 54484 264636
rect 46808 264596 46814 264608
rect 54478 264596 54484 264608
rect 54536 264596 54542 264648
rect 233142 264596 233148 264648
rect 233200 264636 233206 264648
rect 259454 264636 259460 264648
rect 233200 264608 259460 264636
rect 233200 264596 233206 264608
rect 259454 264596 259460 264608
rect 259512 264596 259518 264648
rect 391934 264596 391940 264648
rect 391992 264636 391998 264648
rect 418154 264636 418160 264648
rect 391992 264608 418160 264636
rect 391992 264596 391998 264608
rect 418154 264596 418160 264608
rect 418212 264596 418218 264648
rect 46658 264528 46664 264580
rect 46716 264568 46722 264580
rect 53098 264568 53104 264580
rect 46716 264540 53104 264568
rect 46716 264528 46722 264540
rect 53098 264528 53104 264540
rect 53156 264528 53162 264580
rect 215110 264528 215116 264580
rect 215168 264568 215174 264580
rect 219066 264568 219072 264580
rect 215168 264540 219072 264568
rect 215168 264528 215174 264540
rect 219066 264528 219072 264540
rect 219124 264568 219130 264580
rect 244366 264568 244372 264580
rect 219124 264540 244372 264568
rect 219124 264528 219130 264540
rect 244366 264528 244372 264540
rect 244424 264528 244430 264580
rect 46566 264460 46572 264512
rect 46624 264500 46630 264512
rect 54570 264500 54576 264512
rect 46624 264472 54576 264500
rect 46624 264460 46630 264472
rect 54570 264460 54576 264472
rect 54628 264460 54634 264512
rect 210234 264256 210240 264308
rect 210292 264296 210298 264308
rect 217134 264296 217140 264308
rect 210292 264268 217140 264296
rect 210292 264256 210298 264268
rect 217134 264256 217140 264268
rect 217192 264296 217198 264308
rect 256694 264296 256700 264308
rect 217192 264268 256700 264296
rect 217192 264256 217198 264268
rect 256694 264256 256700 264268
rect 256752 264256 256758 264308
rect 57790 264188 57796 264240
rect 57848 264228 57854 264240
rect 80054 264228 80060 264240
rect 57848 264200 80060 264228
rect 57848 264188 57854 264200
rect 80054 264188 80060 264200
rect 80112 264188 80118 264240
rect 213546 264188 213552 264240
rect 213604 264228 213610 264240
rect 269114 264228 269120 264240
rect 213604 264200 269120 264228
rect 213604 264188 213610 264200
rect 269114 264188 269120 264200
rect 269172 264188 269178 264240
rect 379330 264188 379336 264240
rect 379388 264228 379394 264240
rect 413002 264228 413008 264240
rect 379388 264200 413008 264228
rect 379388 264188 379394 264200
rect 413002 264188 413008 264200
rect 413060 264188 413066 264240
rect 210326 263644 210332 263696
rect 210384 263684 210390 263696
rect 213546 263684 213552 263696
rect 210384 263656 213552 263684
rect 210384 263644 210390 263656
rect 213546 263644 213552 263656
rect 213604 263644 213610 263696
rect 211706 263576 211712 263628
rect 211764 263616 211770 263628
rect 212074 263616 212080 263628
rect 211764 263588 212080 263616
rect 211764 263576 211770 263588
rect 212074 263576 212080 263588
rect 212132 263576 212138 263628
rect 376478 263576 376484 263628
rect 376536 263616 376542 263628
rect 378686 263616 378692 263628
rect 376536 263588 378692 263616
rect 376536 263576 376542 263588
rect 378686 263576 378692 263588
rect 378744 263576 378750 263628
rect 379330 263576 379336 263628
rect 379388 263616 379394 263628
rect 379882 263616 379888 263628
rect 379388 263588 379888 263616
rect 379388 263576 379394 263588
rect 379882 263576 379888 263588
rect 379940 263576 379946 263628
rect 42426 263508 42432 263560
rect 42484 263548 42490 263560
rect 57238 263548 57244 263560
rect 42484 263520 57244 263548
rect 42484 263508 42490 263520
rect 57238 263508 57244 263520
rect 57296 263548 57302 263560
rect 57790 263548 57796 263560
rect 57296 263520 57796 263548
rect 57296 263508 57302 263520
rect 57790 263508 57796 263520
rect 57848 263508 57854 263560
rect 375098 263508 375104 263560
rect 375156 263548 375162 263560
rect 436094 263548 436100 263560
rect 375156 263520 436100 263548
rect 375156 263508 375162 263520
rect 436094 263508 436100 263520
rect 436152 263508 436158 263560
rect 214374 262964 214380 263016
rect 214432 262964 214438 263016
rect 214392 262732 214420 262964
rect 378962 262828 378968 262880
rect 379020 262868 379026 262880
rect 426434 262868 426440 262880
rect 379020 262840 426440 262868
rect 379020 262828 379026 262840
rect 426434 262828 426440 262840
rect 426492 262828 426498 262880
rect 214466 262732 214472 262744
rect 214392 262704 214472 262732
rect 214466 262692 214472 262704
rect 214524 262692 214530 262744
rect 369670 262148 369676 262200
rect 369728 262188 369734 262200
rect 378962 262188 378968 262200
rect 369728 262160 378968 262188
rect 369728 262148 369734 262160
rect 378962 262148 378968 262160
rect 379020 262148 379026 262200
rect 220814 251132 220820 251184
rect 220872 251172 220878 251184
rect 221366 251172 221372 251184
rect 220872 251144 221372 251172
rect 220872 251132 220878 251144
rect 221366 251132 221372 251144
rect 221424 251172 221430 251184
rect 266446 251172 266452 251184
rect 221424 251144 266452 251172
rect 221424 251132 221430 251144
rect 266446 251132 266452 251144
rect 266504 251132 266510 251184
rect 369762 251132 369768 251184
rect 369820 251172 369826 251184
rect 370406 251172 370412 251184
rect 369820 251144 370412 251172
rect 369820 251132 369826 251144
rect 370406 251132 370412 251144
rect 370464 251132 370470 251184
rect 374546 251132 374552 251184
rect 374604 251172 374610 251184
rect 395338 251172 395344 251184
rect 374604 251144 395344 251172
rect 374604 251132 374610 251144
rect 395338 251132 395344 251144
rect 395396 251132 395402 251184
rect 197354 251064 197360 251116
rect 197412 251104 197418 251116
rect 197630 251104 197636 251116
rect 197412 251076 197636 251104
rect 197412 251064 197418 251076
rect 197630 251064 197636 251076
rect 197688 251064 197694 251116
rect 368382 251064 368388 251116
rect 368440 251104 368446 251116
rect 370958 251104 370964 251116
rect 368440 251076 370964 251104
rect 368440 251064 368446 251076
rect 370958 251064 370964 251076
rect 371016 251064 371022 251116
rect 379146 251064 379152 251116
rect 379204 251104 379210 251116
rect 379422 251104 379428 251116
rect 379204 251076 379428 251104
rect 379204 251064 379210 251076
rect 379422 251064 379428 251076
rect 379480 251104 379486 251116
rect 396718 251104 396724 251116
rect 379480 251076 396724 251104
rect 379480 251064 379486 251076
rect 396718 251064 396724 251076
rect 396776 251064 396782 251116
rect 368290 250996 368296 251048
rect 368348 251036 368354 251048
rect 370866 251036 370872 251048
rect 368348 251008 370872 251036
rect 368348 250996 368354 251008
rect 370866 250996 370872 251008
rect 370924 250996 370930 251048
rect 500034 250656 500040 250708
rect 500092 250696 500098 250708
rect 517606 250696 517612 250708
rect 500092 250668 517612 250696
rect 500092 250656 500098 250668
rect 517606 250656 517612 250668
rect 517664 250656 517670 250708
rect 204162 250588 204168 250640
rect 204220 250628 204226 250640
rect 204220 250600 216076 250628
rect 204220 250588 204226 250600
rect 58710 250520 58716 250572
rect 58768 250560 58774 250572
rect 79318 250560 79324 250572
rect 58768 250532 79324 250560
rect 58768 250520 58774 250532
rect 79318 250520 79324 250532
rect 79376 250520 79382 250572
rect 85850 250520 85856 250572
rect 85908 250560 85914 250572
rect 106918 250560 106924 250572
rect 85908 250532 106924 250560
rect 85908 250520 85914 250532
rect 106918 250520 106924 250532
rect 106976 250520 106982 250572
rect 179782 250520 179788 250572
rect 179840 250560 179846 250572
rect 197630 250560 197636 250572
rect 179840 250532 197636 250560
rect 179840 250520 179846 250532
rect 197630 250520 197636 250532
rect 197688 250520 197694 250572
rect 58618 250452 58624 250504
rect 58676 250492 58682 250504
rect 106274 250492 106280 250504
rect 58676 250464 106280 250492
rect 58676 250452 58682 250464
rect 106274 250452 106280 250464
rect 106332 250452 106338 250504
rect 179322 250452 179328 250504
rect 179380 250492 179386 250504
rect 197538 250492 197544 250504
rect 179380 250464 197544 250492
rect 179380 250452 179386 250464
rect 197538 250452 197544 250464
rect 197596 250452 197602 250504
rect 203518 250452 203524 250504
rect 203576 250492 203582 250504
rect 215938 250492 215944 250504
rect 203576 250464 215944 250492
rect 203576 250452 203582 250464
rect 215938 250452 215944 250464
rect 215996 250452 216002 250504
rect 216048 250492 216076 250600
rect 340046 250588 340052 250640
rect 340104 250628 340110 250640
rect 356882 250628 356888 250640
rect 340104 250600 356888 250628
rect 340104 250588 340110 250600
rect 356882 250588 356888 250600
rect 356940 250588 356946 250640
rect 370406 250588 370412 250640
rect 370464 250628 370470 250640
rect 421558 250628 421564 250640
rect 370464 250600 421564 250628
rect 370464 250588 370470 250600
rect 421558 250588 421564 250600
rect 421616 250588 421622 250640
rect 219066 250520 219072 250572
rect 219124 250560 219130 250572
rect 235994 250560 236000 250572
rect 219124 250532 236000 250560
rect 219124 250520 219130 250532
rect 235994 250520 236000 250532
rect 236052 250520 236058 250572
rect 338482 250520 338488 250572
rect 338540 250560 338546 250572
rect 357618 250560 357624 250572
rect 338540 250532 357624 250560
rect 338540 250520 338546 250532
rect 357618 250520 357624 250532
rect 357676 250520 357682 250572
rect 370958 250520 370964 250572
rect 371016 250560 371022 250572
rect 425698 250560 425704 250572
rect 371016 250532 425704 250560
rect 371016 250520 371022 250532
rect 425698 250520 425704 250532
rect 425756 250520 425762 250572
rect 499022 250520 499028 250572
rect 499080 250560 499086 250572
rect 517698 250560 517704 250572
rect 499080 250532 517704 250560
rect 499080 250520 499086 250532
rect 517698 250520 517704 250532
rect 517756 250520 517762 250572
rect 219526 250492 219532 250504
rect 216048 250464 219532 250492
rect 219526 250452 219532 250464
rect 219584 250492 219590 250504
rect 267734 250492 267740 250504
rect 219584 250464 267740 250492
rect 219584 250452 219590 250464
rect 267734 250452 267740 250464
rect 267792 250452 267798 250504
rect 351730 250452 351736 250504
rect 351788 250492 351794 250504
rect 358078 250492 358084 250504
rect 351788 250464 358084 250492
rect 351788 250452 351794 250464
rect 358078 250452 358084 250464
rect 358136 250452 358142 250504
rect 370866 250452 370872 250504
rect 370924 250492 370930 250504
rect 427078 250492 427084 250504
rect 370924 250464 427084 250492
rect 370924 250452 370930 250464
rect 427078 250452 427084 250464
rect 427136 250452 427142 250504
rect 517606 250248 517612 250300
rect 517664 250288 517670 250300
rect 518066 250288 518072 250300
rect 517664 250260 518072 250288
rect 517664 250248 517670 250260
rect 518066 250248 518072 250260
rect 518124 250248 518130 250300
rect 510890 249908 510896 249960
rect 510948 249948 510954 249960
rect 517514 249948 517520 249960
rect 510948 249920 517520 249948
rect 510948 249908 510954 249920
rect 517514 249908 517520 249920
rect 517572 249908 517578 249960
rect 190914 249772 190920 249824
rect 190972 249812 190978 249824
rect 203518 249812 203524 249824
rect 190972 249784 203524 249812
rect 190972 249772 190978 249784
rect 203518 249772 203524 249784
rect 203576 249772 203582 249824
rect 218514 249772 218520 249824
rect 218572 249812 218578 249824
rect 221366 249812 221372 249824
rect 218572 249784 221372 249812
rect 218572 249772 218578 249784
rect 221366 249772 221372 249784
rect 221424 249772 221430 249824
rect 43898 249704 43904 249756
rect 43956 249744 43962 249756
rect 58710 249744 58716 249756
rect 43956 249716 58716 249744
rect 43956 249704 43962 249716
rect 58710 249704 58716 249716
rect 58768 249704 58774 249756
rect 56962 248956 56968 249008
rect 57020 248996 57026 249008
rect 62114 248996 62120 249008
rect 57020 248968 62120 248996
rect 57020 248956 57026 248968
rect 62114 248956 62120 248968
rect 62172 248956 62178 249008
rect 3050 202784 3056 202836
rect 3108 202824 3114 202836
rect 42058 202824 42064 202836
rect 3108 202796 42064 202824
rect 3108 202784 3114 202796
rect 42058 202784 42064 202796
rect 42116 202784 42122 202836
rect 520182 182180 520188 182232
rect 520240 182220 520246 182232
rect 580258 182220 580264 182232
rect 520240 182192 580264 182220
rect 520240 182180 520246 182192
rect 580258 182180 580264 182192
rect 580316 182180 580322 182232
rect 519538 182112 519544 182164
rect 519596 182152 519602 182164
rect 580350 182152 580356 182164
rect 519596 182124 580356 182152
rect 519596 182112 519602 182124
rect 580350 182112 580356 182124
rect 580408 182112 580414 182164
rect 368014 175176 368020 175228
rect 368072 175216 368078 175228
rect 376846 175216 376852 175228
rect 368072 175188 376852 175216
rect 368072 175176 368078 175188
rect 376846 175176 376852 175188
rect 376904 175176 376910 175228
rect 43990 173816 43996 173868
rect 44048 173856 44054 173868
rect 57790 173856 57796 173868
rect 44048 173828 57796 173856
rect 44048 173816 44054 173828
rect 57790 173816 57796 173828
rect 57848 173816 57854 173868
rect 203518 173816 203524 173868
rect 203576 173856 203582 173868
rect 204162 173856 204168 173868
rect 203576 173828 204168 173856
rect 203576 173816 203582 173828
rect 204162 173816 204168 173828
rect 204220 173856 204226 173868
rect 216674 173856 216680 173868
rect 204220 173828 216680 173856
rect 204220 173816 204226 173828
rect 216674 173816 216680 173828
rect 216732 173816 216738 173868
rect 366726 173816 366732 173868
rect 366784 173856 366790 173868
rect 377122 173856 377128 173868
rect 366784 173828 377128 173856
rect 366784 173816 366790 173828
rect 377122 173816 377128 173828
rect 377180 173816 377186 173868
rect 206462 173748 206468 173800
rect 206520 173788 206526 173800
rect 217042 173788 217048 173800
rect 206520 173760 217048 173788
rect 206520 173748 206526 173760
rect 217042 173748 217048 173760
rect 217100 173748 217106 173800
rect 197998 173136 198004 173188
rect 198056 173176 198062 173188
rect 204162 173176 204168 173188
rect 198056 173148 204168 173176
rect 198056 173136 198062 173148
rect 204162 173136 204168 173148
rect 204220 173136 204226 173188
rect 358078 173136 358084 173188
rect 358136 173176 358142 173188
rect 376846 173176 376852 173188
rect 358136 173148 376852 173176
rect 358136 173136 358142 173148
rect 376846 173136 376852 173148
rect 376904 173136 376910 173188
rect 54386 165520 54392 165572
rect 54444 165560 54450 165572
rect 56502 165560 56508 165572
rect 54444 165532 56508 165560
rect 54444 165520 54450 165532
rect 56502 165520 56508 165532
rect 56560 165520 56566 165572
rect 50614 164636 50620 164688
rect 50672 164676 50678 164688
rect 96062 164676 96068 164688
rect 50672 164648 96068 164676
rect 50672 164636 50678 164648
rect 96062 164636 96068 164648
rect 96120 164636 96126 164688
rect 55674 164568 55680 164620
rect 55732 164608 55738 164620
rect 56502 164608 56508 164620
rect 55732 164580 56508 164608
rect 55732 164568 55738 164580
rect 56502 164568 56508 164580
rect 56560 164608 56566 164620
rect 115750 164608 115756 164620
rect 56560 164580 115756 164608
rect 56560 164568 56566 164580
rect 115750 164568 115756 164580
rect 115808 164568 115814 164620
rect 59170 164500 59176 164552
rect 59228 164540 59234 164552
rect 140866 164540 140872 164552
rect 59228 164512 140872 164540
rect 59228 164500 59234 164512
rect 140866 164500 140872 164512
rect 140924 164500 140930 164552
rect 55950 164432 55956 164484
rect 56008 164472 56014 164484
rect 138474 164472 138480 164484
rect 56008 164444 138480 164472
rect 56008 164432 56014 164444
rect 138474 164432 138480 164444
rect 138532 164432 138538 164484
rect 42518 164364 42524 164416
rect 42576 164404 42582 164416
rect 143534 164404 143540 164416
rect 42576 164376 143540 164404
rect 42576 164364 42582 164376
rect 143534 164364 143540 164376
rect 143592 164364 143598 164416
rect 373442 164364 373448 164416
rect 373500 164404 373506 164416
rect 425974 164404 425980 164416
rect 373500 164376 425980 164404
rect 373500 164364 373506 164376
rect 425974 164364 425980 164376
rect 426032 164364 426038 164416
rect 39850 164296 39856 164348
rect 39908 164336 39914 164348
rect 163314 164336 163320 164348
rect 39908 164308 163320 164336
rect 39908 164296 39914 164308
rect 163314 164296 163320 164308
rect 163372 164296 163378 164348
rect 210694 164296 210700 164348
rect 210752 164336 210758 164348
rect 261018 164336 261024 164348
rect 210752 164308 261024 164336
rect 210752 164296 210758 164308
rect 261018 164296 261024 164308
rect 261076 164296 261082 164348
rect 369394 164296 369400 164348
rect 369452 164336 369458 164348
rect 450998 164336 451004 164348
rect 369452 164308 451004 164336
rect 369452 164296 369458 164308
rect 450998 164296 451004 164308
rect 451056 164296 451062 164348
rect 41322 164228 41328 164280
rect 41380 164268 41386 164280
rect 165890 164268 165896 164280
rect 41380 164240 165896 164268
rect 41380 164228 41386 164240
rect 165890 164228 165896 164240
rect 165948 164228 165954 164280
rect 203610 164228 203616 164280
rect 203668 164268 203674 164280
rect 288250 164268 288256 164280
rect 203668 164240 288256 164268
rect 203668 164228 203674 164240
rect 288250 164228 288256 164240
rect 288308 164228 288314 164280
rect 365254 164228 365260 164280
rect 365312 164268 365318 164280
rect 480898 164268 480904 164280
rect 365312 164240 480904 164268
rect 365312 164228 365318 164240
rect 480898 164228 480904 164240
rect 480956 164228 480962 164280
rect 357526 164160 357532 164212
rect 357584 164200 357590 164212
rect 360194 164200 360200 164212
rect 357584 164172 360200 164200
rect 357584 164160 357590 164172
rect 360194 164160 360200 164172
rect 360252 164160 360258 164212
rect 374914 164160 374920 164212
rect 374972 164200 374978 164212
rect 375742 164200 375748 164212
rect 374972 164172 375748 164200
rect 374972 164160 374978 164172
rect 375742 164160 375748 164172
rect 375800 164160 375806 164212
rect 375926 164160 375932 164212
rect 375984 164200 375990 164212
rect 393958 164200 393964 164212
rect 375984 164172 393964 164200
rect 375984 164160 375990 164172
rect 393958 164160 393964 164172
rect 394016 164160 394022 164212
rect 356698 164092 356704 164144
rect 356756 164132 356762 164144
rect 418430 164132 418436 164144
rect 356756 164104 418436 164132
rect 356756 164092 356762 164104
rect 418430 164092 418436 164104
rect 418488 164092 418494 164144
rect 52270 164024 52276 164076
rect 52328 164064 52334 164076
rect 101030 164064 101036 164076
rect 52328 164036 101036 164064
rect 52328 164024 52334 164036
rect 101030 164024 101036 164036
rect 101088 164024 101094 164076
rect 358262 164024 358268 164076
rect 358320 164064 358326 164076
rect 421006 164064 421012 164076
rect 358320 164036 421012 164064
rect 358320 164024 358326 164036
rect 421006 164024 421012 164036
rect 421064 164024 421070 164076
rect 49418 163956 49424 164008
rect 49476 163996 49482 164008
rect 98454 163996 98460 164008
rect 49476 163968 98460 163996
rect 49476 163956 49482 163968
rect 98454 163956 98460 163968
rect 98512 163956 98518 164008
rect 367830 163956 367836 164008
rect 367888 163996 367894 164008
rect 430942 163996 430948 164008
rect 367888 163968 430948 163996
rect 367888 163956 367894 163968
rect 430942 163956 430948 163968
rect 431000 163956 431006 164008
rect 50890 163888 50896 163940
rect 50948 163928 50954 163940
rect 103514 163928 103520 163940
rect 50948 163900 103520 163928
rect 50948 163888 50954 163900
rect 103514 163888 103520 163900
rect 103572 163888 103578 163940
rect 211982 163888 211988 163940
rect 212040 163928 212046 163940
rect 265894 163928 265900 163940
rect 212040 163900 265900 163928
rect 212040 163888 212046 163900
rect 265894 163888 265900 163900
rect 265952 163888 265958 163940
rect 358354 163888 358360 163940
rect 358412 163928 358418 163940
rect 423490 163928 423496 163940
rect 358412 163900 423496 163928
rect 358412 163888 358418 163900
rect 423490 163888 423496 163900
rect 423548 163888 423554 163940
rect 52178 163820 52184 163872
rect 52236 163860 52242 163872
rect 105906 163860 105912 163872
rect 52236 163832 105912 163860
rect 52236 163820 52242 163832
rect 105906 163820 105912 163832
rect 105964 163820 105970 163872
rect 110782 163820 110788 163872
rect 110840 163860 110846 163872
rect 111150 163860 111156 163872
rect 110840 163832 111156 163860
rect 110840 163820 110846 163832
rect 111150 163820 111156 163832
rect 111208 163860 111214 163872
rect 196618 163860 196624 163872
rect 111208 163832 196624 163860
rect 111208 163820 111214 163832
rect 196618 163820 196624 163832
rect 196676 163820 196682 163872
rect 204898 163820 204904 163872
rect 204956 163860 204962 163872
rect 285950 163860 285956 163872
rect 204956 163832 285956 163860
rect 204956 163820 204962 163832
rect 285950 163820 285956 163832
rect 286008 163820 286014 163872
rect 362494 163820 362500 163872
rect 362552 163860 362558 163872
rect 428182 163860 428188 163872
rect 362552 163832 428188 163860
rect 362552 163820 362558 163832
rect 428182 163820 428188 163832
rect 428240 163820 428246 163872
rect 438854 163820 438860 163872
rect 438912 163860 438918 163872
rect 516594 163860 516600 163872
rect 438912 163832 516600 163860
rect 438912 163820 438918 163832
rect 516594 163820 516600 163832
rect 516652 163820 516658 163872
rect 47946 163752 47952 163804
rect 48004 163792 48010 163804
rect 52270 163792 52276 163804
rect 48004 163764 52276 163792
rect 48004 163752 48010 163764
rect 52270 163752 52276 163764
rect 52328 163752 52334 163804
rect 59906 163752 59912 163804
rect 59964 163792 59970 163804
rect 145926 163792 145932 163804
rect 59964 163764 145932 163792
rect 59964 163752 59970 163764
rect 145926 163752 145932 163764
rect 145984 163752 145990 163804
rect 213178 163752 213184 163804
rect 213236 163792 213242 163804
rect 303430 163792 303436 163804
rect 213236 163764 303436 163792
rect 213236 163752 213242 163764
rect 303430 163752 303436 163764
rect 303488 163752 303494 163804
rect 373534 163752 373540 163804
rect 373592 163792 373598 163804
rect 475838 163792 475844 163804
rect 373592 163764 475844 163792
rect 373592 163752 373598 163764
rect 475838 163752 475844 163764
rect 475896 163752 475902 163804
rect 50798 163684 50804 163736
rect 50856 163724 50862 163736
rect 108206 163724 108212 163736
rect 50856 163696 108212 163724
rect 50856 163684 50862 163696
rect 108206 163684 108212 163696
rect 108264 163684 108270 163736
rect 110506 163684 110512 163736
rect 110564 163724 110570 163736
rect 196802 163724 196808 163736
rect 110564 163696 196808 163724
rect 110564 163684 110570 163696
rect 196802 163684 196808 163696
rect 196860 163684 196866 163736
rect 206370 163684 206376 163736
rect 206428 163724 206434 163736
rect 298462 163724 298468 163736
rect 206428 163696 298468 163724
rect 206428 163684 206434 163696
rect 298462 163684 298468 163696
rect 298520 163684 298526 163736
rect 370774 163684 370780 163736
rect 370832 163724 370838 163736
rect 473446 163724 473452 163736
rect 370832 163696 473452 163724
rect 370832 163684 370838 163696
rect 473446 163684 473452 163696
rect 473504 163684 473510 163736
rect 59078 163616 59084 163668
rect 59136 163656 59142 163668
rect 148502 163656 148508 163668
rect 59136 163628 148508 163656
rect 59136 163616 59142 163628
rect 148502 163616 148508 163628
rect 148560 163616 148566 163668
rect 207750 163616 207756 163668
rect 207808 163656 207814 163668
rect 300854 163656 300860 163668
rect 207808 163628 300860 163656
rect 207808 163616 207814 163628
rect 300854 163616 300860 163628
rect 300912 163616 300918 163668
rect 367922 163616 367928 163668
rect 367980 163656 367986 163668
rect 470962 163656 470968 163668
rect 367980 163628 470968 163656
rect 367980 163616 367986 163628
rect 470962 163616 470968 163628
rect 471020 163616 471026 163668
rect 510522 163616 510528 163668
rect 510580 163656 510586 163668
rect 517514 163656 517520 163668
rect 510580 163628 517520 163656
rect 510580 163616 510586 163628
rect 517514 163616 517520 163628
rect 517572 163616 517578 163668
rect 58894 163548 58900 163600
rect 58952 163588 58958 163600
rect 150894 163588 150900 163600
rect 58952 163560 150900 163588
rect 58952 163548 58958 163560
rect 150894 163548 150900 163560
rect 150952 163548 150958 163600
rect 209130 163548 209136 163600
rect 209188 163588 209194 163600
rect 305914 163588 305920 163600
rect 209188 163560 305920 163588
rect 209188 163548 209194 163560
rect 305914 163548 305920 163560
rect 305972 163548 305978 163600
rect 372062 163548 372068 163600
rect 372120 163588 372126 163600
rect 478414 163588 478420 163600
rect 372120 163560 478420 163588
rect 372120 163548 372126 163560
rect 478414 163548 478420 163560
rect 478472 163548 478478 163600
rect 59998 163480 60004 163532
rect 60056 163520 60062 163532
rect 153378 163520 153384 163532
rect 60056 163492 153384 163520
rect 60056 163480 60062 163492
rect 153378 163480 153384 163492
rect 153436 163480 153442 163532
rect 214742 163480 214748 163532
rect 214800 163520 214806 163532
rect 313366 163520 313372 163532
rect 214800 163492 313372 163520
rect 214800 163480 214806 163492
rect 313366 163480 313372 163492
rect 313424 163480 313430 163532
rect 366634 163480 366640 163532
rect 366692 163520 366698 163532
rect 483382 163520 483388 163532
rect 366692 163492 483388 163520
rect 366692 163480 366698 163492
rect 483382 163480 483388 163492
rect 483440 163480 483446 163532
rect 218606 163412 218612 163464
rect 218664 163452 218670 163464
rect 219710 163452 219716 163464
rect 218664 163424 219716 163452
rect 218664 163412 218670 163424
rect 219710 163412 219716 163424
rect 219768 163452 219774 163464
rect 220446 163452 220452 163464
rect 219768 163424 220452 163452
rect 219768 163412 219774 163424
rect 220446 163412 220452 163424
rect 220504 163412 220510 163464
rect 373166 163140 373172 163192
rect 373224 163180 373230 163192
rect 374178 163180 374184 163192
rect 373224 163152 374184 163180
rect 373224 163140 373230 163152
rect 374178 163140 374184 163152
rect 374236 163180 374242 163192
rect 375282 163180 375288 163192
rect 374236 163152 375288 163180
rect 374236 163140 374242 163152
rect 375282 163140 375288 163152
rect 375340 163140 375346 163192
rect 53190 163004 53196 163056
rect 53248 163044 53254 163056
rect 113450 163044 113456 163056
rect 53248 163016 113456 163044
rect 53248 163004 53254 163016
rect 113450 163004 113456 163016
rect 113508 163044 113514 163056
rect 123018 163044 123024 163056
rect 113508 163016 123024 163044
rect 113508 163004 113514 163016
rect 123018 163004 123024 163016
rect 123076 163004 123082 163056
rect 373718 163004 373724 163056
rect 373776 163044 373782 163056
rect 374914 163044 374920 163056
rect 373776 163016 374920 163044
rect 373776 163004 373782 163016
rect 374914 163004 374920 163016
rect 374972 163044 374978 163056
rect 429746 163044 429752 163056
rect 374972 163016 429752 163044
rect 374972 163004 374978 163016
rect 429746 163004 429752 163016
rect 429804 163004 429810 163056
rect 52270 162936 52276 162988
rect 52328 162976 52334 162988
rect 114370 162976 114376 162988
rect 52328 162948 114376 162976
rect 52328 162936 52334 162948
rect 114370 162936 114376 162948
rect 114428 162936 114434 162988
rect 217134 162936 217140 162988
rect 217192 162976 217198 162988
rect 236638 162976 236644 162988
rect 217192 162948 236644 162976
rect 217192 162936 217198 162948
rect 236638 162936 236644 162948
rect 236696 162936 236702 162988
rect 375282 162936 375288 162988
rect 375340 162976 375346 162988
rect 431954 162976 431960 162988
rect 375340 162948 431960 162976
rect 375340 162936 375346 162948
rect 431954 162936 431960 162948
rect 432012 162936 432018 162988
rect 55766 162868 55772 162920
rect 55824 162908 55830 162920
rect 118050 162908 118056 162920
rect 55824 162880 118056 162908
rect 55824 162868 55830 162880
rect 118050 162868 118056 162880
rect 118108 162868 118114 162920
rect 197446 162868 197452 162920
rect 197504 162908 197510 162920
rect 200114 162908 200120 162920
rect 197504 162880 200120 162908
rect 197504 162868 197510 162880
rect 200114 162868 200120 162880
rect 200172 162868 200178 162920
rect 220446 162868 220452 162920
rect 220504 162908 220510 162920
rect 267550 162908 267556 162920
rect 220504 162880 267556 162908
rect 220504 162868 220510 162880
rect 267550 162868 267556 162880
rect 267608 162868 267614 162920
rect 375742 162868 375748 162920
rect 375800 162908 375806 162920
rect 436922 162908 436928 162920
rect 375800 162880 436928 162908
rect 375800 162868 375806 162880
rect 436922 162868 436928 162880
rect 436980 162868 436986 162920
rect 50522 162800 50528 162852
rect 50580 162840 50586 162852
rect 155954 162840 155960 162852
rect 50580 162812 155960 162840
rect 50580 162800 50586 162812
rect 155954 162800 155960 162812
rect 156012 162800 156018 162852
rect 210602 162800 210608 162852
rect 210660 162840 210666 162852
rect 320910 162840 320916 162852
rect 210660 162812 320916 162840
rect 210660 162800 210666 162812
rect 320910 162800 320916 162812
rect 320968 162800 320974 162852
rect 356698 162800 356704 162852
rect 356756 162840 356762 162852
rect 357066 162840 357072 162852
rect 356756 162812 357072 162840
rect 356756 162800 356762 162812
rect 357066 162800 357072 162812
rect 357124 162800 357130 162852
rect 365162 162800 365168 162852
rect 365220 162840 365226 162852
rect 458358 162840 458364 162852
rect 365220 162812 458364 162840
rect 365220 162800 365226 162812
rect 458358 162800 458364 162812
rect 458416 162800 458422 162852
rect 517606 162800 517612 162852
rect 517664 162840 517670 162852
rect 517882 162840 517888 162852
rect 517664 162812 517888 162840
rect 517664 162800 517670 162812
rect 517882 162800 517888 162812
rect 517940 162800 517946 162852
rect 56134 162732 56140 162784
rect 56192 162772 56198 162784
rect 135990 162772 135996 162784
rect 56192 162744 135996 162772
rect 56192 162732 56198 162744
rect 135990 162732 135996 162744
rect 136048 162732 136054 162784
rect 214558 162732 214564 162784
rect 214616 162772 214622 162784
rect 293218 162772 293224 162784
rect 214616 162744 293224 162772
rect 214616 162732 214622 162744
rect 293218 162732 293224 162744
rect 293276 162732 293282 162784
rect 369210 162732 369216 162784
rect 369268 162772 369274 162784
rect 455782 162772 455788 162784
rect 369268 162744 455788 162772
rect 369268 162732 369274 162744
rect 455782 162732 455788 162744
rect 455840 162732 455846 162784
rect 517514 162732 517520 162784
rect 517572 162772 517578 162784
rect 517974 162772 517980 162784
rect 517572 162744 517980 162772
rect 517572 162732 517578 162744
rect 517974 162732 517980 162744
rect 518032 162732 518038 162784
rect 55122 162664 55128 162716
rect 55180 162704 55186 162716
rect 133414 162704 133420 162716
rect 55180 162676 133420 162704
rect 55180 162664 55186 162676
rect 133414 162664 133420 162676
rect 133472 162664 133478 162716
rect 211798 162664 211804 162716
rect 211856 162704 211862 162716
rect 280798 162704 280804 162716
rect 211856 162676 280804 162704
rect 211856 162664 211862 162676
rect 280798 162664 280804 162676
rect 280856 162664 280862 162716
rect 370682 162664 370688 162716
rect 370740 162704 370746 162716
rect 453390 162704 453396 162716
rect 370740 162676 453396 162704
rect 370740 162664 370746 162676
rect 453390 162664 453396 162676
rect 453448 162664 453454 162716
rect 56318 162596 56324 162648
rect 56376 162636 56382 162648
rect 130838 162636 130844 162648
rect 56376 162608 130844 162636
rect 56376 162596 56382 162608
rect 130838 162596 130844 162608
rect 130896 162596 130902 162648
rect 218790 162596 218796 162648
rect 218848 162636 218854 162648
rect 283742 162636 283748 162648
rect 218848 162608 283748 162636
rect 218848 162596 218854 162608
rect 283742 162596 283748 162608
rect 283800 162596 283806 162648
rect 366542 162596 366548 162648
rect 366600 162636 366606 162648
rect 448238 162636 448244 162648
rect 366600 162608 448244 162636
rect 366600 162596 366606 162608
rect 448238 162596 448244 162608
rect 448296 162596 448302 162648
rect 55030 162528 55036 162580
rect 55088 162568 55094 162580
rect 128354 162568 128360 162580
rect 55088 162540 128360 162568
rect 55088 162528 55094 162540
rect 128354 162528 128360 162540
rect 128412 162528 128418 162580
rect 204990 162528 204996 162580
rect 205048 162568 205054 162580
rect 263686 162568 263692 162580
rect 205048 162540 263692 162568
rect 205048 162528 205054 162540
rect 263686 162528 263692 162540
rect 263744 162528 263750 162580
rect 360930 162528 360936 162580
rect 360988 162568 360994 162580
rect 435910 162568 435916 162580
rect 360988 162540 435916 162568
rect 360988 162528 360994 162540
rect 435910 162528 435916 162540
rect 435968 162528 435974 162580
rect 54938 162460 54944 162512
rect 54996 162500 55002 162512
rect 122742 162500 122748 162512
rect 54996 162472 122748 162500
rect 54996 162460 55002 162472
rect 122742 162460 122748 162472
rect 122800 162460 122806 162512
rect 123018 162460 123024 162512
rect 123076 162500 123082 162512
rect 196710 162500 196716 162512
rect 123076 162472 196716 162500
rect 123076 162460 123082 162472
rect 196710 162460 196716 162472
rect 196768 162460 196774 162512
rect 214650 162460 214656 162512
rect 214708 162500 214714 162512
rect 273438 162500 273444 162512
rect 214708 162472 273444 162500
rect 214708 162460 214714 162472
rect 273438 162460 273444 162472
rect 273496 162460 273502 162512
rect 371970 162460 371976 162512
rect 372028 162500 372034 162512
rect 445846 162500 445852 162512
rect 372028 162472 445852 162500
rect 372028 162460 372034 162472
rect 445846 162460 445852 162472
rect 445904 162460 445910 162512
rect 56226 162392 56232 162444
rect 56284 162432 56290 162444
rect 125870 162432 125876 162444
rect 56284 162404 125876 162432
rect 56284 162392 56290 162404
rect 125870 162392 125876 162404
rect 125928 162392 125934 162444
rect 210418 162392 210424 162444
rect 210476 162432 210482 162444
rect 268286 162432 268292 162444
rect 210476 162404 268292 162432
rect 210476 162392 210482 162404
rect 268286 162392 268292 162404
rect 268344 162392 268350 162444
rect 363782 162392 363788 162444
rect 363840 162432 363846 162444
rect 438486 162432 438492 162444
rect 363840 162404 438492 162432
rect 363840 162392 363846 162404
rect 438486 162392 438492 162404
rect 438544 162392 438550 162444
rect 53374 162324 53380 162376
rect 53432 162364 53438 162376
rect 120718 162364 120724 162376
rect 53432 162336 120724 162364
rect 53432 162324 53438 162336
rect 120718 162324 120724 162336
rect 120776 162324 120782 162376
rect 183462 162324 183468 162376
rect 183520 162364 183526 162376
rect 197354 162364 197360 162376
rect 183520 162336 197360 162364
rect 183520 162324 183526 162336
rect 197354 162324 197360 162336
rect 197412 162324 197418 162376
rect 218882 162324 218888 162376
rect 218940 162364 218946 162376
rect 276106 162364 276112 162376
rect 218940 162336 276112 162364
rect 218940 162324 218946 162336
rect 276106 162324 276112 162336
rect 276164 162324 276170 162376
rect 373350 162324 373356 162376
rect 373408 162364 373414 162376
rect 443454 162364 443460 162376
rect 373408 162336 443460 162364
rect 373408 162324 373414 162336
rect 443454 162324 443460 162336
rect 443512 162324 443518 162376
rect 53282 162256 53288 162308
rect 53340 162296 53346 162308
rect 116026 162296 116032 162308
rect 53340 162268 116032 162296
rect 53340 162256 53346 162268
rect 116026 162256 116032 162268
rect 116084 162256 116090 162308
rect 202138 162256 202144 162308
rect 202196 162296 202202 162308
rect 256142 162296 256148 162308
rect 202196 162268 256148 162296
rect 202196 162256 202202 162268
rect 256142 162256 256148 162268
rect 256200 162256 256206 162308
rect 343450 162256 343456 162308
rect 343508 162296 343514 162308
rect 356698 162296 356704 162308
rect 343508 162268 356704 162296
rect 343508 162256 343514 162268
rect 356698 162256 356704 162268
rect 356756 162256 356762 162308
rect 374822 162256 374828 162308
rect 374880 162296 374886 162308
rect 440878 162296 440884 162308
rect 374880 162268 440884 162296
rect 374880 162256 374886 162268
rect 440878 162256 440884 162268
rect 440936 162256 440942 162308
rect 503254 162256 503260 162308
rect 503312 162296 503318 162308
rect 517514 162296 517520 162308
rect 503312 162268 517520 162296
rect 503312 162256 503318 162268
rect 517514 162256 517520 162268
rect 517572 162256 517578 162308
rect 56042 162188 56048 162240
rect 56100 162228 56106 162240
rect 118326 162228 118332 162240
rect 56100 162200 118332 162228
rect 56100 162188 56106 162200
rect 118326 162188 118332 162200
rect 118384 162188 118390 162240
rect 183186 162188 183192 162240
rect 183244 162228 183250 162240
rect 197446 162228 197452 162240
rect 183244 162200 197452 162228
rect 183244 162188 183250 162200
rect 197446 162188 197452 162200
rect 197504 162188 197510 162240
rect 211890 162188 211896 162240
rect 211948 162228 211954 162240
rect 258350 162228 258356 162240
rect 211948 162200 258356 162228
rect 211948 162188 211954 162200
rect 258350 162188 258356 162200
rect 258408 162188 258414 162240
rect 369118 162188 369124 162240
rect 369176 162228 369182 162240
rect 433518 162228 433524 162240
rect 369176 162200 433524 162228
rect 369176 162188 369182 162200
rect 433518 162188 433524 162200
rect 433576 162188 433582 162240
rect 100018 162120 100024 162172
rect 100076 162160 100082 162172
rect 100754 162160 100760 162172
rect 100076 162132 100760 162160
rect 100076 162120 100082 162132
rect 100754 162120 100760 162132
rect 100812 162120 100818 162172
rect 112806 162120 112812 162172
rect 112864 162160 112870 162172
rect 113082 162160 113088 162172
rect 112864 162132 113088 162160
rect 112864 162120 112870 162132
rect 113082 162120 113088 162132
rect 113140 162160 113146 162172
rect 197814 162160 197820 162172
rect 113140 162132 197820 162160
rect 113140 162120 113146 162132
rect 197814 162120 197820 162132
rect 197872 162120 197878 162172
rect 209038 162120 209044 162172
rect 209096 162160 209102 162172
rect 253566 162160 253572 162172
rect 209096 162132 253572 162160
rect 209096 162120 209102 162132
rect 253566 162120 253572 162132
rect 253624 162120 253630 162172
rect 343358 162120 343364 162172
rect 343416 162160 343422 162172
rect 357526 162160 357532 162172
rect 343416 162132 357532 162160
rect 343416 162120 343422 162132
rect 357526 162120 357532 162132
rect 357584 162120 357590 162172
rect 362402 162120 362408 162172
rect 362460 162160 362466 162172
rect 410610 162160 410616 162172
rect 362460 162132 410616 162160
rect 362460 162120 362466 162132
rect 410610 162120 410616 162132
rect 410668 162120 410674 162172
rect 415302 162120 415308 162172
rect 415360 162160 415366 162172
rect 418246 162160 418252 162172
rect 415360 162132 418252 162160
rect 415360 162120 415366 162132
rect 418246 162120 418252 162132
rect 418304 162120 418310 162172
rect 503622 162120 503628 162172
rect 503680 162160 503686 162172
rect 517606 162160 517612 162172
rect 503680 162132 517612 162160
rect 503680 162120 503686 162132
rect 517606 162120 517612 162132
rect 517664 162120 517670 162172
rect 53466 162052 53472 162104
rect 53524 162092 53530 162104
rect 110966 162092 110972 162104
rect 53524 162064 110972 162092
rect 53524 162052 53530 162064
rect 110966 162052 110972 162064
rect 111024 162052 111030 162104
rect 210510 162052 210516 162104
rect 210568 162092 210574 162104
rect 250622 162092 250628 162104
rect 210568 162064 250628 162092
rect 210568 162052 210574 162064
rect 250622 162052 250628 162064
rect 250680 162052 250686 162104
rect 367738 162052 367744 162104
rect 367796 162092 367802 162104
rect 408310 162092 408316 162104
rect 367796 162064 408316 162092
rect 367796 162052 367802 162064
rect 408310 162052 408316 162064
rect 408368 162052 408374 162104
rect 49326 161984 49332 162036
rect 49384 162024 49390 162036
rect 90726 162024 90732 162036
rect 49384 161996 90732 162024
rect 49384 161984 49390 161996
rect 90726 161984 90732 161996
rect 90784 161984 90790 162036
rect 216030 161984 216036 162036
rect 216088 162024 216094 162036
rect 248230 162024 248236 162036
rect 216088 161996 248236 162024
rect 216088 161984 216094 161996
rect 248230 161984 248236 161996
rect 248288 161984 248294 162036
rect 374730 161984 374736 162036
rect 374788 162024 374794 162036
rect 413554 162024 413560 162036
rect 374788 161996 413560 162024
rect 374788 161984 374794 161996
rect 413554 161984 413560 161996
rect 413612 161984 413618 162036
rect 56410 161916 56416 161968
rect 56468 161956 56474 161968
rect 88334 161956 88340 161968
rect 56468 161928 88340 161956
rect 56468 161916 56474 161928
rect 88334 161916 88340 161928
rect 88392 161916 88398 161968
rect 378778 161916 378784 161968
rect 378836 161956 378842 161968
rect 416038 161956 416044 161968
rect 378836 161928 416044 161956
rect 378836 161916 378842 161928
rect 416038 161916 416044 161928
rect 416096 161916 416102 161968
rect 54846 161848 54852 161900
rect 54904 161888 54910 161900
rect 113174 161888 113180 161900
rect 54904 161860 113180 161888
rect 54904 161848 54910 161860
rect 113174 161848 113180 161860
rect 113232 161848 113238 161900
rect 428734 161508 428740 161560
rect 428792 161548 428798 161560
rect 435726 161548 435732 161560
rect 428792 161520 435732 161548
rect 428792 161508 428798 161520
rect 435726 161508 435732 161520
rect 435784 161508 435790 161560
rect 98638 161440 98644 161492
rect 98696 161480 98702 161492
rect 103790 161480 103796 161492
rect 98696 161452 103796 161480
rect 98696 161440 98702 161452
rect 103790 161440 103796 161452
rect 103848 161440 103854 161492
rect 56870 161372 56876 161424
rect 56928 161412 56934 161424
rect 115934 161412 115940 161424
rect 56928 161384 115940 161412
rect 56928 161372 56934 161384
rect 115934 161372 115940 161384
rect 115992 161372 115998 161424
rect 219526 161372 219532 161424
rect 219584 161412 219590 161424
rect 267734 161412 267740 161424
rect 219584 161384 267740 161412
rect 219584 161372 219590 161384
rect 267734 161372 267740 161384
rect 267792 161372 267798 161424
rect 379974 161372 379980 161424
rect 380032 161412 380038 161424
rect 426434 161412 426440 161424
rect 380032 161384 426440 161412
rect 380032 161372 380038 161384
rect 426434 161372 426440 161384
rect 426492 161372 426498 161424
rect 58618 161304 58624 161356
rect 58676 161344 58682 161356
rect 106366 161344 106372 161356
rect 58676 161316 106372 161344
rect 58676 161304 58682 161316
rect 106366 161304 106372 161316
rect 106424 161304 106430 161356
rect 218514 161304 218520 161356
rect 218572 161344 218578 161356
rect 266354 161344 266360 161356
rect 218572 161316 266360 161344
rect 218572 161304 218578 161316
rect 266354 161304 266360 161316
rect 266412 161304 266418 161356
rect 379698 161304 379704 161356
rect 379756 161344 379762 161356
rect 425054 161344 425060 161356
rect 379756 161316 425060 161344
rect 379756 161304 379762 161316
rect 425054 161304 425060 161316
rect 425112 161304 425118 161356
rect 54202 161236 54208 161288
rect 54260 161276 54266 161288
rect 55030 161276 55036 161288
rect 54260 161248 55036 161276
rect 54260 161236 54266 161248
rect 55030 161236 55036 161248
rect 55088 161276 55094 161288
rect 99374 161276 99380 161288
rect 55088 161248 99380 161276
rect 55088 161236 55094 161248
rect 99374 161236 99380 161248
rect 99432 161236 99438 161288
rect 214282 161236 214288 161288
rect 214340 161276 214346 161288
rect 260834 161276 260840 161288
rect 214340 161248 260840 161276
rect 214340 161236 214346 161248
rect 260834 161236 260840 161248
rect 260892 161236 260898 161288
rect 219618 161168 219624 161220
rect 219676 161208 219682 161220
rect 264974 161208 264980 161220
rect 219676 161180 264980 161208
rect 219676 161168 219682 161180
rect 264974 161168 264980 161180
rect 265032 161168 265038 161220
rect 218974 161100 218980 161152
rect 219032 161140 219038 161152
rect 219342 161140 219348 161152
rect 219032 161112 219348 161140
rect 219032 161100 219038 161112
rect 219342 161100 219348 161112
rect 219400 161140 219406 161152
rect 263594 161140 263600 161152
rect 219400 161112 263600 161140
rect 219400 161100 219406 161112
rect 263594 161100 263600 161112
rect 263652 161100 263658 161152
rect 217870 161032 217876 161084
rect 217928 161072 217934 161084
rect 258074 161072 258080 161084
rect 217928 161044 258080 161072
rect 217928 161032 217934 161044
rect 258074 161032 258080 161044
rect 258132 161032 258138 161084
rect 52914 160964 52920 161016
rect 52972 161004 52978 161016
rect 57790 161004 57796 161016
rect 52972 160976 57796 161004
rect 52972 160964 52978 160976
rect 57790 160964 57796 160976
rect 57848 161004 57854 161016
rect 95234 161004 95240 161016
rect 57848 160976 95240 161004
rect 57848 160964 57854 160976
rect 95234 160964 95240 160976
rect 95292 160964 95298 161016
rect 54294 160896 54300 160948
rect 54352 160936 54358 160948
rect 59078 160936 59084 160948
rect 54352 160908 59084 160936
rect 54352 160896 54358 160908
rect 59078 160896 59084 160908
rect 59136 160936 59142 160948
rect 96614 160936 96620 160948
rect 59136 160908 96620 160936
rect 59136 160896 59142 160908
rect 96614 160896 96620 160908
rect 96672 160896 96678 160948
rect 51442 160828 51448 160880
rect 51500 160868 51506 160880
rect 55122 160868 55128 160880
rect 51500 160840 55128 160868
rect 51500 160828 51506 160840
rect 55122 160828 55128 160840
rect 55180 160868 55186 160880
rect 97994 160868 98000 160880
rect 55180 160840 98000 160868
rect 55180 160828 55186 160840
rect 97994 160828 98000 160840
rect 98052 160828 98058 160880
rect 373810 160828 373816 160880
rect 373868 160868 373874 160880
rect 374730 160868 374736 160880
rect 373868 160840 374736 160868
rect 373868 160828 373874 160840
rect 374730 160828 374736 160840
rect 374788 160868 374794 160880
rect 430574 160868 430580 160880
rect 374788 160840 430580 160868
rect 374788 160828 374794 160840
rect 430574 160828 430580 160840
rect 430632 160828 430638 160880
rect 59998 160760 60004 160812
rect 60056 160800 60062 160812
rect 106274 160800 106280 160812
rect 60056 160772 106280 160800
rect 60056 160760 60062 160772
rect 106274 160760 106280 160772
rect 106332 160760 106338 160812
rect 371694 160760 371700 160812
rect 371752 160800 371758 160812
rect 373626 160800 373632 160812
rect 371752 160772 373632 160800
rect 371752 160760 371758 160772
rect 373626 160760 373632 160772
rect 373684 160800 373690 160812
rect 433334 160800 433340 160812
rect 373684 160772 433340 160800
rect 373684 160760 373690 160772
rect 433334 160760 433340 160772
rect 433392 160760 433398 160812
rect 47854 160692 47860 160744
rect 47912 160732 47918 160744
rect 59354 160732 59360 160744
rect 47912 160704 59360 160732
rect 47912 160692 47918 160704
rect 59354 160692 59360 160704
rect 59412 160732 59418 160744
rect 118694 160732 118700 160744
rect 59412 160704 118700 160732
rect 59412 160692 59418 160704
rect 118694 160692 118700 160704
rect 118752 160692 118758 160744
rect 213270 160692 213276 160744
rect 213328 160732 213334 160744
rect 273254 160732 273260 160744
rect 213328 160704 273260 160732
rect 213328 160692 213334 160704
rect 273254 160692 273260 160704
rect 273312 160692 273318 160744
rect 370406 160692 370412 160744
rect 370464 160732 370470 160744
rect 374546 160732 374552 160744
rect 370464 160704 374552 160732
rect 370464 160692 370470 160704
rect 374546 160692 374552 160704
rect 374604 160732 374610 160744
rect 437382 160732 437388 160744
rect 374604 160704 437388 160732
rect 374604 160692 374610 160704
rect 437382 160692 437388 160704
rect 437440 160692 437446 160744
rect 58710 160556 58716 160608
rect 58768 160596 58774 160608
rect 59998 160596 60004 160608
rect 58768 160568 60004 160596
rect 58768 160556 58774 160568
rect 59998 160556 60004 160568
rect 60056 160556 60062 160608
rect 212166 160420 212172 160472
rect 212224 160460 212230 160472
rect 213270 160460 213276 160472
rect 212224 160432 213276 160460
rect 212224 160420 212230 160432
rect 213270 160420 213276 160432
rect 213328 160420 213334 160472
rect 58618 160080 58624 160132
rect 58676 160120 58682 160132
rect 59170 160120 59176 160132
rect 58676 160092 59176 160120
rect 58676 160080 58682 160092
rect 59170 160080 59176 160092
rect 59228 160080 59234 160132
rect 214282 160080 214288 160132
rect 214340 160120 214346 160132
rect 214742 160120 214748 160132
rect 214340 160092 214748 160120
rect 214340 160080 214346 160092
rect 214742 160080 214748 160092
rect 214800 160080 214806 160132
rect 218238 160080 218244 160132
rect 218296 160120 218302 160132
rect 218514 160120 218520 160132
rect 218296 160092 218520 160120
rect 218296 160080 218302 160092
rect 218514 160080 218520 160092
rect 218572 160080 218578 160132
rect 379790 160080 379796 160132
rect 379848 160120 379854 160132
rect 379974 160120 379980 160132
rect 379848 160092 379980 160120
rect 379848 160080 379854 160092
rect 379974 160080 379980 160092
rect 380032 160080 380038 160132
rect 214834 160012 214840 160064
rect 214892 160052 214898 160064
rect 259546 160052 259552 160064
rect 214892 160024 259552 160052
rect 214892 160012 214898 160024
rect 259546 160012 259552 160024
rect 259604 160012 259610 160064
rect 376294 160012 376300 160064
rect 376352 160052 376358 160064
rect 420914 160052 420920 160064
rect 376352 160024 420920 160052
rect 376352 160012 376358 160024
rect 420914 160012 420920 160024
rect 420972 160012 420978 160064
rect 216398 159944 216404 159996
rect 216456 159984 216462 159996
rect 259454 159984 259460 159996
rect 216456 159956 259460 159984
rect 216456 159944 216462 159956
rect 259454 159944 259460 159956
rect 259512 159944 259518 159996
rect 377674 159944 377680 159996
rect 377732 159984 377738 159996
rect 419534 159984 419540 159996
rect 377732 159956 419540 159984
rect 377732 159944 377738 159956
rect 419534 159944 419540 159956
rect 419592 159944 419598 159996
rect 215754 159536 215760 159588
rect 215812 159576 215818 159588
rect 216398 159576 216404 159588
rect 215812 159548 216404 159576
rect 215812 159536 215818 159548
rect 216398 159536 216404 159548
rect 216456 159536 216462 159588
rect 376386 159400 376392 159452
rect 376444 159440 376450 159452
rect 379606 159440 379612 159452
rect 376444 159412 379612 159440
rect 376444 159400 376450 159412
rect 379606 159400 379612 159412
rect 379664 159440 379670 159452
rect 418154 159440 418160 159452
rect 379664 159412 418160 159440
rect 379664 159400 379670 159412
rect 418154 159400 418160 159412
rect 418212 159400 418218 159452
rect 370866 159332 370872 159384
rect 370924 159372 370930 159384
rect 372246 159372 372252 159384
rect 370924 159344 372252 159372
rect 370924 159332 370930 159344
rect 372246 159332 372252 159344
rect 372304 159372 372310 159384
rect 428734 159372 428740 159384
rect 372304 159344 428740 159372
rect 372304 159332 372310 159344
rect 428734 159332 428740 159344
rect 428792 159332 428798 159384
rect 376662 158720 376668 158772
rect 376720 158760 376726 158772
rect 377674 158760 377680 158772
rect 376720 158732 377680 158760
rect 376720 158720 376726 158732
rect 377674 158720 377680 158732
rect 377732 158720 377738 158772
rect 217134 156612 217140 156664
rect 217192 156652 217198 156664
rect 217870 156652 217876 156664
rect 217192 156624 217876 156652
rect 217192 156612 217198 156624
rect 217870 156612 217876 156624
rect 217928 156612 217934 156664
rect 215018 148996 215024 149048
rect 215076 149036 215082 149048
rect 274726 149036 274732 149048
rect 215076 149008 274732 149036
rect 215076 148996 215082 149008
rect 274726 148996 274732 149008
rect 274784 148996 274790 149048
rect 380802 148996 380808 149048
rect 380860 149036 380866 149048
rect 429194 149036 429200 149048
rect 380860 149008 429200 149036
rect 380860 148996 380866 149008
rect 429194 148996 429200 149008
rect 429252 148996 429258 149048
rect 213362 148928 213368 148980
rect 213420 148968 213426 148980
rect 240134 148968 240140 148980
rect 213420 148940 240140 148968
rect 213420 148928 213426 148940
rect 240134 148928 240140 148940
rect 240192 148928 240198 148980
rect 379882 148928 379888 148980
rect 379940 148968 379946 148980
rect 412726 148968 412732 148980
rect 379940 148940 412732 148968
rect 379940 148928 379946 148940
rect 412726 148928 412732 148940
rect 412784 148928 412790 148980
rect 214926 148860 214932 148912
rect 214984 148900 214990 148912
rect 241514 148900 241520 148912
rect 214984 148872 241520 148900
rect 214984 148860 214990 148872
rect 241514 148860 241520 148872
rect 241572 148860 241578 148912
rect 373718 148860 373724 148912
rect 373776 148900 373782 148912
rect 375006 148900 375012 148912
rect 373776 148872 375012 148900
rect 373776 148860 373782 148872
rect 375006 148860 375012 148872
rect 375064 148900 375070 148912
rect 400214 148900 400220 148912
rect 375064 148872 400220 148900
rect 375064 148860 375070 148872
rect 400214 148860 400220 148872
rect 400272 148860 400278 148912
rect 215662 148792 215668 148844
rect 215720 148832 215726 148844
rect 238754 148832 238760 148844
rect 215720 148804 238760 148832
rect 215720 148792 215726 148804
rect 238754 148792 238760 148804
rect 238812 148792 238818 148844
rect 48038 148656 48044 148708
rect 48096 148696 48102 148708
rect 52086 148696 52092 148708
rect 48096 148668 52092 148696
rect 48096 148656 48102 148668
rect 52086 148656 52092 148668
rect 52144 148696 52150 148708
rect 78674 148696 78680 148708
rect 52144 148668 78680 148696
rect 52144 148656 52150 148668
rect 78674 148656 78680 148668
rect 78732 148656 78738 148708
rect 46474 148588 46480 148640
rect 46532 148628 46538 148640
rect 53374 148628 53380 148640
rect 46532 148600 53380 148628
rect 46532 148588 46538 148600
rect 53374 148588 53380 148600
rect 53432 148628 53438 148640
rect 80054 148628 80060 148640
rect 53432 148600 80060 148628
rect 53432 148588 53438 148600
rect 80054 148588 80060 148600
rect 80112 148588 80118 148640
rect 49142 148520 49148 148572
rect 49200 148560 49206 148572
rect 53282 148560 53288 148572
rect 49200 148532 53288 148560
rect 49200 148520 49206 148532
rect 53282 148520 53288 148532
rect 53340 148560 53346 148572
rect 81434 148560 81440 148572
rect 53340 148532 81440 148560
rect 53340 148520 53346 148532
rect 81434 148520 81440 148532
rect 81492 148520 81498 148572
rect 372338 148520 372344 148572
rect 372396 148560 372402 148572
rect 375006 148560 375012 148572
rect 372396 148532 375012 148560
rect 372396 148520 372402 148532
rect 375006 148520 375012 148532
rect 375064 148560 375070 148572
rect 401594 148560 401600 148572
rect 375064 148532 401600 148560
rect 375064 148520 375070 148532
rect 401594 148520 401600 148532
rect 401652 148520 401658 148572
rect 54754 148452 54760 148504
rect 54812 148492 54818 148504
rect 110782 148492 110788 148504
rect 54812 148464 110788 148492
rect 54812 148452 54818 148464
rect 110782 148452 110788 148464
rect 110840 148452 110846 148504
rect 370222 148452 370228 148504
rect 370280 148492 370286 148504
rect 371970 148492 371976 148504
rect 370280 148464 371976 148492
rect 370280 148452 370286 148464
rect 371970 148452 371976 148464
rect 372028 148492 372034 148504
rect 398834 148492 398840 148504
rect 372028 148464 398840 148492
rect 372028 148452 372034 148464
rect 398834 148452 398840 148464
rect 398892 148452 398898 148504
rect 54938 148384 54944 148436
rect 54996 148424 55002 148436
rect 113174 148424 113180 148436
rect 54996 148396 113180 148424
rect 54996 148384 55002 148396
rect 113174 148384 113180 148396
rect 113232 148384 113238 148436
rect 370314 148384 370320 148436
rect 370372 148424 370378 148436
rect 370372 148396 373994 148424
rect 370372 148384 370378 148396
rect 52178 148316 52184 148368
rect 52236 148356 52242 148368
rect 110506 148356 110512 148368
rect 52236 148328 110512 148356
rect 52236 148316 52242 148328
rect 110506 148316 110512 148328
rect 110564 148316 110570 148368
rect 213454 148316 213460 148368
rect 213512 148356 213518 148368
rect 215938 148356 215944 148368
rect 213512 148328 215944 148356
rect 213512 148316 213518 148328
rect 215938 148316 215944 148328
rect 215996 148356 216002 148368
rect 271874 148356 271880 148368
rect 215996 148328 271880 148356
rect 215996 148316 216002 148328
rect 271874 148316 271880 148328
rect 271932 148316 271938 148368
rect 373966 148288 373994 148396
rect 380250 148384 380256 148436
rect 380308 148424 380314 148436
rect 423674 148424 423680 148436
rect 380308 148396 423680 148424
rect 380308 148384 380314 148396
rect 423674 148384 423680 148396
rect 423732 148384 423738 148436
rect 376386 148316 376392 148368
rect 376444 148356 376450 148368
rect 434714 148356 434720 148368
rect 376444 148328 380480 148356
rect 376444 148316 376450 148328
rect 377674 148288 377680 148300
rect 373966 148260 377680 148288
rect 377674 148248 377680 148260
rect 377732 148288 377738 148300
rect 380250 148288 380256 148300
rect 377732 148260 380256 148288
rect 377732 148248 377738 148260
rect 380250 148248 380256 148260
rect 380308 148248 380314 148300
rect 380452 148288 380480 148328
rect 386386 148328 434720 148356
rect 386386 148288 386414 148328
rect 434714 148316 434720 148328
rect 434772 148316 434778 148368
rect 380452 148260 386414 148288
rect 213178 147636 213184 147688
rect 213236 147676 213242 147688
rect 215018 147676 215024 147688
rect 213236 147648 215024 147676
rect 213236 147636 213242 147648
rect 215018 147636 215024 147648
rect 215076 147636 215082 147688
rect 374362 147636 374368 147688
rect 374420 147676 374426 147688
rect 376386 147676 376392 147688
rect 374420 147648 376392 147676
rect 374420 147636 374426 147648
rect 376386 147636 376392 147648
rect 376444 147636 376450 147688
rect 379422 147636 379428 147688
rect 379480 147676 379486 147688
rect 379882 147676 379888 147688
rect 379480 147648 379888 147676
rect 379480 147636 379486 147648
rect 379882 147636 379888 147648
rect 379940 147636 379946 147688
rect 59722 147568 59728 147620
rect 59780 147608 59786 147620
rect 107654 147608 107660 147620
rect 59780 147580 107660 147608
rect 59780 147568 59786 147580
rect 107654 147568 107660 147580
rect 107712 147568 107718 147620
rect 379330 147568 379336 147620
rect 379388 147608 379394 147620
rect 426526 147608 426532 147620
rect 379388 147580 426532 147608
rect 379388 147568 379394 147580
rect 426526 147568 426532 147580
rect 426584 147568 426590 147620
rect 57054 147500 57060 147552
rect 57112 147540 57118 147552
rect 104894 147540 104900 147552
rect 57112 147512 104900 147540
rect 57112 147500 57118 147512
rect 104894 147500 104900 147512
rect 104952 147500 104958 147552
rect 378962 147364 378968 147416
rect 379020 147404 379026 147416
rect 379330 147404 379336 147416
rect 379020 147376 379336 147404
rect 379020 147364 379026 147376
rect 379330 147364 379336 147376
rect 379388 147364 379394 147416
rect 213454 146276 213460 146328
rect 213512 146316 213518 146328
rect 213512 146288 274680 146316
rect 213512 146276 213518 146288
rect 47762 146208 47768 146260
rect 47820 146248 47826 146260
rect 51810 146248 51816 146260
rect 47820 146220 51816 146248
rect 47820 146208 47826 146220
rect 51810 146208 51816 146220
rect 51868 146208 51874 146260
rect 56226 146208 56232 146260
rect 56284 146248 56290 146260
rect 57974 146248 57980 146260
rect 56284 146220 57980 146248
rect 56284 146208 56290 146220
rect 57974 146208 57980 146220
rect 58032 146208 58038 146260
rect 58894 146208 58900 146260
rect 58952 146248 58958 146260
rect 59814 146248 59820 146260
rect 58952 146220 59820 146248
rect 58952 146208 58958 146220
rect 59814 146208 59820 146220
rect 59872 146248 59878 146260
rect 102134 146248 102140 146260
rect 59872 146220 102140 146248
rect 59872 146208 59878 146220
rect 102134 146208 102140 146220
rect 102192 146208 102198 146260
rect 179046 146208 179052 146260
rect 179104 146248 179110 146260
rect 197538 146248 197544 146260
rect 179104 146220 197544 146248
rect 179104 146208 179110 146220
rect 197538 146208 197544 146220
rect 197596 146208 197602 146260
rect 219066 146208 219072 146260
rect 219124 146248 219130 146260
rect 255314 146248 255320 146260
rect 219124 146220 255320 146248
rect 219124 146208 219130 146220
rect 255314 146208 255320 146220
rect 255372 146208 255378 146260
rect 274652 146248 274680 146288
rect 274818 146248 274824 146260
rect 274652 146220 274824 146248
rect 274818 146208 274824 146220
rect 274876 146248 274882 146260
rect 356790 146248 356796 146260
rect 274876 146220 356796 146248
rect 274876 146208 274882 146220
rect 356790 146208 356796 146220
rect 356848 146208 356854 146260
rect 376202 146208 376208 146260
rect 376260 146248 376266 146260
rect 376846 146248 376852 146260
rect 376260 146220 376852 146248
rect 376260 146208 376266 146220
rect 376846 146208 376852 146220
rect 376904 146208 376910 146260
rect 377950 146208 377956 146260
rect 378008 146248 378014 146260
rect 411254 146248 411260 146260
rect 378008 146220 411260 146248
rect 378008 146208 378014 146220
rect 411254 146208 411260 146220
rect 411312 146208 411318 146260
rect 53098 146140 53104 146192
rect 53156 146180 53162 146192
rect 86954 146180 86960 146192
rect 53156 146152 86960 146180
rect 53156 146140 53162 146152
rect 86954 146140 86960 146152
rect 87012 146140 87018 146192
rect 179690 146140 179696 146192
rect 179748 146180 179754 146192
rect 197630 146180 197636 146192
rect 179748 146152 197636 146180
rect 179748 146140 179754 146152
rect 197630 146140 197636 146152
rect 197688 146140 197694 146192
rect 236638 146140 236644 146192
rect 236696 146180 236702 146192
rect 256694 146180 256700 146192
rect 236696 146152 256700 146180
rect 236696 146140 236702 146152
rect 256694 146140 256700 146152
rect 256752 146140 256758 146192
rect 276014 146140 276020 146192
rect 276072 146180 276078 146192
rect 356606 146180 356612 146192
rect 276072 146152 356612 146180
rect 276072 146140 276078 146152
rect 356606 146140 356612 146152
rect 356664 146140 356670 146192
rect 375834 146140 375840 146192
rect 375892 146180 375898 146192
rect 379054 146180 379060 146192
rect 375892 146152 379060 146180
rect 375892 146140 375898 146152
rect 379054 146140 379060 146152
rect 379112 146140 379118 146192
rect 379238 146140 379244 146192
rect 379296 146180 379302 146192
rect 411346 146180 411352 146192
rect 379296 146152 411352 146180
rect 379296 146140 379302 146152
rect 411346 146140 411352 146152
rect 411404 146140 411410 146192
rect 500218 146140 500224 146192
rect 500276 146180 500282 146192
rect 518066 146180 518072 146192
rect 500276 146152 518072 146180
rect 500276 146140 500282 146152
rect 518066 146140 518072 146152
rect 518124 146180 518130 146192
rect 518250 146180 518256 146192
rect 518124 146152 518256 146180
rect 518124 146140 518130 146152
rect 518250 146140 518256 146152
rect 518308 146140 518314 146192
rect 56962 146072 56968 146124
rect 57020 146112 57026 146124
rect 58986 146112 58992 146124
rect 57020 146084 58992 146112
rect 57020 146072 57026 146084
rect 58986 146072 58992 146084
rect 59044 146072 59050 146124
rect 59446 146072 59452 146124
rect 59504 146112 59510 146124
rect 88426 146112 88432 146124
rect 59504 146084 88432 146112
rect 59504 146072 59510 146084
rect 88426 146072 88432 146084
rect 88484 146072 88490 146124
rect 219802 146072 219808 146124
rect 219860 146112 219866 146124
rect 253934 146112 253940 146124
rect 219860 146084 253940 146112
rect 219860 146072 219866 146084
rect 253934 146072 253940 146084
rect 253992 146072 253998 146124
rect 338482 146072 338488 146124
rect 338540 146112 338546 146124
rect 357618 146112 357624 146124
rect 338540 146084 357624 146112
rect 338540 146072 338546 146084
rect 357618 146072 357624 146084
rect 357676 146072 357682 146124
rect 378594 146072 378600 146124
rect 378652 146112 378658 146124
rect 409874 146112 409880 146124
rect 378652 146084 409880 146112
rect 378652 146072 378658 146084
rect 409874 146072 409880 146084
rect 409932 146072 409938 146124
rect 498654 146072 498660 146124
rect 498712 146112 498718 146124
rect 517698 146112 517704 146124
rect 498712 146084 517704 146112
rect 498712 146072 498718 146084
rect 517698 146072 517704 146084
rect 517756 146072 517762 146124
rect 57974 146004 57980 146056
rect 58032 146044 58038 146056
rect 89806 146044 89812 146056
rect 58032 146016 89812 146044
rect 58032 146004 58038 146016
rect 89806 146004 89812 146016
rect 89864 146004 89870 146056
rect 219894 146004 219900 146056
rect 219952 146044 219958 146056
rect 252554 146044 252560 146056
rect 219952 146016 252560 146044
rect 219952 146004 219958 146016
rect 252554 146004 252560 146016
rect 252612 146004 252618 146056
rect 340230 146004 340236 146056
rect 340288 146044 340294 146056
rect 356882 146044 356888 146056
rect 340288 146016 356888 146044
rect 340288 146004 340294 146016
rect 356882 146004 356888 146016
rect 356940 146004 356946 146056
rect 376846 146004 376852 146056
rect 376904 146044 376910 146056
rect 408494 146044 408500 146056
rect 376904 146016 408500 146044
rect 376904 146004 376910 146016
rect 408494 146004 408500 146016
rect 408552 146004 408558 146056
rect 54846 145936 54852 145988
rect 54904 145976 54910 145988
rect 85574 145976 85580 145988
rect 54904 145948 85580 145976
rect 54904 145936 54910 145948
rect 85574 145936 85580 145948
rect 85632 145936 85638 145988
rect 219250 145936 219256 145988
rect 219308 145976 219314 145988
rect 251174 145976 251180 145988
rect 219308 145948 251180 145976
rect 219308 145936 219314 145948
rect 251174 145936 251180 145948
rect 251232 145936 251238 145988
rect 376478 145936 376484 145988
rect 376536 145976 376542 145988
rect 405734 145976 405740 145988
rect 376536 145948 405740 145976
rect 376536 145936 376542 145948
rect 405734 145936 405740 145948
rect 405792 145936 405798 145988
rect 58710 145868 58716 145920
rect 58768 145908 58774 145920
rect 84286 145908 84292 145920
rect 58768 145880 84292 145908
rect 58768 145868 58774 145880
rect 84286 145868 84292 145880
rect 84344 145868 84350 145920
rect 217962 145868 217968 145920
rect 218020 145908 218026 145920
rect 249794 145908 249800 145920
rect 218020 145880 249800 145908
rect 218020 145868 218026 145880
rect 249794 145868 249800 145880
rect 249852 145868 249858 145920
rect 374270 145868 374276 145920
rect 374328 145908 374334 145920
rect 403066 145908 403072 145920
rect 374328 145880 403072 145908
rect 374328 145868 374334 145880
rect 403066 145868 403072 145880
rect 403124 145868 403130 145920
rect 56502 145800 56508 145852
rect 56560 145840 56566 145852
rect 84194 145840 84200 145852
rect 56560 145812 84200 145840
rect 56560 145800 56566 145812
rect 84194 145800 84200 145812
rect 84252 145800 84258 145852
rect 219158 145800 219164 145852
rect 219216 145840 219222 145852
rect 248414 145840 248420 145852
rect 219216 145812 248420 145840
rect 219216 145800 219222 145812
rect 248414 145800 248420 145812
rect 248472 145800 248478 145852
rect 376570 145800 376576 145852
rect 376628 145840 376634 145852
rect 402974 145840 402980 145852
rect 376628 145812 402980 145840
rect 376628 145800 376634 145812
rect 402974 145800 402980 145812
rect 403032 145800 403038 145852
rect 48958 145732 48964 145784
rect 49016 145772 49022 145784
rect 54386 145772 54392 145784
rect 49016 145744 54392 145772
rect 49016 145732 49022 145744
rect 54386 145732 54392 145744
rect 54444 145772 54450 145784
rect 82814 145772 82820 145784
rect 54444 145744 82820 145772
rect 54444 145732 54450 145744
rect 82814 145732 82820 145744
rect 82872 145732 82878 145784
rect 215110 145732 215116 145784
rect 215168 145772 215174 145784
rect 244366 145772 244372 145784
rect 215168 145744 244372 145772
rect 215168 145732 215174 145744
rect 244366 145732 244372 145744
rect 244424 145732 244430 145784
rect 375190 145732 375196 145784
rect 375248 145772 375254 145784
rect 378502 145772 378508 145784
rect 375248 145744 378508 145772
rect 375248 145732 375254 145744
rect 378502 145732 378508 145744
rect 378560 145772 378566 145784
rect 404354 145772 404360 145784
rect 378560 145744 404360 145772
rect 378560 145732 378566 145744
rect 404354 145732 404360 145744
rect 404412 145732 404418 145784
rect 58986 145664 58992 145716
rect 59044 145704 59050 145716
rect 91186 145704 91192 145716
rect 59044 145676 91192 145704
rect 59044 145664 59050 145676
rect 91186 145664 91192 145676
rect 91244 145664 91250 145716
rect 216122 145664 216128 145716
rect 216180 145704 216186 145716
rect 244274 145704 244280 145716
rect 216180 145676 244280 145704
rect 216180 145664 216186 145676
rect 244274 145664 244280 145676
rect 244332 145664 244338 145716
rect 375282 145664 375288 145716
rect 375340 145704 375346 145716
rect 397454 145704 397460 145716
rect 375340 145676 397460 145704
rect 375340 145664 375346 145676
rect 397454 145664 397460 145676
rect 397512 145664 397518 145716
rect 57054 145596 57060 145648
rect 57112 145636 57118 145648
rect 91094 145636 91100 145648
rect 57112 145608 91100 145636
rect 57112 145596 57118 145608
rect 91094 145596 91100 145608
rect 91152 145596 91158 145648
rect 216582 145596 216588 145648
rect 216640 145636 216646 145648
rect 247034 145636 247040 145648
rect 216640 145608 247040 145636
rect 216640 145596 216646 145608
rect 247034 145596 247040 145608
rect 247092 145596 247098 145648
rect 280062 145596 280068 145648
rect 280120 145636 280126 145648
rect 356606 145636 356612 145648
rect 280120 145608 356612 145636
rect 280120 145596 280126 145608
rect 356606 145596 356612 145608
rect 356664 145636 356670 145648
rect 358814 145636 358820 145648
rect 356664 145608 358820 145636
rect 356664 145596 356670 145608
rect 358814 145596 358820 145608
rect 358872 145596 358878 145648
rect 378042 145596 378048 145648
rect 378100 145636 378106 145648
rect 378594 145636 378600 145648
rect 378100 145608 378600 145636
rect 378100 145596 378106 145608
rect 378594 145596 378600 145608
rect 378652 145596 378658 145648
rect 378778 145596 378784 145648
rect 378836 145636 378842 145648
rect 407206 145636 407212 145648
rect 378836 145608 407212 145636
rect 378836 145596 378842 145608
rect 407206 145596 407212 145608
rect 407264 145596 407270 145648
rect 517698 145596 517704 145648
rect 517756 145636 517762 145648
rect 580350 145636 580356 145648
rect 517756 145608 580356 145636
rect 517756 145596 517762 145608
rect 580350 145596 580356 145608
rect 580408 145596 580414 145648
rect 46198 145528 46204 145580
rect 46256 145568 46262 145580
rect 59814 145568 59820 145580
rect 46256 145540 59820 145568
rect 46256 145528 46262 145540
rect 59814 145528 59820 145540
rect 59872 145568 59878 145580
rect 93854 145568 93860 145580
rect 59872 145540 93860 145568
rect 59872 145528 59878 145540
rect 93854 145528 93860 145540
rect 93912 145528 93918 145580
rect 191742 145528 191748 145580
rect 191800 145568 191806 145580
rect 197998 145568 198004 145580
rect 191800 145540 198004 145568
rect 191800 145528 191806 145540
rect 197998 145528 198004 145540
rect 198056 145568 198062 145580
rect 204898 145568 204904 145580
rect 198056 145540 204904 145568
rect 198056 145528 198062 145540
rect 204898 145528 204904 145540
rect 204956 145528 204962 145580
rect 214650 145528 214656 145580
rect 214708 145568 214714 145580
rect 245654 145568 245660 145580
rect 214708 145540 245660 145568
rect 214708 145528 214714 145540
rect 245654 145528 245660 145540
rect 245712 145528 245718 145580
rect 351638 145528 351644 145580
rect 351696 145568 351702 145580
rect 358078 145568 358084 145580
rect 351696 145540 358084 145568
rect 351696 145528 351702 145540
rect 358078 145528 358084 145540
rect 358136 145568 358142 145580
rect 358722 145568 358728 145580
rect 358136 145540 358728 145568
rect 358136 145528 358142 145540
rect 358722 145528 358728 145540
rect 358780 145568 358786 145580
rect 510522 145568 510528 145580
rect 358780 145540 510528 145568
rect 358780 145528 358786 145540
rect 510522 145528 510528 145540
rect 510580 145528 510586 145580
rect 518250 145528 518256 145580
rect 518308 145568 518314 145580
rect 580258 145568 580264 145580
rect 518308 145540 580264 145568
rect 518308 145528 518314 145540
rect 580258 145528 580264 145540
rect 580316 145528 580322 145580
rect 51810 145460 51816 145512
rect 51868 145500 51874 145512
rect 77294 145500 77300 145512
rect 51868 145472 77300 145500
rect 51868 145460 51874 145472
rect 77294 145460 77300 145472
rect 77352 145460 77358 145512
rect 215386 145460 215392 145512
rect 215444 145500 215450 145512
rect 242894 145500 242900 145512
rect 215444 145472 242900 145500
rect 215444 145460 215450 145472
rect 242894 145460 242900 145472
rect 242952 145460 242958 145512
rect 378870 145460 378876 145512
rect 378928 145500 378934 145512
rect 396074 145500 396080 145512
rect 378928 145472 396080 145500
rect 378928 145460 378934 145472
rect 396074 145460 396080 145472
rect 396132 145460 396138 145512
rect 48130 145392 48136 145444
rect 48188 145432 48194 145444
rect 54570 145432 54576 145444
rect 48188 145404 54576 145432
rect 48188 145392 48194 145404
rect 54570 145392 54576 145404
rect 54628 145432 54634 145444
rect 75914 145432 75920 145444
rect 54628 145404 75920 145432
rect 54628 145392 54634 145404
rect 75914 145392 75920 145404
rect 75972 145392 75978 145444
rect 218606 145392 218612 145444
rect 218664 145432 218670 145444
rect 236086 145432 236092 145444
rect 218664 145404 236092 145432
rect 218664 145392 218670 145404
rect 236086 145392 236092 145404
rect 236144 145392 236150 145444
rect 376110 145392 376116 145444
rect 376168 145432 376174 145444
rect 376570 145432 376576 145444
rect 376168 145404 376576 145432
rect 376168 145392 376174 145404
rect 376570 145392 376576 145404
rect 376628 145392 376634 145444
rect 379054 145392 379060 145444
rect 379112 145432 379118 145444
rect 396166 145432 396172 145444
rect 379112 145404 396172 145432
rect 379112 145392 379118 145404
rect 396166 145392 396172 145404
rect 396224 145392 396230 145444
rect 46382 145324 46388 145376
rect 46440 145364 46446 145376
rect 54662 145364 54668 145376
rect 46440 145336 54668 145364
rect 46440 145324 46446 145336
rect 54662 145324 54668 145336
rect 54720 145364 54726 145376
rect 76006 145364 76012 145376
rect 54720 145336 76012 145364
rect 54720 145324 54726 145336
rect 76006 145324 76012 145336
rect 76064 145324 76070 145376
rect 216214 145324 216220 145376
rect 216272 145364 216278 145376
rect 218974 145364 218980 145376
rect 216272 145336 218980 145364
rect 216272 145324 216278 145336
rect 218974 145324 218980 145336
rect 219032 145364 219038 145376
rect 235994 145364 236000 145376
rect 219032 145336 236000 145364
rect 219032 145324 219038 145336
rect 235994 145324 236000 145336
rect 236052 145324 236058 145376
rect 378962 145324 378968 145376
rect 379020 145364 379026 145376
rect 393958 145364 393964 145376
rect 379020 145336 393964 145364
rect 379020 145324 379026 145336
rect 393958 145324 393964 145336
rect 394016 145324 394022 145376
rect 56134 145256 56140 145308
rect 56192 145296 56198 145308
rect 59446 145296 59452 145308
rect 56192 145268 59452 145296
rect 56192 145256 56198 145268
rect 59446 145256 59452 145268
rect 59504 145256 59510 145308
rect 251266 145296 251272 145308
rect 229066 145268 251272 145296
rect 217134 145120 217140 145172
rect 217192 145160 217198 145172
rect 229066 145160 229094 145268
rect 251266 145256 251272 145268
rect 251324 145256 251330 145308
rect 217192 145132 229094 145160
rect 217192 145120 217198 145132
rect 218514 145052 218520 145104
rect 218572 145092 218578 145104
rect 219066 145092 219072 145104
rect 218572 145064 219072 145092
rect 218572 145052 218578 145064
rect 219066 145052 219072 145064
rect 219124 145052 219130 145104
rect 215386 144984 215392 145036
rect 215444 145024 215450 145036
rect 216214 145024 216220 145036
rect 215444 144996 216220 145024
rect 215444 144984 215450 144996
rect 216214 144984 216220 144996
rect 216272 144984 216278 145036
rect 218790 144984 218796 145036
rect 218848 145024 218854 145036
rect 219894 145024 219900 145036
rect 218848 144996 219900 145024
rect 218848 144984 218854 144996
rect 219894 144984 219900 144996
rect 219952 144984 219958 145036
rect 215846 144916 215852 144968
rect 215904 144956 215910 144968
rect 216122 144956 216128 144968
rect 215904 144928 216128 144956
rect 215904 144916 215910 144928
rect 216122 144916 216128 144928
rect 216180 144916 216186 144968
rect 217042 144916 217048 144968
rect 217100 144956 217106 144968
rect 217962 144956 217968 144968
rect 217100 144928 217968 144956
rect 217100 144916 217106 144928
rect 217962 144916 217968 144928
rect 218020 144916 218026 144968
rect 218882 144916 218888 144968
rect 218940 144956 218946 144968
rect 219250 144956 219256 144968
rect 218940 144928 219256 144956
rect 218940 144916 218946 144928
rect 219250 144916 219256 144928
rect 219308 144916 219314 144968
rect 375098 144956 375104 144968
rect 373828 144928 375104 144956
rect 54478 144848 54484 144900
rect 54536 144888 54542 144900
rect 55950 144888 55956 144900
rect 54536 144860 55956 144888
rect 54536 144848 54542 144860
rect 55950 144848 55956 144860
rect 56008 144888 56014 144900
rect 56502 144888 56508 144900
rect 56008 144860 56508 144888
rect 56008 144848 56014 144860
rect 56502 144848 56508 144860
rect 56560 144848 56566 144900
rect 209590 144848 209596 144900
rect 209648 144888 209654 144900
rect 214558 144888 214564 144900
rect 209648 144860 214564 144888
rect 209648 144848 209654 144860
rect 214558 144848 214564 144860
rect 214616 144848 214622 144900
rect 372430 144848 372436 144900
rect 372488 144888 372494 144900
rect 373828 144888 373856 144928
rect 375098 144916 375104 144928
rect 375156 144956 375162 144968
rect 375282 144956 375288 144968
rect 375156 144928 375288 144956
rect 375156 144916 375162 144928
rect 375282 144916 375288 144928
rect 375340 144916 375346 144968
rect 372488 144860 373856 144888
rect 372488 144848 372494 144860
rect 373902 144848 373908 144900
rect 373960 144888 373966 144900
rect 378778 144888 378784 144900
rect 373960 144860 378784 144888
rect 373960 144848 373966 144860
rect 378778 144848 378784 144860
rect 378836 144848 378842 144900
rect 51994 144780 52000 144832
rect 52052 144820 52058 144832
rect 58710 144820 58716 144832
rect 52052 144792 58716 144820
rect 52052 144780 52058 144792
rect 58710 144780 58716 144792
rect 58768 144780 58774 144832
rect 213730 144780 213736 144832
rect 213788 144820 213794 144832
rect 216030 144820 216036 144832
rect 213788 144792 216036 144820
rect 213788 144780 213794 144792
rect 216030 144780 216036 144792
rect 216088 144820 216094 144832
rect 216582 144820 216588 144832
rect 216088 144792 216588 144820
rect 216088 144780 216094 144792
rect 216582 144780 216588 144792
rect 216640 144780 216646 144832
rect 374086 144780 374092 144832
rect 374144 144820 374150 144832
rect 378870 144820 378876 144832
rect 374144 144792 378876 144820
rect 374144 144780 374150 144792
rect 378870 144780 378876 144792
rect 378928 144780 378934 144832
rect 51902 144712 51908 144764
rect 51960 144752 51966 144764
rect 57054 144752 57060 144764
rect 51960 144724 57060 144752
rect 51960 144712 51966 144724
rect 57054 144712 57060 144724
rect 57112 144712 57118 144764
rect 213638 144712 213644 144764
rect 213696 144752 213702 144764
rect 214650 144752 214656 144764
rect 213696 144724 214656 144752
rect 213696 144712 213702 144724
rect 214650 144712 214656 144724
rect 214708 144712 214714 144764
rect 50338 144644 50344 144696
rect 50396 144684 50402 144696
rect 55858 144684 55864 144696
rect 50396 144656 55864 144684
rect 50396 144644 50402 144656
rect 55858 144644 55864 144656
rect 55916 144684 55922 144696
rect 56410 144684 56416 144696
rect 55916 144656 56416 144684
rect 55916 144644 55922 144656
rect 56410 144644 56416 144656
rect 56468 144644 56474 144696
rect 213546 144644 213552 144696
rect 213604 144684 213610 144696
rect 216122 144684 216128 144696
rect 213604 144656 216128 144684
rect 213604 144644 213610 144656
rect 216122 144644 216128 144656
rect 216180 144684 216186 144696
rect 216306 144684 216312 144696
rect 216180 144656 216312 144684
rect 216180 144644 216186 144656
rect 216306 144644 216312 144656
rect 216364 144644 216370 144696
rect 374270 144644 374276 144696
rect 374328 144684 374334 144696
rect 375190 144684 375196 144696
rect 374328 144656 375196 144684
rect 374328 144644 374334 144656
rect 375190 144644 375196 144656
rect 375248 144644 375254 144696
rect 49234 144576 49240 144628
rect 49292 144616 49298 144628
rect 58618 144616 58624 144628
rect 49292 144588 58624 144616
rect 49292 144576 49298 144588
rect 58618 144576 58624 144588
rect 58676 144576 58682 144628
rect 212074 144576 212080 144628
rect 212132 144616 212138 144628
rect 215018 144616 215024 144628
rect 212132 144588 215024 144616
rect 212132 144576 212138 144588
rect 215018 144576 215024 144588
rect 215076 144576 215082 144628
rect 520182 79976 520188 80028
rect 520240 80016 520246 80028
rect 580442 80016 580448 80028
rect 520240 79988 580448 80016
rect 520240 79976 520246 79988
rect 580442 79976 580448 79988
rect 580500 79976 580506 80028
rect 207658 70320 207664 70372
rect 207716 70360 207722 70372
rect 216674 70360 216680 70372
rect 207716 70332 216680 70360
rect 207716 70320 207722 70332
rect 216674 70320 216680 70332
rect 216732 70320 216738 70372
rect 365070 70320 365076 70372
rect 365128 70360 365134 70372
rect 376938 70360 376944 70372
rect 365128 70332 376944 70360
rect 365128 70320 365134 70332
rect 376938 70320 376944 70332
rect 376996 70320 377002 70372
rect 46842 68960 46848 69012
rect 46900 69000 46906 69012
rect 56870 69000 56876 69012
rect 46900 68972 56876 69000
rect 46900 68960 46906 68972
rect 56870 68960 56876 68972
rect 56928 68960 56934 69012
rect 358078 68416 358084 68468
rect 358136 68456 358142 68468
rect 358722 68456 358728 68468
rect 358136 68428 358728 68456
rect 358136 68416 358142 68428
rect 358722 68416 358728 68428
rect 358780 68456 358786 68468
rect 358780 68428 364334 68456
rect 358780 68416 358786 68428
rect 364306 68320 364334 68428
rect 376938 68320 376944 68332
rect 364306 68292 376944 68320
rect 376938 68280 376944 68292
rect 376996 68280 377002 68332
rect 204898 67600 204904 67652
rect 204956 67640 204962 67652
rect 216674 67640 216680 67652
rect 204956 67612 216680 67640
rect 204956 67600 204962 67612
rect 216674 67600 216680 67612
rect 216732 67600 216738 67652
rect 218790 61072 218796 61124
rect 218848 61112 218854 61124
rect 219066 61112 219072 61124
rect 218848 61084 219072 61112
rect 218848 61072 218854 61084
rect 219066 61072 219072 61084
rect 219124 61072 219130 61124
rect 379054 59712 379060 59764
rect 379112 59752 379118 59764
rect 397086 59752 397092 59764
rect 379112 59724 397092 59752
rect 379112 59712 379118 59724
rect 397086 59712 397092 59724
rect 397144 59712 397150 59764
rect 218606 59644 218612 59696
rect 218664 59684 218670 59696
rect 237098 59684 237104 59696
rect 218664 59656 237104 59684
rect 218664 59644 218670 59656
rect 237098 59644 237104 59656
rect 237156 59644 237162 59696
rect 378870 59644 378876 59696
rect 378928 59684 378934 59696
rect 396074 59684 396080 59696
rect 378928 59656 396080 59684
rect 378928 59644 378934 59656
rect 396074 59644 396080 59656
rect 396132 59644 396138 59696
rect 54570 59576 54576 59628
rect 54628 59616 54634 59628
rect 77110 59616 77116 59628
rect 54628 59588 77116 59616
rect 54628 59576 54634 59588
rect 77110 59576 77116 59588
rect 77168 59576 77174 59628
rect 218514 59576 218520 59628
rect 218572 59616 218578 59628
rect 255866 59616 255872 59628
rect 218572 59588 255872 59616
rect 218572 59576 218578 59588
rect 255866 59576 255872 59588
rect 255924 59576 255930 59628
rect 378962 59576 378968 59628
rect 379020 59616 379026 59628
rect 418154 59616 418160 59628
rect 379020 59588 418160 59616
rect 379020 59576 379026 59588
rect 418154 59576 418160 59588
rect 418212 59576 418218 59628
rect 54386 59508 54392 59560
rect 54444 59548 54450 59560
rect 83090 59548 83096 59560
rect 54444 59520 83096 59548
rect 54444 59508 54450 59520
rect 83090 59508 83096 59520
rect 83148 59508 83154 59560
rect 217870 59508 217876 59560
rect 217928 59548 217934 59560
rect 256970 59548 256976 59560
rect 217928 59520 256976 59548
rect 217928 59508 217934 59520
rect 256970 59508 256976 59520
rect 257028 59508 257034 59560
rect 375926 59508 375932 59560
rect 375984 59548 375990 59560
rect 416958 59548 416964 59560
rect 375984 59520 416964 59548
rect 375984 59508 375990 59520
rect 416958 59508 416964 59520
rect 417016 59508 417022 59560
rect 55030 59440 55036 59492
rect 55088 59480 55094 59492
rect 99466 59480 99472 59492
rect 55088 59452 99472 59480
rect 55088 59440 55094 59452
rect 99466 59440 99472 59452
rect 99524 59440 99530 59492
rect 219342 59440 219348 59492
rect 219400 59480 219406 59492
rect 263870 59480 263876 59492
rect 219400 59452 263876 59480
rect 219400 59440 219406 59452
rect 263870 59440 263876 59452
rect 263928 59440 263934 59492
rect 377674 59440 377680 59492
rect 377732 59480 377738 59492
rect 423950 59480 423956 59492
rect 377732 59452 423956 59480
rect 377732 59440 377738 59452
rect 423950 59440 423956 59452
rect 424008 59440 424014 59492
rect 49510 59372 49516 59424
rect 49568 59412 49574 59424
rect 113542 59412 113548 59424
rect 49568 59384 113548 59412
rect 49568 59372 49574 59384
rect 113542 59372 113548 59384
rect 113600 59372 113606 59424
rect 214742 59372 214748 59424
rect 214800 59412 214806 59424
rect 261754 59412 261760 59424
rect 214800 59384 261760 59412
rect 214800 59372 214806 59384
rect 261754 59372 261760 59384
rect 261812 59372 261818 59424
rect 362218 59372 362224 59424
rect 362276 59412 362282 59424
rect 418430 59412 418436 59424
rect 362276 59384 418436 59412
rect 362276 59372 362282 59384
rect 418430 59372 418436 59384
rect 418488 59372 418494 59424
rect 55950 59304 55956 59356
rect 56008 59344 56014 59356
rect 84194 59344 84200 59356
rect 56008 59316 84200 59344
rect 56008 59304 56014 59316
rect 84194 59304 84200 59316
rect 84252 59304 84258 59356
rect 217962 59304 217968 59356
rect 218020 59344 218026 59356
rect 358078 59344 358084 59356
rect 218020 59316 358084 59344
rect 218020 59304 218026 59316
rect 358078 59304 358084 59316
rect 358136 59304 358142 59356
rect 59814 59236 59820 59288
rect 59872 59276 59878 59288
rect 94498 59276 94504 59288
rect 59872 59248 94504 59276
rect 59872 59236 59878 59248
rect 94498 59236 94504 59248
rect 94556 59236 94562 59288
rect 375190 59236 375196 59288
rect 375248 59276 375254 59288
rect 403066 59276 403072 59288
rect 375248 59248 403072 59276
rect 375248 59236 375254 59248
rect 403066 59236 403072 59248
rect 403124 59236 403130 59288
rect 57790 59168 57796 59220
rect 57848 59208 57854 59220
rect 95878 59208 95884 59220
rect 57848 59180 95884 59208
rect 57848 59168 57854 59180
rect 95878 59168 95884 59180
rect 95936 59168 95942 59220
rect 214834 59168 214840 59220
rect 214892 59208 214898 59220
rect 260650 59208 260656 59220
rect 214892 59180 260656 59208
rect 214892 59168 214898 59180
rect 260650 59168 260656 59180
rect 260708 59168 260714 59220
rect 379606 59168 379612 59220
rect 379664 59208 379670 59220
rect 419442 59208 419448 59220
rect 379664 59180 419448 59208
rect 379664 59168 379670 59180
rect 419442 59168 419448 59180
rect 419500 59168 419506 59220
rect 59078 59100 59084 59152
rect 59136 59140 59142 59152
rect 96982 59140 96988 59152
rect 59136 59112 96988 59140
rect 59136 59100 59142 59112
rect 96982 59100 96988 59112
rect 97040 59100 97046 59152
rect 215754 59100 215760 59152
rect 215812 59140 215818 59152
rect 262766 59140 262772 59152
rect 215812 59112 262772 59140
rect 215812 59100 215818 59112
rect 262766 59100 262772 59112
rect 262824 59100 262830 59152
rect 279234 59100 279240 59152
rect 279292 59140 279298 59152
rect 356606 59140 356612 59152
rect 279292 59112 356612 59140
rect 279292 59100 279298 59112
rect 356606 59100 356612 59112
rect 356664 59100 356670 59152
rect 376662 59100 376668 59152
rect 376720 59140 376726 59152
rect 420638 59140 420644 59152
rect 376720 59112 420644 59140
rect 376720 59100 376726 59112
rect 420638 59100 420644 59112
rect 420696 59100 420702 59152
rect 58894 59032 58900 59084
rect 58952 59072 58958 59084
rect 102778 59072 102784 59084
rect 58952 59044 102784 59072
rect 58952 59032 58958 59044
rect 102778 59032 102784 59044
rect 102836 59032 102842 59084
rect 205542 59032 205548 59084
rect 205600 59072 205606 59084
rect 290918 59072 290924 59084
rect 205600 59044 290924 59072
rect 205600 59032 205606 59044
rect 290918 59032 290924 59044
rect 290976 59032 290982 59084
rect 376294 59032 376300 59084
rect 376352 59072 376358 59084
rect 421742 59072 421748 59084
rect 376352 59044 421748 59072
rect 376352 59032 376358 59044
rect 421742 59032 421748 59044
rect 421800 59032 421806 59084
rect 56042 58964 56048 59016
rect 56100 59004 56106 59016
rect 101766 59004 101772 59016
rect 56100 58976 101772 59004
rect 56100 58964 56106 58976
rect 101766 58964 101772 58976
rect 101824 58964 101830 59016
rect 208946 58964 208952 59016
rect 209004 59004 209010 59016
rect 298462 59004 298468 59016
rect 209004 58976 298468 59004
rect 209004 58964 209010 58976
rect 298462 58964 298468 58976
rect 298520 58964 298526 59016
rect 379698 58964 379704 59016
rect 379756 59004 379762 59016
rect 425238 59004 425244 59016
rect 379756 58976 425244 59004
rect 379756 58964 379762 58976
rect 425238 58964 425244 58976
rect 425296 58964 425302 59016
rect 55858 58896 55864 58948
rect 55916 58936 55922 58948
rect 103882 58936 103888 58948
rect 55916 58908 103888 58936
rect 55916 58896 55922 58908
rect 103882 58896 103888 58908
rect 103940 58896 103946 58948
rect 215202 58896 215208 58948
rect 215260 58936 215266 58948
rect 313366 58936 313372 58948
rect 215260 58908 313372 58936
rect 215260 58896 215266 58908
rect 313366 58896 313372 58908
rect 313424 58896 313430 58948
rect 373258 58896 373264 58948
rect 373316 58936 373322 58948
rect 423490 58936 423496 58948
rect 373316 58908 423496 58936
rect 373316 58896 373322 58908
rect 423490 58896 423496 58908
rect 423548 58896 423554 58948
rect 54754 58828 54760 58880
rect 54812 58868 54818 58880
rect 111150 58868 111156 58880
rect 54812 58840 111156 58868
rect 54812 58828 54818 58840
rect 111150 58828 111156 58840
rect 111208 58828 111214 58880
rect 206830 58828 206836 58880
rect 206888 58868 206894 58880
rect 305914 58868 305920 58880
rect 206888 58840 305920 58868
rect 206888 58828 206894 58840
rect 305914 58828 305920 58840
rect 305972 58828 305978 58880
rect 363598 58828 363604 58880
rect 363656 58868 363662 58880
rect 425974 58868 425980 58880
rect 363656 58840 425980 58868
rect 363656 58828 363662 58840
rect 425974 58828 425980 58840
rect 426032 58828 426038 58880
rect 42610 58760 42616 58812
rect 42668 58800 42674 58812
rect 115934 58800 115940 58812
rect 42668 58772 115940 58800
rect 42668 58760 42674 58772
rect 115934 58760 115940 58772
rect 115992 58760 115998 58812
rect 201402 58760 201408 58812
rect 201460 58800 201466 58812
rect 318426 58800 318432 58812
rect 201460 58772 318432 58800
rect 201460 58760 201466 58772
rect 318426 58760 318432 58772
rect 318484 58760 318490 58812
rect 366450 58760 366456 58812
rect 366508 58800 366514 58812
rect 465902 58800 465908 58812
rect 366508 58772 465908 58800
rect 366508 58760 366514 58772
rect 465902 58760 465908 58772
rect 465960 58760 465966 58812
rect 50062 58692 50068 58744
rect 50120 58732 50126 58744
rect 148502 58732 148508 58744
rect 50120 58704 148508 58732
rect 50120 58692 50126 58704
rect 148502 58692 148508 58704
rect 148560 58692 148566 58744
rect 202782 58692 202788 58744
rect 202840 58732 202846 58744
rect 325878 58732 325884 58744
rect 202840 58704 325884 58732
rect 202840 58692 202846 58704
rect 325878 58692 325884 58704
rect 325936 58692 325942 58744
rect 358630 58692 358636 58744
rect 358688 58732 358694 58744
rect 485958 58732 485964 58744
rect 358688 58704 485964 58732
rect 358688 58692 358694 58704
rect 485958 58692 485964 58704
rect 486016 58692 486022 58744
rect 53558 58624 53564 58676
rect 53616 58664 53622 58676
rect 150894 58664 150900 58676
rect 53616 58636 150900 58664
rect 53616 58624 53622 58636
rect 150894 58624 150900 58636
rect 150952 58624 150958 58676
rect 219250 58624 219256 58676
rect 219308 58664 219314 58676
rect 428182 58664 428188 58676
rect 219308 58636 428188 58664
rect 219308 58624 219314 58636
rect 428182 58624 428188 58636
rect 428240 58624 428246 58676
rect 216398 58556 216404 58608
rect 216456 58596 216462 58608
rect 259454 58596 259460 58608
rect 216456 58568 259460 58596
rect 216456 58556 216462 58568
rect 259454 58556 259460 58568
rect 259512 58556 259518 58608
rect 376110 58556 376116 58608
rect 376168 58596 376174 58608
rect 404170 58596 404176 58608
rect 376168 58568 404176 58596
rect 376168 58556 376174 58568
rect 404170 58556 404176 58568
rect 404228 58556 404234 58608
rect 57882 57876 57888 57928
rect 57940 57916 57946 57928
rect 204898 57916 204904 57928
rect 57940 57888 204904 57916
rect 57940 57876 57946 57888
rect 204898 57876 204904 57888
rect 204956 57876 204962 57928
rect 210970 57876 210976 57928
rect 211028 57916 211034 57928
rect 323302 57916 323308 57928
rect 211028 57888 323308 57916
rect 211028 57876 211034 57888
rect 323302 57876 323308 57888
rect 323360 57876 323366 57928
rect 343174 57876 343180 57928
rect 343232 57916 343238 57928
rect 357526 57916 357532 57928
rect 343232 57888 357532 57916
rect 343232 57876 343238 57888
rect 357526 57876 357532 57888
rect 357584 57876 357590 57928
rect 364978 57876 364984 57928
rect 365036 57916 365042 57928
rect 478414 57916 478420 57928
rect 365036 57888 478420 57916
rect 365036 57876 365042 57888
rect 478414 57876 478420 57888
rect 478472 57876 478478 57928
rect 503346 57876 503352 57928
rect 503404 57916 503410 57928
rect 517606 57916 517612 57928
rect 503404 57888 517612 57916
rect 503404 57876 503410 57888
rect 517606 57876 517612 57888
rect 517664 57876 517670 57928
rect 52362 57808 52368 57860
rect 52420 57848 52426 57860
rect 145558 57848 145564 57860
rect 52420 57820 145564 57848
rect 52420 57808 52426 57820
rect 145558 57808 145564 57820
rect 145616 57808 145622 57860
rect 183278 57808 183284 57860
rect 183336 57848 183342 57860
rect 197446 57848 197452 57860
rect 183336 57820 197452 57848
rect 183336 57808 183342 57820
rect 197446 57808 197452 57820
rect 197504 57808 197510 57860
rect 212350 57808 212356 57860
rect 212408 57848 212414 57860
rect 315758 57848 315764 57860
rect 212408 57820 315764 57848
rect 212408 57808 212414 57820
rect 315758 57808 315764 57820
rect 315816 57808 315822 57860
rect 343450 57808 343456 57860
rect 343508 57848 343514 57860
rect 356698 57848 356704 57860
rect 343508 57820 356704 57848
rect 343508 57808 343514 57820
rect 356698 57808 356704 57820
rect 356756 57808 356762 57860
rect 360838 57808 360844 57860
rect 360896 57848 360902 57860
rect 443454 57848 443460 57860
rect 360896 57820 443460 57848
rect 360896 57808 360902 57820
rect 443454 57808 443460 57820
rect 443512 57808 443518 57860
rect 503254 57808 503260 57860
rect 503312 57848 503318 57860
rect 517514 57848 517520 57860
rect 503312 57820 517520 57848
rect 503312 57808 503318 57820
rect 517514 57808 517520 57820
rect 517572 57808 517578 57860
rect 44082 57740 44088 57792
rect 44140 57780 44146 57792
rect 123478 57780 123484 57792
rect 44140 57752 123484 57780
rect 44140 57740 44146 57752
rect 123478 57740 123484 57752
rect 123536 57740 123542 57792
rect 183462 57740 183468 57792
rect 183520 57780 183526 57792
rect 197354 57780 197360 57792
rect 183520 57752 197360 57780
rect 183520 57740 183526 57752
rect 197354 57740 197360 57752
rect 197412 57740 197418 57792
rect 218698 57740 218704 57792
rect 218756 57780 218762 57792
rect 320910 57780 320916 57792
rect 218756 57752 320916 57780
rect 218756 57740 218762 57752
rect 320910 57740 320916 57752
rect 320968 57740 320974 57792
rect 358170 57740 358176 57792
rect 358228 57780 358234 57792
rect 440878 57780 440884 57792
rect 358228 57752 440884 57780
rect 358228 57740 358234 57752
rect 440878 57740 440884 57752
rect 440936 57740 440942 57792
rect 52822 57672 52828 57724
rect 52880 57712 52886 57724
rect 130838 57712 130844 57724
rect 52880 57684 130844 57712
rect 52880 57672 52886 57684
rect 130838 57672 130844 57684
rect 130896 57672 130902 57724
rect 208302 57672 208308 57724
rect 208360 57712 208366 57724
rect 308490 57712 308496 57724
rect 208360 57684 308496 57712
rect 208360 57672 208366 57684
rect 308490 57672 308496 57684
rect 308548 57672 308554 57724
rect 363690 57672 363696 57724
rect 363748 57712 363754 57724
rect 445846 57712 445852 57724
rect 363748 57684 445852 57712
rect 363748 57672 363754 57684
rect 445846 57672 445852 57684
rect 445904 57672 445910 57724
rect 54938 57604 54944 57656
rect 54996 57644 55002 57656
rect 54996 57616 58020 57644
rect 54996 57604 55002 57616
rect 57238 57536 57244 57588
rect 57296 57576 57302 57588
rect 57882 57576 57888 57588
rect 57296 57548 57888 57576
rect 57296 57536 57302 57548
rect 57882 57536 57888 57548
rect 57940 57536 57946 57588
rect 57992 57576 58020 57616
rect 58066 57604 58072 57656
rect 58124 57644 58130 57656
rect 133230 57644 133236 57656
rect 58124 57616 133236 57644
rect 58124 57604 58130 57616
rect 133230 57604 133236 57616
rect 133288 57604 133294 57656
rect 216490 57604 216496 57656
rect 216548 57644 216554 57656
rect 310974 57644 310980 57656
rect 216548 57616 310980 57644
rect 216548 57604 216554 57616
rect 310974 57604 310980 57616
rect 311032 57604 311038 57656
rect 374638 57604 374644 57656
rect 374696 57644 374702 57656
rect 450998 57644 451004 57656
rect 374696 57616 451004 57644
rect 374696 57604 374702 57616
rect 450998 57604 451004 57616
rect 451056 57604 451062 57656
rect 112070 57576 112076 57588
rect 57992 57548 112076 57576
rect 112070 57536 112076 57548
rect 112128 57536 112134 57588
rect 213822 57536 213828 57588
rect 213880 57576 213886 57588
rect 303430 57576 303436 57588
rect 213880 57548 303436 57576
rect 213880 57536 213886 57548
rect 303430 57536 303436 57548
rect 303488 57536 303494 57588
rect 362310 57536 362316 57588
rect 362368 57576 362374 57588
rect 438486 57576 438492 57588
rect 362368 57548 438492 57576
rect 362368 57536 362374 57548
rect 438486 57536 438492 57548
rect 438544 57536 438550 57588
rect 39942 57468 39948 57520
rect 40000 57508 40006 57520
rect 90726 57508 90732 57520
rect 40000 57480 90732 57508
rect 40000 57468 40006 57480
rect 90726 57468 90732 57480
rect 90784 57468 90790 57520
rect 211062 57468 211068 57520
rect 211120 57508 211126 57520
rect 295886 57508 295892 57520
rect 211120 57480 295892 57508
rect 211120 57468 211126 57480
rect 295886 57468 295892 57480
rect 295944 57468 295950 57520
rect 371878 57468 371884 57520
rect 371936 57508 371942 57520
rect 435910 57508 435916 57520
rect 371936 57480 435916 57508
rect 371936 57468 371942 57480
rect 435910 57468 435916 57480
rect 435968 57468 435974 57520
rect 55122 57400 55128 57452
rect 55180 57440 55186 57452
rect 98086 57440 98092 57452
rect 55180 57412 98092 57440
rect 55180 57400 55186 57412
rect 98086 57400 98092 57412
rect 98144 57400 98150 57452
rect 218330 57400 218336 57452
rect 218388 57440 218394 57452
rect 300854 57440 300860 57452
rect 218388 57412 300860 57440
rect 218388 57400 218394 57412
rect 300854 57400 300860 57412
rect 300912 57400 300918 57452
rect 370590 57400 370596 57452
rect 370648 57440 370654 57452
rect 433518 57440 433524 57452
rect 370648 57412 433524 57440
rect 370648 57400 370654 57412
rect 433518 57400 433524 57412
rect 433576 57400 433582 57452
rect 53650 57332 53656 57384
rect 53708 57372 53714 57384
rect 88334 57372 88340 57384
rect 53708 57344 88340 57372
rect 53708 57332 53714 57344
rect 88334 57332 88340 57344
rect 88392 57332 88398 57384
rect 212442 57332 212448 57384
rect 212500 57372 212506 57384
rect 293310 57372 293316 57384
rect 212500 57344 293316 57372
rect 212500 57332 212506 57344
rect 293310 57332 293316 57344
rect 293368 57332 293374 57384
rect 376018 57332 376024 57384
rect 376076 57372 376082 57384
rect 430942 57372 430948 57384
rect 376076 57344 430948 57372
rect 376076 57332 376082 57344
rect 430942 57332 430948 57344
rect 431000 57332 431006 57384
rect 55490 57264 55496 57316
rect 55548 57304 55554 57316
rect 58066 57304 58072 57316
rect 55548 57276 58072 57304
rect 55548 57264 55554 57276
rect 58066 57264 58072 57276
rect 58124 57264 58130 57316
rect 59262 57264 59268 57316
rect 59320 57304 59326 57316
rect 93670 57304 93676 57316
rect 59320 57276 93676 57304
rect 59320 57264 59326 57276
rect 93670 57264 93676 57276
rect 93728 57264 93734 57316
rect 215294 57264 215300 57316
rect 215352 57304 215358 57316
rect 287606 57304 287612 57316
rect 215352 57276 287612 57304
rect 215352 57264 215358 57276
rect 287606 57264 287612 57276
rect 287664 57264 287670 57316
rect 370498 57264 370504 57316
rect 370556 57304 370562 57316
rect 416038 57304 416044 57316
rect 370556 57276 416044 57304
rect 370556 57264 370562 57276
rect 416038 57264 416044 57276
rect 416096 57264 416102 57316
rect 51810 57196 51816 57248
rect 51868 57236 51874 57248
rect 78214 57236 78220 57248
rect 51868 57208 78220 57236
rect 51868 57196 51874 57208
rect 78214 57196 78220 57208
rect 78272 57196 78278 57248
rect 218790 57196 218796 57248
rect 218848 57236 218854 57248
rect 265894 57236 265900 57248
rect 218848 57208 265900 57236
rect 218848 57196 218854 57208
rect 265894 57196 265900 57208
rect 265952 57196 265958 57248
rect 379146 57196 379152 57248
rect 379204 57236 379210 57248
rect 415486 57236 415492 57248
rect 379204 57208 415492 57236
rect 379204 57196 379210 57208
rect 415486 57196 415492 57208
rect 415544 57196 415550 57248
rect 54662 57128 54668 57180
rect 54720 57168 54726 57180
rect 76006 57168 76012 57180
rect 54720 57140 76012 57168
rect 54720 57128 54726 57140
rect 76006 57128 76012 57140
rect 76064 57128 76070 57180
rect 58710 56516 58716 56568
rect 58768 56556 58774 56568
rect 85390 56556 85396 56568
rect 58768 56528 85396 56556
rect 58768 56516 58774 56528
rect 85390 56516 85396 56528
rect 85448 56516 85454 56568
rect 214926 56516 214932 56568
rect 214984 56556 214990 56568
rect 241606 56556 241612 56568
rect 214984 56528 241612 56556
rect 214984 56516 214990 56528
rect 241606 56516 241612 56528
rect 241664 56516 241670 56568
rect 375006 56516 375012 56568
rect 375064 56556 375070 56568
rect 401686 56556 401692 56568
rect 375064 56528 401692 56556
rect 375064 56516 375070 56528
rect 401686 56516 401692 56528
rect 401744 56516 401750 56568
rect 53190 56448 53196 56500
rect 53248 56488 53254 56500
rect 113174 56488 113180 56500
rect 53248 56460 113180 56488
rect 53248 56448 53254 56460
rect 113174 56448 113180 56460
rect 113232 56448 113238 56500
rect 215662 56448 215668 56500
rect 215720 56488 215726 56500
rect 239214 56488 239220 56500
rect 215720 56460 239220 56488
rect 215720 56448 215726 56460
rect 239214 56448 239220 56460
rect 239272 56448 239278 56500
rect 374546 56448 374552 56500
rect 374604 56488 374610 56500
rect 438302 56488 438308 56500
rect 374604 56460 438308 56488
rect 374604 56448 374610 56460
rect 438302 56448 438308 56460
rect 438360 56448 438366 56500
rect 59906 56380 59912 56432
rect 59964 56420 59970 56432
rect 108022 56420 108028 56432
rect 59964 56392 108028 56420
rect 59964 56380 59970 56392
rect 108022 56380 108028 56392
rect 108080 56380 108086 56432
rect 218974 56380 218980 56432
rect 219032 56420 219038 56432
rect 235994 56420 236000 56432
rect 219032 56392 236000 56420
rect 219032 56380 219038 56392
rect 235994 56380 236000 56392
rect 236052 56380 236058 56432
rect 372246 56380 372252 56432
rect 372304 56420 372310 56432
rect 435726 56420 435732 56432
rect 372304 56392 435732 56420
rect 372304 56380 372310 56392
rect 435726 56380 435732 56392
rect 435784 56380 435790 56432
rect 59170 56312 59176 56364
rect 59228 56352 59234 56364
rect 107378 56352 107384 56364
rect 59228 56324 107384 56352
rect 59228 56312 59234 56324
rect 107378 56312 107384 56324
rect 107436 56312 107442 56364
rect 215018 56312 215024 56364
rect 215076 56352 215082 56364
rect 271230 56352 271236 56364
rect 215076 56324 271236 56352
rect 215076 56312 215082 56324
rect 271230 56312 271236 56324
rect 271288 56312 271294 56364
rect 376386 56312 376392 56364
rect 376444 56352 376450 56364
rect 433334 56352 433340 56364
rect 376444 56324 433340 56352
rect 376444 56312 376450 56324
rect 433334 56312 433340 56324
rect 433392 56312 433398 56364
rect 59998 56244 60004 56296
rect 60056 56284 60062 56296
rect 106366 56284 106372 56296
rect 60056 56256 106372 56284
rect 60056 56244 60062 56256
rect 106366 56244 106372 56256
rect 106424 56244 106430 56296
rect 219526 56244 219532 56296
rect 219584 56284 219590 56296
rect 268470 56284 268476 56296
rect 219584 56256 268476 56284
rect 219584 56244 219590 56256
rect 268470 56244 268476 56256
rect 268528 56244 268534 56296
rect 379330 56244 379336 56296
rect 379388 56284 379394 56296
rect 427630 56284 427636 56296
rect 379388 56256 427636 56284
rect 379388 56244 379394 56256
rect 427630 56244 427636 56256
rect 427688 56244 427694 56296
rect 57054 56176 57060 56228
rect 57112 56216 57118 56228
rect 92106 56216 92112 56228
rect 57112 56188 92112 56216
rect 57112 56176 57118 56188
rect 92106 56176 92112 56188
rect 92164 56176 92170 56228
rect 218238 56176 218244 56228
rect 218296 56216 218302 56228
rect 266354 56216 266360 56228
rect 218296 56188 266360 56216
rect 218296 56176 218302 56188
rect 266354 56176 266360 56188
rect 266412 56176 266418 56228
rect 379790 56176 379796 56228
rect 379848 56216 379854 56228
rect 426434 56216 426440 56228
rect 379848 56188 426440 56216
rect 379848 56176 379854 56188
rect 426434 56176 426440 56188
rect 426492 56176 426498 56228
rect 56134 56108 56140 56160
rect 56192 56148 56198 56160
rect 88702 56148 88708 56160
rect 56192 56120 88708 56148
rect 56192 56108 56198 56120
rect 88702 56108 88708 56120
rect 88760 56108 88766 56160
rect 219066 56108 219072 56160
rect 219124 56148 219130 56160
rect 253382 56148 253388 56160
rect 219124 56120 253388 56148
rect 219124 56108 219130 56120
rect 253382 56108 253388 56120
rect 253440 56108 253446 56160
rect 379974 56108 379980 56160
rect 380032 56148 380038 56160
rect 414566 56148 414572 56160
rect 380032 56120 414572 56148
rect 380032 56108 380038 56120
rect 414566 56108 414572 56120
rect 414624 56108 414630 56160
rect 54846 56040 54852 56092
rect 54904 56080 54910 56092
rect 86494 56080 86500 56092
rect 54904 56052 86500 56080
rect 54904 56040 54910 56052
rect 86494 56040 86500 56052
rect 86552 56040 86558 56092
rect 218882 56040 218888 56092
rect 218940 56080 218946 56092
rect 251174 56080 251180 56092
rect 218940 56052 251180 56080
rect 218940 56040 218946 56052
rect 251174 56040 251180 56052
rect 251232 56040 251238 56092
rect 379422 56040 379428 56092
rect 379480 56080 379486 56092
rect 412634 56080 412640 56092
rect 379480 56052 412640 56080
rect 379480 56040 379486 56052
rect 412634 56040 412640 56052
rect 412692 56040 412698 56092
rect 53282 55972 53288 56024
rect 53340 56012 53346 56024
rect 81802 56012 81808 56024
rect 53340 55984 81808 56012
rect 53340 55972 53346 55984
rect 81802 55972 81808 55984
rect 81860 55972 81866 56024
rect 219158 55972 219164 56024
rect 219216 56012 219222 56024
rect 248598 56012 248604 56024
rect 219216 55984 248604 56012
rect 219216 55972 219222 55984
rect 248598 55972 248604 55984
rect 248656 55972 248662 56024
rect 376202 55972 376208 56024
rect 376260 56012 376266 56024
rect 408678 56012 408684 56024
rect 376260 55984 408684 56012
rect 376260 55972 376266 55984
rect 408678 55972 408684 55984
rect 408736 55972 408742 56024
rect 52086 55904 52092 55956
rect 52144 55944 52150 55956
rect 79502 55944 79508 55956
rect 52144 55916 79508 55944
rect 52144 55904 52150 55916
rect 79502 55904 79508 55916
rect 79560 55904 79566 55956
rect 215846 55904 215852 55956
rect 215904 55944 215910 55956
rect 245286 55944 245292 55956
rect 215904 55916 245292 55944
rect 215904 55904 215910 55916
rect 245286 55904 245292 55916
rect 245344 55904 245350 55956
rect 379238 55904 379244 55956
rect 379296 55944 379302 55956
rect 411254 55944 411260 55956
rect 379296 55916 411260 55944
rect 379296 55904 379302 55916
rect 411254 55904 411260 55916
rect 411312 55904 411318 55956
rect 49602 55836 49608 55888
rect 49660 55876 49666 55888
rect 157426 55876 157432 55888
rect 49660 55848 157432 55876
rect 49660 55836 49666 55848
rect 157426 55836 157432 55848
rect 157484 55836 157490 55888
rect 213454 55836 213460 55888
rect 213512 55876 213518 55888
rect 275462 55876 275468 55888
rect 213512 55848 275468 55876
rect 213512 55836 213518 55848
rect 275462 55836 275468 55848
rect 275520 55836 275526 55888
rect 371970 55836 371976 55888
rect 372028 55876 372034 55888
rect 399478 55876 399484 55888
rect 372028 55848 399484 55876
rect 372028 55836 372034 55848
rect 399478 55836 399484 55848
rect 399536 55836 399542 55888
rect 219986 55768 219992 55820
rect 220044 55808 220050 55820
rect 408310 55808 408316 55820
rect 220044 55780 408316 55808
rect 220044 55768 220050 55780
rect 408310 55768 408316 55780
rect 408368 55768 408374 55820
rect 213178 55700 213184 55752
rect 213236 55740 213242 55752
rect 273254 55740 273260 55752
rect 213236 55712 273260 55740
rect 213236 55700 213242 55712
rect 273254 55700 273260 55712
rect 273312 55700 273318 55752
rect 55766 55156 55772 55208
rect 55824 55196 55830 55208
rect 117314 55196 117320 55208
rect 55824 55168 117320 55196
rect 55824 55156 55830 55168
rect 117314 55156 117320 55168
rect 117372 55156 117378 55208
rect 216214 55156 216220 55208
rect 216272 55196 216278 55208
rect 242894 55196 242900 55208
rect 216272 55168 242900 55196
rect 216272 55156 216278 55168
rect 242894 55156 242900 55168
rect 242952 55156 242958 55208
rect 375742 55156 375748 55208
rect 375800 55196 375806 55208
rect 436094 55196 436100 55208
rect 375800 55168 436100 55196
rect 375800 55156 375806 55168
rect 436094 55156 436100 55168
rect 436152 55156 436158 55208
rect 52270 55088 52276 55140
rect 52328 55128 52334 55140
rect 113266 55128 113272 55140
rect 52328 55100 113272 55128
rect 52328 55088 52334 55100
rect 113266 55088 113272 55100
rect 113324 55088 113330 55140
rect 215938 55088 215944 55140
rect 215996 55128 216002 55140
rect 271874 55128 271880 55140
rect 215996 55100 271880 55128
rect 215996 55088 216002 55100
rect 271874 55088 271880 55100
rect 271932 55088 271938 55140
rect 375098 55088 375104 55140
rect 375156 55128 375162 55140
rect 397454 55128 397460 55140
rect 375156 55100 397460 55128
rect 375156 55088 375162 55100
rect 397454 55088 397460 55100
rect 397512 55088 397518 55140
rect 55674 55020 55680 55072
rect 55732 55060 55738 55072
rect 114554 55060 114560 55072
rect 55732 55032 114560 55060
rect 55732 55020 55738 55032
rect 114554 55020 114560 55032
rect 114612 55020 114618 55072
rect 216122 55020 216128 55072
rect 216180 55060 216186 55072
rect 269114 55060 269120 55072
rect 216180 55032 269120 55060
rect 216180 55020 216186 55032
rect 269114 55020 269120 55032
rect 269172 55020 269178 55072
rect 374178 55020 374184 55072
rect 374236 55060 374242 55072
rect 431954 55060 431960 55072
rect 374236 55032 431960 55060
rect 374236 55020 374242 55032
rect 431954 55020 431960 55032
rect 432012 55020 432018 55072
rect 52178 54952 52184 55004
rect 52236 54992 52242 55004
rect 109034 54992 109040 55004
rect 52236 54964 109040 54992
rect 52236 54952 52242 54964
rect 109034 54952 109040 54964
rect 109092 54952 109098 55004
rect 219710 54952 219716 55004
rect 219768 54992 219774 55004
rect 266446 54992 266452 55004
rect 219768 54964 266452 54992
rect 219768 54952 219774 54964
rect 266446 54952 266452 54964
rect 266504 54952 266510 55004
rect 374730 54952 374736 55004
rect 374788 54992 374794 55004
rect 430574 54992 430580 55004
rect 374788 54964 430580 54992
rect 374788 54952 374794 54964
rect 430574 54952 430580 54964
rect 430632 54952 430638 55004
rect 53098 54884 53104 54936
rect 53156 54924 53162 54936
rect 86954 54924 86960 54936
rect 53156 54896 86960 54924
rect 53156 54884 53162 54896
rect 86954 54884 86960 54896
rect 87012 54884 87018 54936
rect 219618 54884 219624 54936
rect 219676 54924 219682 54936
rect 264974 54924 264980 54936
rect 219676 54896 264980 54924
rect 219676 54884 219682 54896
rect 264974 54884 264980 54896
rect 265032 54884 265038 54936
rect 374914 54884 374920 54936
rect 374972 54924 374978 54936
rect 429194 54924 429200 54936
rect 374972 54896 429200 54924
rect 374972 54884 374978 54896
rect 429194 54884 429200 54896
rect 429252 54884 429258 54936
rect 58618 54816 58624 54868
rect 58676 54856 58682 54868
rect 92474 54856 92480 54868
rect 58676 54828 92480 54856
rect 58676 54816 58682 54828
rect 92474 54816 92480 54828
rect 92532 54816 92538 54868
rect 219802 54816 219808 54868
rect 219860 54856 219866 54868
rect 253934 54856 253940 54868
rect 219860 54828 253940 54856
rect 219860 54816 219866 54828
rect 253934 54816 253940 54828
rect 253992 54816 253998 54868
rect 377950 54816 377956 54868
rect 378008 54856 378014 54868
rect 411346 54856 411352 54868
rect 378008 54828 411352 54856
rect 378008 54816 378014 54828
rect 411346 54816 411352 54828
rect 411404 54816 411410 54868
rect 56226 54748 56232 54800
rect 56284 54788 56290 54800
rect 89714 54788 89720 54800
rect 56284 54760 89720 54788
rect 56284 54748 56290 54760
rect 89714 54748 89720 54760
rect 89772 54748 89778 54800
rect 217134 54748 217140 54800
rect 217192 54788 217198 54800
rect 251358 54788 251364 54800
rect 217192 54760 251364 54788
rect 217192 54748 217198 54760
rect 251358 54748 251364 54760
rect 251416 54748 251422 54800
rect 378042 54748 378048 54800
rect 378100 54788 378106 54800
rect 409874 54788 409880 54800
rect 378100 54760 409880 54788
rect 378100 54748 378106 54760
rect 409874 54748 409880 54760
rect 409932 54748 409938 54800
rect 58986 54680 58992 54732
rect 59044 54720 59050 54732
rect 91186 54720 91192 54732
rect 59044 54692 91192 54720
rect 59044 54680 59050 54692
rect 91186 54680 91192 54692
rect 91244 54680 91250 54732
rect 217042 54680 217048 54732
rect 217100 54720 217106 54732
rect 249794 54720 249800 54732
rect 217100 54692 249800 54720
rect 217100 54680 217106 54692
rect 249794 54680 249800 54692
rect 249852 54680 249858 54732
rect 376478 54680 376484 54732
rect 376536 54720 376542 54732
rect 405826 54720 405832 54732
rect 376536 54692 405832 54720
rect 376536 54680 376542 54692
rect 405826 54680 405832 54692
rect 405884 54680 405890 54732
rect 53374 54612 53380 54664
rect 53432 54652 53438 54664
rect 80054 54652 80060 54664
rect 53432 54624 80060 54652
rect 53432 54612 53438 54624
rect 80054 54612 80060 54624
rect 80112 54612 80118 54664
rect 216030 54612 216036 54664
rect 216088 54652 216094 54664
rect 247034 54652 247040 54664
rect 216088 54624 247040 54652
rect 216088 54612 216094 54624
rect 247034 54612 247040 54624
rect 247092 54612 247098 54664
rect 375282 54612 375288 54664
rect 375340 54652 375346 54664
rect 404354 54652 404360 54664
rect 375340 54624 404360 54652
rect 375340 54612 375346 54624
rect 404354 54612 404360 54624
rect 404412 54612 404418 54664
rect 214650 54544 214656 54596
rect 214708 54584 214714 54596
rect 245654 54584 245660 54596
rect 214708 54556 245660 54584
rect 214708 54544 214714 54556
rect 245654 54544 245660 54556
rect 245712 54544 245718 54596
rect 378778 54544 378784 54596
rect 378836 54584 378842 54596
rect 407206 54584 407212 54596
rect 378836 54556 407212 54584
rect 378836 54544 378842 54556
rect 407206 54544 407212 54556
rect 407264 54544 407270 54596
rect 215110 54476 215116 54528
rect 215168 54516 215174 54528
rect 244366 54516 244372 54528
rect 215168 54488 244372 54516
rect 215168 54476 215174 54488
rect 244366 54476 244372 54488
rect 244424 54476 244430 54528
rect 373718 54476 373724 54528
rect 373776 54516 373782 54528
rect 400214 54516 400220 54528
rect 373776 54488 400220 54516
rect 373776 54476 373782 54488
rect 400214 54476 400220 54488
rect 400272 54476 400278 54528
rect 213270 54408 213276 54460
rect 213328 54448 213334 54460
rect 273346 54448 273352 54460
rect 213328 54420 273352 54448
rect 213328 54408 213334 54420
rect 273346 54408 273352 54420
rect 273404 54408 273410 54460
rect 373626 54408 373632 54460
rect 373684 54448 373690 54460
rect 433426 54448 433432 54460
rect 373684 54420 433432 54448
rect 373684 54408 373690 54420
rect 433426 54408 433432 54420
rect 433484 54408 433490 54460
rect 213362 54340 213368 54392
rect 213420 54380 213426 54392
rect 240134 54380 240140 54392
rect 213420 54352 240140 54380
rect 213420 54340 213426 54352
rect 240134 54340 240140 54352
rect 240192 54340 240198 54392
rect 214558 54272 214564 54324
rect 214616 54312 214622 54324
rect 237374 54312 237380 54324
rect 214616 54284 237380 54312
rect 214616 54272 214622 54284
rect 237374 54272 237380 54284
rect 237432 54272 237438 54324
rect 2774 20340 2780 20392
rect 2832 20380 2838 20392
rect 4798 20380 4804 20392
rect 2832 20352 4804 20380
rect 2832 20340 2838 20352
rect 4798 20340 4804 20352
rect 4856 20340 4862 20392
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 57238 3448 57244 3460
rect 624 3420 57244 3448
rect 624 3408 630 3420
rect 57238 3408 57244 3420
rect 57296 3408 57302 3460
rect 125870 3408 125876 3460
rect 125928 3448 125934 3460
rect 366358 3448 366364 3460
rect 125928 3420 366364 3448
rect 125928 3408 125934 3420
rect 366358 3408 366364 3420
rect 366416 3408 366422 3460
<< via1 >>
rect 235172 700340 235224 700392
rect 305644 700340 305696 700392
rect 57888 700272 57940 700324
rect 543464 700272 543516 700324
rect 137836 683136 137888 683188
rect 580172 683136 580224 683188
rect 299480 640976 299532 641028
rect 400680 640976 400732 641028
rect 3424 639548 3476 639600
rect 317052 639548 317104 639600
rect 104900 636828 104952 636880
rect 429384 636828 429436 636880
rect 169760 635468 169812 635520
rect 430948 635468 431000 635520
rect 316868 634856 316920 634908
rect 430580 634856 430632 634908
rect 316960 634788 317012 634840
rect 430856 634788 430908 634840
rect 318800 634040 318852 634092
rect 494060 634040 494112 634092
rect 298100 633632 298152 633684
rect 435364 633632 435416 633684
rect 289820 633564 289872 633616
rect 432604 633564 432656 633616
rect 296720 633496 296772 633548
rect 494336 633496 494388 633548
rect 288440 633428 288492 633480
rect 510712 633428 510764 633480
rect 316684 632952 316736 633004
rect 396632 632952 396684 633004
rect 300124 632884 300176 632936
rect 378600 632884 378652 632936
rect 318248 632816 318300 632868
rect 428188 632816 428240 632868
rect 312544 632748 312596 632800
rect 337384 632748 337436 632800
rect 319444 632680 319496 632732
rect 355416 632680 355468 632732
rect 364340 632680 364392 632732
rect 423680 632680 423732 632732
rect 318156 632612 318208 632664
rect 359924 632612 359976 632664
rect 307024 632544 307076 632596
rect 350908 632544 350960 632596
rect 313924 632476 313976 632528
rect 364432 632476 364484 632528
rect 319720 632408 319772 632460
rect 373448 632408 373500 632460
rect 316776 632340 316828 632392
rect 383108 632340 383160 632392
rect 314016 632272 314068 632324
rect 387616 632272 387668 632324
rect 315304 632204 315356 632256
rect 332876 632204 332928 632256
rect 320364 632136 320416 632188
rect 341892 632136 341944 632188
rect 319628 632068 319680 632120
rect 323860 632068 323912 632120
rect 414664 632068 414716 632120
rect 457444 632068 457496 632120
rect 284944 631320 284996 631372
rect 368940 631320 368992 631372
rect 285036 631252 285088 631304
rect 419172 631252 419224 631304
rect 298192 631184 298244 631236
rect 432696 631184 432748 631236
rect 319812 631116 319864 631168
rect 457536 631116 457588 631168
rect 291200 631048 291252 631100
rect 429844 631048 429896 631100
rect 318064 630980 318116 631032
rect 471152 630980 471204 631032
rect 293960 630912 294012 630964
rect 510620 630912 510672 630964
rect 287060 630844 287112 630896
rect 512000 630844 512052 630896
rect 319076 630776 319128 630828
rect 580172 630776 580224 630828
rect 18604 630708 18656 630760
rect 409880 630708 409932 630760
rect 218704 630640 218756 630692
rect 414572 630640 414624 630692
rect 280712 629960 280764 630012
rect 320364 630436 320416 630488
rect 217784 629892 217836 629944
rect 319076 629892 319128 629944
rect 309784 629280 309836 629332
rect 317788 629280 317840 629332
rect 100576 625744 100628 625796
rect 124680 625744 124732 625796
rect 213920 625744 213972 625796
rect 225420 625744 225472 625796
rect 115388 625676 115440 625728
rect 124588 625676 124640 625728
rect 137744 625676 137796 625728
rect 186504 625676 186556 625728
rect 206468 625676 206520 625728
rect 231308 625676 231360 625728
rect 112168 625608 112220 625660
rect 124496 625608 124548 625660
rect 139308 625608 139360 625660
rect 162860 625608 162912 625660
rect 212540 625608 212592 625660
rect 271880 625608 271932 625660
rect 83188 625540 83240 625592
rect 125692 625540 125744 625592
rect 135168 625540 135220 625592
rect 160284 625540 160336 625592
rect 217876 625540 217928 625592
rect 242900 625540 242952 625592
rect 109592 625472 109644 625524
rect 122840 625472 122892 625524
rect 136364 625472 136416 625524
rect 166172 625472 166224 625524
rect 218888 625472 218940 625524
rect 251916 625472 251968 625524
rect 106372 625404 106424 625456
rect 120908 625404 120960 625456
rect 139124 625404 139176 625456
rect 174452 625404 174504 625456
rect 218796 625404 218848 625456
rect 263600 625404 263652 625456
rect 103796 625336 103848 625388
rect 122288 625336 122340 625388
rect 134892 625336 134944 625388
rect 180340 625336 180392 625388
rect 190000 625336 190052 625388
rect 204444 625336 204496 625388
rect 209780 625336 209832 625388
rect 260196 625336 260248 625388
rect 54852 625268 54904 625320
rect 88984 625268 89036 625320
rect 124220 625268 124272 625320
rect 171876 625268 171928 625320
rect 214012 625268 214064 625320
rect 269212 625268 269264 625320
rect 55128 625200 55180 625252
rect 92204 625200 92256 625252
rect 94780 625200 94832 625252
rect 121644 625200 121696 625252
rect 135260 625200 135312 625252
rect 183652 625200 183704 625252
rect 192576 625200 192628 625252
rect 201684 625200 201736 625252
rect 219348 625200 219400 625252
rect 275100 625200 275152 625252
rect 56508 625132 56560 625184
rect 77392 625132 77444 625184
rect 133880 625132 133932 625184
rect 139860 625132 139912 625184
rect 157524 625132 157576 625184
rect 195704 625132 195756 625184
rect 200856 625132 200908 625184
rect 289084 625132 289136 625184
rect 317604 625132 317656 625184
rect 140136 625064 140188 625116
rect 215300 624044 215352 624096
rect 234620 624044 234672 624096
rect 219624 623976 219676 624028
rect 246028 623976 246080 624028
rect 59360 623908 59412 623960
rect 98000 623908 98052 623960
rect 210424 623908 210476 623960
rect 237564 623908 237616 623960
rect 57796 623840 57848 623892
rect 80612 623840 80664 623892
rect 86408 623840 86460 623892
rect 124312 623840 124364 623892
rect 133144 623840 133196 623892
rect 151268 623840 151320 623892
rect 206284 623840 206336 623892
rect 254492 623840 254544 623892
rect 69020 623772 69072 623824
rect 124404 623772 124456 623824
rect 136640 623772 136692 623824
rect 168748 623772 168800 623824
rect 204260 623772 204312 623824
rect 277676 623772 277728 623824
rect 217968 622820 218020 622872
rect 228732 622820 228784 622872
rect 135076 622752 135128 622804
rect 145564 622752 145616 622804
rect 214564 622752 214616 622804
rect 257620 622752 257672 622804
rect 126244 622684 126296 622736
rect 177856 622684 177908 622736
rect 204352 622684 204404 622736
rect 222844 622684 222896 622736
rect 55036 622616 55088 622668
rect 62948 622616 63000 622668
rect 136456 622616 136508 622668
rect 149152 622616 149204 622668
rect 208400 622616 208452 622668
rect 240324 622616 240376 622668
rect 54944 622548 54996 622600
rect 65524 622548 65576 622600
rect 136548 622548 136600 622600
rect 154580 622548 154632 622600
rect 206376 622548 206428 622600
rect 248696 622548 248748 622600
rect 56324 622480 56376 622532
rect 71228 622480 71280 622532
rect 134984 622480 135036 622532
rect 142988 622480 143040 622532
rect 211804 622480 211856 622532
rect 266268 622480 266320 622532
rect 280712 622480 280764 622532
rect 56416 622412 56468 622464
rect 74632 622412 74684 622464
rect 137928 622412 137980 622464
rect 218704 622412 218756 622464
rect 118240 622344 118292 622396
rect 121552 622344 121604 622396
rect 198280 622344 198332 622396
rect 202236 622344 202288 622396
rect 217324 622344 217376 622396
rect 219716 622344 219768 622396
rect 280712 622276 280764 622328
rect 432604 621732 432656 621784
rect 483204 621732 483256 621784
rect 432696 621664 432748 621716
rect 501236 621664 501288 621716
rect 465172 620984 465224 621036
rect 515404 620984 515456 621036
rect 429844 620916 429896 620968
rect 456800 620916 456852 620968
rect 213184 619624 213236 619676
rect 216680 619624 216732 619676
rect 311164 619624 311216 619676
rect 317972 619624 318024 619676
rect 208492 616836 208544 616888
rect 216680 616836 216732 616888
rect 286324 615476 286376 615528
rect 317972 615476 318024 615528
rect 287704 609968 287756 610020
rect 317880 609968 317932 610020
rect 435364 608540 435416 608592
rect 456800 608540 456852 608592
rect 132500 607180 132552 607232
rect 136732 607180 136784 607232
rect 204904 607180 204956 607232
rect 216680 607180 216732 607232
rect 304264 605820 304316 605872
rect 317972 605820 318024 605872
rect 294604 600312 294656 600364
rect 317604 600312 317656 600364
rect 200948 598000 201000 598052
rect 203064 598000 203116 598052
rect 287796 596164 287848 596216
rect 317604 596164 317656 596216
rect 207020 593376 207072 593428
rect 216680 593376 216732 593428
rect 302240 589908 302292 589960
rect 319812 589908 319864 589960
rect 124128 589364 124180 589416
rect 134616 589364 134668 589416
rect 134524 589296 134576 589348
rect 136732 589296 136784 589348
rect 203248 589296 203300 589348
rect 204536 589296 204588 589348
rect 210516 589296 210568 589348
rect 216680 589296 216732 589348
rect 283656 589296 283708 589348
rect 302240 589296 302292 589348
rect 211160 586848 211212 586900
rect 216680 586848 216732 586900
rect 293224 586508 293276 586560
rect 317420 586508 317472 586560
rect 515404 585760 515456 585812
rect 580172 585760 580224 585812
rect 57520 583720 57572 583772
rect 58624 583720 58676 583772
rect 304356 582360 304408 582412
rect 317972 582360 318024 582412
rect 217692 581680 217744 581732
rect 218704 581680 218756 581732
rect 125600 576852 125652 576904
rect 136732 576852 136784 576904
rect 300216 576852 300268 576904
rect 317880 576852 317932 576904
rect 206560 574064 206612 574116
rect 216680 574064 216732 574116
rect 513288 572704 513340 572756
rect 560944 572704 560996 572756
rect 57336 572296 57388 572348
rect 58716 572296 58768 572348
rect 210608 571344 210660 571396
rect 216680 571344 216732 571396
rect 289176 571344 289228 571396
rect 317972 571344 318024 571396
rect 209044 562300 209096 562352
rect 217416 562300 217468 562352
rect 57888 561144 57940 561196
rect 137284 561144 137336 561196
rect 3424 561076 3476 561128
rect 304356 561076 304408 561128
rect 201040 560464 201092 560516
rect 202880 560464 202932 560516
rect 217692 560260 217744 560312
rect 220176 560260 220228 560312
rect 57152 560192 57204 560244
rect 62120 560192 62172 560244
rect 137652 560192 137704 560244
rect 140780 560192 140832 560244
rect 106280 560124 106332 560176
rect 124588 560124 124640 560176
rect 134616 560124 134668 560176
rect 204536 560192 204588 560244
rect 302240 560192 302292 560244
rect 98092 560056 98144 560108
rect 122840 560056 122892 560108
rect 96804 559988 96856 560040
rect 124496 559988 124548 560040
rect 164332 559988 164384 560040
rect 200856 559988 200908 560040
rect 93860 559920 93912 559972
rect 124680 559920 124732 559972
rect 182364 559920 182416 559972
rect 218888 559920 218940 559972
rect 260840 559920 260892 559972
rect 316960 559920 317012 559972
rect 57060 559852 57112 559904
rect 67732 559852 67784 559904
rect 86960 559852 87012 559904
rect 120908 559852 120960 559904
rect 137744 559852 137796 559904
rect 145104 559852 145156 559904
rect 157984 559852 158036 559904
rect 203340 559852 203392 559904
rect 258080 559852 258132 559904
rect 316868 559852 316920 559904
rect 59084 559784 59136 559836
rect 82912 559784 82964 559836
rect 87052 559784 87104 559836
rect 121552 559784 121604 559836
rect 139032 559784 139084 559836
rect 150624 559784 150676 559836
rect 154580 559784 154632 559836
rect 201684 559784 201736 559836
rect 216128 559784 216180 559836
rect 282920 559784 282972 559836
rect 54852 559716 54904 559768
rect 78680 559716 78732 559768
rect 85580 559716 85632 559768
rect 121736 559716 121788 559768
rect 134892 559716 134944 559768
rect 151820 559716 151872 559768
rect 156052 559716 156104 559768
rect 204444 559716 204496 559768
rect 247040 559716 247092 559768
rect 319720 559716 319772 559768
rect 67640 559648 67692 559700
rect 121920 559648 121972 559700
rect 136364 559648 136416 559700
rect 161664 559648 161716 559700
rect 179696 559648 179748 559700
rect 281540 559648 281592 559700
rect 63500 559580 63552 559632
rect 122932 559580 122984 559632
rect 138848 559580 138900 559632
rect 165620 559580 165672 559632
rect 180800 559580 180852 559632
rect 283196 559580 283248 559632
rect 3424 559512 3476 559564
rect 286324 559512 286376 559564
rect 217876 559308 217928 559360
rect 222200 559308 222252 559360
rect 219348 559036 219400 559088
rect 223580 559036 223632 559088
rect 139124 558900 139176 558952
rect 142160 558900 142212 558952
rect 57428 558832 57480 558884
rect 60740 558832 60792 558884
rect 100760 558764 100812 558816
rect 102876 558764 102928 558816
rect 116584 558764 116636 558816
rect 120172 558764 120224 558816
rect 161572 558764 161624 558816
rect 168472 558764 168524 558816
rect 173900 558764 173952 558816
rect 179604 558764 179656 558816
rect 225144 558764 225196 558816
rect 227996 558764 228048 558816
rect 260104 558764 260156 558816
rect 262772 558764 262824 558816
rect 278044 558764 278096 558816
rect 280252 558764 280304 558816
rect 60280 558696 60332 558748
rect 62764 558696 62816 558748
rect 119344 558696 119396 558748
rect 120724 558696 120776 558748
rect 147680 558628 147732 558680
rect 162308 558628 162360 558680
rect 151360 558560 151412 558612
rect 164884 558560 164936 558612
rect 231952 558560 232004 558612
rect 259644 558560 259696 558612
rect 142896 558492 142948 558544
rect 160744 558492 160796 558544
rect 222292 558492 222344 558544
rect 253940 558492 253992 558544
rect 68744 558424 68796 558476
rect 71044 558424 71096 558476
rect 82728 558424 82780 558476
rect 88984 558424 89036 558476
rect 140320 558424 140372 558476
rect 159364 558424 159416 558476
rect 188344 558424 188396 558476
rect 200212 558424 200264 558476
rect 212632 558424 212684 558476
rect 251180 558424 251232 558476
rect 77024 558356 77076 558408
rect 85672 558356 85724 558408
rect 94504 558356 94556 558408
rect 104164 558356 104216 558408
rect 112444 558356 112496 558408
rect 117412 558356 117464 558408
rect 129740 558356 129792 558408
rect 153844 558356 153896 558408
rect 154672 558356 154724 558408
rect 171324 558356 171376 558408
rect 187884 558356 187936 558408
rect 233884 558356 233936 558408
rect 62856 558288 62908 558340
rect 80704 558288 80756 558340
rect 86040 558288 86092 558340
rect 108304 558288 108356 558340
rect 111892 558288 111944 558340
rect 123116 558288 123168 558340
rect 133972 558288 134024 558340
rect 197452 558288 197504 558340
rect 227720 558288 227772 558340
rect 245660 558288 245712 558340
rect 249800 558288 249852 558340
rect 294604 558288 294656 558340
rect 71320 558220 71372 558272
rect 93952 558220 94004 558272
rect 100208 558220 100260 558272
rect 115204 558220 115256 558272
rect 118700 558220 118752 558272
rect 144920 558220 144972 558272
rect 158720 558220 158772 558272
rect 182916 558220 182968 558272
rect 190460 558220 190512 558272
rect 257068 558220 257120 558272
rect 273260 558220 273312 558272
rect 318248 558220 318300 558272
rect 58900 558152 58952 558204
rect 74540 558152 74592 558204
rect 79876 558152 79928 558204
rect 114560 558152 114612 558204
rect 132592 558152 132644 558204
rect 177028 558152 177080 558204
rect 177304 558152 177356 558204
rect 188620 558152 188672 558204
rect 191840 558152 191892 558204
rect 276940 558152 276992 558204
rect 71780 557880 71832 557932
rect 73804 557880 73856 557932
rect 184204 557880 184256 557932
rect 185492 557880 185544 557932
rect 264244 557880 264296 557932
rect 265348 557880 265400 557932
rect 262864 557608 262916 557660
rect 268660 557608 268712 557660
rect 64144 557540 64196 557592
rect 65064 557540 65116 557592
rect 222936 557540 222988 557592
rect 224408 557540 224460 557592
rect 267740 557540 267792 557592
rect 317420 557540 317472 557592
rect 219256 557472 219308 557524
rect 223672 557472 223724 557524
rect 178040 557064 178092 557116
rect 206560 557064 206612 557116
rect 269488 557064 269540 557116
rect 300216 557064 300268 557116
rect 57336 556996 57388 557048
rect 81716 556996 81768 557048
rect 122840 556996 122892 557048
rect 202144 556996 202196 557048
rect 229284 556996 229336 557048
rect 281264 556996 281316 557048
rect 78864 556928 78916 556980
rect 121460 556928 121512 556980
rect 143540 556928 143592 556980
rect 156420 556928 156472 556980
rect 159824 556928 159876 556980
rect 173440 556928 173492 556980
rect 194600 556928 194652 556980
rect 283656 556928 283708 556980
rect 63776 556860 63828 556912
rect 123576 556860 123628 556912
rect 138940 556860 138992 556912
rect 160100 556860 160152 556912
rect 179512 556860 179564 556912
rect 281908 556860 281960 556912
rect 4804 556792 4856 556844
rect 318340 556792 318392 556844
rect 219532 556724 219584 556776
rect 219900 556724 219952 556776
rect 193220 555704 193272 555756
rect 218796 555704 218848 555756
rect 266544 555704 266596 555756
rect 307024 555704 307076 555756
rect 168380 555636 168432 555688
rect 200672 555636 200724 555688
rect 240784 555636 240836 555688
rect 283472 555636 283524 555688
rect 59268 555568 59320 555620
rect 92572 555568 92624 555620
rect 100392 555568 100444 555620
rect 123484 555568 123536 555620
rect 137836 555568 137888 555620
rect 149060 555568 149112 555620
rect 157892 555568 157944 555620
rect 203248 555568 203300 555620
rect 245108 555568 245160 555620
rect 318156 555568 318208 555620
rect 64880 555500 64932 555552
rect 122196 555500 122248 555552
rect 138572 555500 138624 555552
rect 169116 555500 169168 555552
rect 181352 555500 181404 555552
rect 281724 555500 281776 555552
rect 3516 555432 3568 555484
rect 319720 555432 319772 555484
rect 129832 554208 129884 554260
rect 202972 554208 203024 554260
rect 246488 554208 246540 554260
rect 287704 554208 287756 554260
rect 73252 554140 73304 554192
rect 108580 554140 108632 554192
rect 122932 554140 122984 554192
rect 201868 554140 201920 554192
rect 263692 554140 263744 554192
rect 315304 554140 315356 554192
rect 58532 554072 58584 554124
rect 110420 554072 110472 554124
rect 195980 554072 196032 554124
rect 283380 554072 283432 554124
rect 66720 554004 66772 554056
rect 121184 554004 121236 554056
rect 182272 554004 182324 554056
rect 282000 554004 282052 554056
rect 3516 553392 3568 553444
rect 317972 553392 318024 553444
rect 226432 552916 226484 552968
rect 280804 552916 280856 552968
rect 59452 552848 59504 552900
rect 75920 552848 75972 552900
rect 88616 552848 88668 552900
rect 103520 552848 103572 552900
rect 106924 552848 106976 552900
rect 123392 552848 123444 552900
rect 129004 552848 129056 552900
rect 203156 552848 203208 552900
rect 256700 552848 256752 552900
rect 316776 552848 316828 552900
rect 75276 552780 75328 552832
rect 96988 552780 97040 552832
rect 121460 552780 121512 552832
rect 201132 552780 201184 552832
rect 250812 552780 250864 552832
rect 319628 552780 319680 552832
rect 57704 552712 57756 552764
rect 77392 552712 77444 552764
rect 80060 552712 80112 552764
rect 120816 552712 120868 552764
rect 138480 552712 138532 552764
rect 160652 552712 160704 552764
rect 196348 552712 196400 552764
rect 283288 552712 283340 552764
rect 69020 552644 69072 552696
rect 114652 552644 114704 552696
rect 138664 552644 138716 552696
rect 174912 552644 174964 552696
rect 179144 552644 179196 552696
rect 271236 552644 271288 552696
rect 192116 551624 192168 551676
rect 217324 551624 217376 551676
rect 281540 551624 281592 551676
rect 293224 551624 293276 551676
rect 176660 551556 176712 551608
rect 210516 551556 210568 551608
rect 260012 551556 260064 551608
rect 289176 551556 289228 551608
rect 80980 551488 81032 551540
rect 122104 551488 122156 551540
rect 144092 551488 144144 551540
rect 201776 551488 201828 551540
rect 253664 551488 253716 551540
rect 316684 551488 316736 551540
rect 57520 551420 57572 551472
rect 89812 551420 89864 551472
rect 93952 551420 94004 551472
rect 114652 551420 114704 551472
rect 121552 551420 121604 551472
rect 201592 551420 201644 551472
rect 211620 551420 211672 551472
rect 280988 551420 281040 551472
rect 282920 551420 282972 551472
rect 304264 551420 304316 551472
rect 58992 551352 59044 551404
rect 102508 551352 102560 551404
rect 200672 551352 200724 551404
rect 281816 551352 281868 551404
rect 65984 551284 66036 551336
rect 123208 551284 123260 551336
rect 139400 551284 139452 551336
rect 159088 551284 159140 551336
rect 186320 551284 186372 551336
rect 283564 551284 283616 551336
rect 176752 550128 176804 550180
rect 225052 550128 225104 550180
rect 228640 550128 228692 550180
rect 280896 550128 280948 550180
rect 80704 550060 80756 550112
rect 109684 550060 109736 550112
rect 142620 550060 142672 550112
rect 202328 550060 202380 550112
rect 251548 550060 251600 550112
rect 313924 550060 313976 550112
rect 59544 549992 59596 550044
rect 101036 549992 101088 550044
rect 120264 549992 120316 550044
rect 190552 549992 190604 550044
rect 193496 549992 193548 550044
rect 213184 549992 213236 550044
rect 242900 549992 242952 550044
rect 314016 549992 314068 550044
rect 69112 549924 69164 549976
rect 121000 549924 121052 549976
rect 138756 549924 138808 549976
rect 153384 549924 153436 549976
rect 189080 549924 189132 549976
rect 262864 549924 262916 549976
rect 271604 549924 271656 549976
rect 289084 549924 289136 549976
rect 70952 549856 71004 549908
rect 121828 549856 121880 549908
rect 147772 549856 147824 549908
rect 167092 549856 167144 549908
rect 187056 549856 187108 549908
rect 283104 549856 283156 549908
rect 40040 549176 40092 549228
rect 317972 549176 318024 549228
rect 199200 548700 199252 548752
rect 215944 548700 215996 548752
rect 88432 548632 88484 548684
rect 104900 548632 104952 548684
rect 189908 548632 189960 548684
rect 206468 548632 206520 548684
rect 76748 548564 76800 548616
rect 112444 548564 112496 548616
rect 205640 548564 205692 548616
rect 264244 548564 264296 548616
rect 59176 548496 59228 548548
rect 108212 548496 108264 548548
rect 136916 548496 136968 548548
rect 201500 548496 201552 548548
rect 210148 548496 210200 548548
rect 281172 548496 281224 548548
rect 57612 547340 57664 547392
rect 91744 547340 91796 547392
rect 140504 547340 140556 547392
rect 188344 547340 188396 547392
rect 190644 547340 190696 547392
rect 204904 547340 204956 547392
rect 211068 547340 211120 547392
rect 236000 547340 236052 547392
rect 259552 547340 259604 547392
rect 309784 547340 309836 547392
rect 84568 547272 84620 547324
rect 122012 547272 122064 547324
rect 124680 547272 124732 547324
rect 201224 547272 201276 547324
rect 235080 547272 235132 547324
rect 319536 547272 319588 547324
rect 62764 547204 62816 547256
rect 105360 547204 105412 547256
rect 185584 547204 185636 547256
rect 274640 547204 274692 547256
rect 63132 547136 63184 547188
rect 110512 547136 110564 547188
rect 122656 547136 122708 547188
rect 137468 547136 137520 547188
rect 147680 547136 147732 547188
rect 184204 547136 184256 547188
rect 187792 547136 187844 547188
rect 283012 547136 283064 547188
rect 273260 547068 273312 547120
rect 274456 547068 274508 547120
rect 139860 546456 139912 546508
rect 141884 546456 141936 546508
rect 184940 545980 184992 546032
rect 216036 545980 216088 546032
rect 138296 545912 138348 545964
rect 200764 545912 200816 545964
rect 206376 545912 206428 545964
rect 241520 545912 241572 545964
rect 267280 545912 267332 545964
rect 300124 545912 300176 545964
rect 82452 545844 82504 545896
rect 116584 545844 116636 545896
rect 139032 545844 139084 545896
rect 202052 545844 202104 545896
rect 217876 545844 217928 545896
rect 260104 545844 260156 545896
rect 275192 545844 275244 545896
rect 312544 545844 312596 545896
rect 57244 545776 57296 545828
rect 103244 545776 103296 545828
rect 198556 545776 198608 545828
rect 278044 545776 278096 545828
rect 71688 545708 71740 545760
rect 123024 545708 123076 545760
rect 127624 545708 127676 545760
rect 194692 545708 194744 545760
rect 197820 545708 197872 545760
rect 210608 545708 210660 545760
rect 234344 545708 234396 545760
rect 319444 545708 319496 545760
rect 289544 545096 289596 545148
rect 313924 545096 313976 545148
rect 154580 544756 154632 544808
rect 155500 544756 155552 544808
rect 171324 544552 171376 544604
rect 203432 544552 203484 544604
rect 161388 544484 161440 544536
rect 203064 544484 203116 544536
rect 219164 544484 219216 544536
rect 227168 544484 227220 544536
rect 270132 544484 270184 544536
rect 287796 544484 287848 544536
rect 94596 544416 94648 544468
rect 123300 544416 123352 544468
rect 137928 544416 137980 544468
rect 149796 544416 149848 544468
rect 152648 544416 152700 544468
rect 201960 544416 202012 544468
rect 220728 544416 220780 544468
rect 247132 544416 247184 544468
rect 279516 544416 279568 544468
rect 311164 544416 311216 544468
rect 71044 544348 71096 544400
rect 108948 544348 109000 544400
rect 131212 544348 131264 544400
rect 177304 544348 177356 544400
rect 184204 544348 184256 544400
rect 281632 544348 281684 544400
rect 290924 544144 290976 544196
rect 287428 544076 287480 544128
rect 69112 544008 69164 544060
rect 70308 544008 70360 544060
rect 104164 544008 104216 544060
rect 113272 544008 113324 544060
rect 121092 544008 121144 544060
rect 121552 544008 121604 544060
rect 122564 544008 122616 544060
rect 63500 543872 63552 543924
rect 64512 543872 64564 543924
rect 78680 543872 78732 543924
rect 79600 543872 79652 543924
rect 88432 543872 88484 543924
rect 89628 543872 89680 543924
rect 89812 543872 89864 543924
rect 91008 543872 91060 543924
rect 100760 543872 100812 543924
rect 101772 543872 101824 543924
rect 61660 543668 61712 543720
rect 64144 543668 64196 543720
rect 88984 543668 89036 543720
rect 90364 543668 90416 543720
rect 291200 543940 291252 543992
rect 292396 543940 292448 543992
rect 293960 543940 294012 543992
rect 295248 543940 295300 543992
rect 314016 544008 314068 544060
rect 314384 543940 314436 543992
rect 106280 543872 106332 543924
rect 107568 543872 107620 543924
rect 114560 543872 114612 543924
rect 115388 543872 115440 543924
rect 124220 543872 124272 543924
rect 125416 543872 125468 543924
rect 125600 543872 125652 543924
rect 126888 543872 126940 543924
rect 129740 543872 129792 543924
rect 130476 543872 130528 543924
rect 136640 543872 136692 543924
rect 137652 543872 137704 543924
rect 142160 543872 142212 543924
rect 143356 543872 143408 543924
rect 143540 543872 143592 543924
rect 144736 543872 144788 543924
rect 158720 543872 158772 543924
rect 159824 543872 159876 543924
rect 161572 543872 161624 543924
rect 162676 543872 162728 543924
rect 164332 543872 164384 543924
rect 165528 543872 165580 543924
rect 179512 543872 179564 543924
rect 180616 543872 180668 543924
rect 180800 543872 180852 543924
rect 181996 543872 182048 543924
rect 191840 543872 191892 543924
rect 192760 543872 192812 543924
rect 193220 543872 193272 543924
rect 194232 543872 194284 543924
rect 195980 543872 196032 543924
rect 197084 543872 197136 543924
rect 208400 543872 208452 543924
rect 209228 543872 209280 543924
rect 212540 543872 212592 543924
rect 213552 543872 213604 543924
rect 213920 543872 213972 543924
rect 215024 543872 215076 543924
rect 222200 543872 222252 543924
rect 222844 543872 222896 543924
rect 256700 543872 256752 543924
rect 257988 543872 258040 543924
rect 285220 543872 285272 543924
rect 314108 543872 314160 543924
rect 137560 543804 137612 543856
rect 139768 543804 139820 543856
rect 252284 543804 252336 543856
rect 317972 543804 318024 543856
rect 237932 543736 237984 543788
rect 316684 543736 316736 543788
rect 106096 543668 106148 543720
rect 108304 543668 108356 543720
rect 111800 543668 111852 543720
rect 115204 543668 115256 543720
rect 116124 543668 116176 543720
rect 135444 543668 135496 543720
rect 137376 543668 137428 543720
rect 146208 543668 146260 543720
rect 55128 543600 55180 543652
rect 67364 543600 67416 543652
rect 91100 543600 91152 543652
rect 96804 543600 96856 543652
rect 134984 543600 135036 543652
rect 146944 543600 146996 543652
rect 159364 543600 159416 543652
rect 163412 543600 163464 543652
rect 165712 543600 165764 543652
rect 169852 543600 169904 543652
rect 201408 543668 201460 543720
rect 206284 543668 206336 543720
rect 207112 543668 207164 543720
rect 209044 543668 209096 543720
rect 217232 543668 217284 543720
rect 218612 543668 218664 543720
rect 219532 543668 219584 543720
rect 221464 543668 221516 543720
rect 224408 543668 224460 543720
rect 225788 543668 225840 543720
rect 202236 543600 202288 543652
rect 203524 543600 203576 543652
rect 211804 543600 211856 543652
rect 217600 543600 217652 543652
rect 219256 543600 219308 543652
rect 55036 543532 55088 543584
rect 88892 543532 88944 543584
rect 96068 543532 96120 543584
rect 106924 543532 106976 543584
rect 118240 543532 118292 543584
rect 126244 543532 126296 543584
rect 131856 543532 131908 543584
rect 133144 543532 133196 543584
rect 135168 543532 135220 543584
rect 151268 543532 151320 543584
rect 164884 543532 164936 543584
rect 172704 543532 172756 543584
rect 57796 543464 57848 543516
rect 93216 543464 93268 543516
rect 110420 543464 110472 543516
rect 119344 543464 119396 543516
rect 120448 543464 120500 543516
rect 122656 543464 122708 543516
rect 136548 543464 136600 543516
rect 157708 543464 157760 543516
rect 237196 543464 237248 543516
rect 284300 543464 284352 543516
rect 58716 543396 58768 543448
rect 95332 543396 95384 543448
rect 114008 543396 114060 543448
rect 124404 543396 124456 543448
rect 135076 543396 135128 543448
rect 156972 543396 157024 543448
rect 164148 543396 164200 543448
rect 173992 543396 174044 543448
rect 277308 543396 277360 543448
rect 303068 543396 303120 543448
rect 56508 543328 56560 543380
rect 83924 543328 83976 543380
rect 85304 543328 85356 543380
rect 121920 543328 121972 543380
rect 139308 543328 139360 543380
rect 164884 543328 164936 543380
rect 199936 543328 199988 543380
rect 210424 543328 210476 543380
rect 252928 543328 252980 543380
rect 301780 543328 301832 543380
rect 56416 543260 56468 543312
rect 99656 543260 99708 543312
rect 106832 543260 106884 543312
rect 125692 543260 125744 543312
rect 139216 543260 139268 543312
rect 175556 543260 175608 543312
rect 195612 543260 195664 543312
rect 206468 543260 206520 543312
rect 242256 543260 242308 543312
rect 301596 543260 301648 543312
rect 54944 543192 54996 543244
rect 98920 543192 98972 543244
rect 103980 543192 104032 543244
rect 56324 543124 56376 543176
rect 73804 543124 73856 543176
rect 78128 543124 78180 543176
rect 58808 543056 58860 543108
rect 116860 543056 116912 543108
rect 58624 542988 58676 543040
rect 117596 542988 117648 543040
rect 128268 543192 128320 543244
rect 157984 543192 158036 543244
rect 160744 543192 160796 543244
rect 167736 543192 167788 543244
rect 170588 543192 170640 543244
rect 201040 543192 201092 543244
rect 202144 543192 202196 543244
rect 216128 543192 216180 543244
rect 217968 543192 218020 543244
rect 230020 543192 230072 543244
rect 231492 543192 231544 543244
rect 238760 543192 238812 543244
rect 278044 543192 278096 543244
rect 319628 543192 319680 543244
rect 136456 543124 136508 543176
rect 171968 543124 172020 543176
rect 176292 543124 176344 543176
rect 214564 543124 214616 543176
rect 220084 543124 220136 543176
rect 232872 543124 232924 543176
rect 238668 543124 238720 543176
rect 319444 543124 319496 543176
rect 118976 543056 119028 543108
rect 134524 543056 134576 543108
rect 202788 543056 202840 543108
rect 211068 543056 211120 543108
rect 216404 543056 216456 543108
rect 240784 543056 240836 543108
rect 245844 543056 245896 543108
rect 281080 543056 281132 543108
rect 124312 542988 124364 543040
rect 126152 542988 126204 543040
rect 200948 542988 201000 543040
rect 218704 542988 218756 543040
rect 233608 542988 233660 543040
rect 284944 542988 284996 543040
rect 299572 542988 299624 543040
rect 318064 542988 318116 543040
rect 122196 542920 122248 542972
rect 240784 542920 240836 542972
rect 275928 542920 275980 542972
rect 301964 542920 302016 542972
rect 270868 542852 270920 542904
rect 300584 542852 300636 542904
rect 273720 542784 273772 542836
rect 304264 542784 304316 542836
rect 276572 542716 276624 542768
rect 318156 542716 318208 542768
rect 257252 542648 257304 542700
rect 300400 542648 300452 542700
rect 283104 542580 283156 542632
rect 300124 542580 300176 542632
rect 284484 542512 284536 542564
rect 301688 542512 301740 542564
rect 280160 542444 280212 542496
rect 301872 542444 301924 542496
rect 154120 542376 154172 542428
rect 161388 542376 161440 542428
rect 296720 542376 296772 542428
rect 302884 542376 302936 542428
rect 235816 541832 235868 541884
rect 268752 541764 268804 541816
rect 302056 541832 302108 541884
rect 319536 541832 319588 541884
rect 298100 541764 298152 541816
rect 298836 541764 298888 541816
rect 281632 541696 281684 541748
rect 316868 541696 316920 541748
rect 265900 541628 265952 541680
rect 300308 541628 300360 541680
rect 260840 541560 260892 541612
rect 317144 541560 317196 541612
rect 243636 541492 243688 541544
rect 300676 541492 300728 541544
rect 244372 541424 244424 541476
rect 302976 541424 303028 541476
rect 255872 541356 255924 541408
rect 317972 541356 318024 541408
rect 240048 541288 240100 541340
rect 303160 541288 303212 541340
rect 254400 541220 254452 541272
rect 319812 541220 319864 541272
rect 236460 541152 236512 541204
rect 304356 541152 304408 541204
rect 319628 541152 319680 541204
rect 249432 541084 249484 541136
rect 318340 541084 318392 541136
rect 319812 541084 319864 541136
rect 247224 541016 247276 541068
rect 319628 541016 319680 541068
rect 272340 540948 272392 541000
rect 300492 540948 300544 541000
rect 295984 540744 296036 540796
rect 317236 540608 317288 540660
rect 293776 540540 293828 540592
rect 314292 540540 314344 540592
rect 293132 540472 293184 540524
rect 314476 540472 314528 540524
rect 278780 540404 278832 540456
rect 300860 540404 300912 540456
rect 265164 540336 265216 540388
rect 318800 540336 318852 540388
rect 263048 540268 263100 540320
rect 307024 540268 307076 540320
rect 273076 540200 273128 540252
rect 319352 540200 319404 540252
rect 262312 540132 262364 540184
rect 318432 540132 318484 540184
rect 3608 540064 3660 540116
rect 312544 540064 312596 540116
rect 300860 539520 300912 539572
rect 318064 539520 318116 539572
rect 304356 535372 304408 535424
rect 317604 535372 317656 535424
rect 302332 532176 302384 532228
rect 304356 532176 304408 532228
rect 300676 529864 300728 529916
rect 317604 529864 317656 529916
rect 303160 525716 303212 525768
rect 317696 525716 317748 525768
rect 431224 525240 431276 525292
rect 431408 525240 431460 525292
rect 430948 525104 431000 525156
rect 431224 525104 431276 525156
rect 430672 524968 430724 525020
rect 430948 524968 431000 525020
rect 319352 524696 319404 524748
rect 319352 524492 319404 524544
rect 319444 524424 319496 524476
rect 319812 524424 319864 524476
rect 319168 523676 319220 523728
rect 319628 523676 319680 523728
rect 318800 520684 318852 520736
rect 319904 520684 319956 520736
rect 314384 520208 314436 520260
rect 476120 520208 476172 520260
rect 317236 520140 317288 520192
rect 457444 520140 457496 520192
rect 300584 520072 300636 520124
rect 430856 520072 430908 520124
rect 300400 520004 300452 520056
rect 431316 520004 431368 520056
rect 301872 519936 301924 519988
rect 430672 519936 430724 519988
rect 303068 519868 303120 519920
rect 431224 519868 431276 519920
rect 319260 519800 319312 519852
rect 430948 519800 431000 519852
rect 319444 519732 319496 519784
rect 431408 519732 431460 519784
rect 301964 519188 302016 519240
rect 351276 519188 351328 519240
rect 305644 519120 305696 519172
rect 369308 519120 369360 519172
rect 304264 519052 304316 519104
rect 396908 519052 396960 519104
rect 318156 518984 318208 519036
rect 414940 518984 414992 519036
rect 324872 518916 324924 518968
rect 429200 518916 429252 518968
rect 319812 518848 319864 518900
rect 346676 518848 346728 518900
rect 319536 518780 319588 518832
rect 333244 518780 333296 518832
rect 318432 518712 318484 518764
rect 328736 518712 328788 518764
rect 318340 518644 318392 518696
rect 423956 518644 424008 518696
rect 307024 518576 307076 518628
rect 401600 518576 401652 518628
rect 318064 518508 318116 518560
rect 406016 518508 406068 518560
rect 302056 518440 302108 518492
rect 387892 518440 387944 518492
rect 300308 518372 300360 518424
rect 383660 518372 383712 518424
rect 319352 518304 319404 518356
rect 364708 518304 364760 518356
rect 319168 518236 319220 518288
rect 360292 518236 360344 518288
rect 317144 518168 317196 518220
rect 342260 518168 342312 518220
rect 301780 518100 301832 518152
rect 431132 518100 431184 518152
rect 302976 518032 303028 518084
rect 419540 518032 419592 518084
rect 300492 517964 300544 518016
rect 410524 517964 410576 518016
rect 314476 517420 314528 517472
rect 512276 517420 512328 517472
rect 317052 517352 317104 517404
rect 495440 517352 495492 517404
rect 302884 517284 302936 517336
rect 459560 517284 459612 517336
rect 314200 517216 314252 517268
rect 457720 517216 457772 517268
rect 300124 517148 300176 517200
rect 430580 517148 430632 517200
rect 301596 517080 301648 517132
rect 431040 517080 431092 517132
rect 301688 517012 301740 517064
rect 430764 517012 430816 517064
rect 302608 516128 302660 516180
rect 519544 516128 519596 516180
rect 301504 516060 301556 516112
rect 512184 516060 512236 516112
rect 316960 515992 317012 516044
rect 500960 515992 501012 516044
rect 314016 515924 314068 515976
rect 488540 515924 488592 515976
rect 314108 515856 314160 515908
rect 470600 515856 470652 515908
rect 314292 515788 314344 515840
rect 465080 515788 465132 515840
rect 313924 515720 313976 515772
rect 457628 515720 457680 515772
rect 316868 515652 316920 515704
rect 429476 515652 429528 515704
rect 304356 515380 304408 515432
rect 580264 515380 580316 515432
rect 316684 514700 316736 514752
rect 428372 514700 428424 514752
rect 316776 514632 316828 514684
rect 427820 514632 427872 514684
rect 560944 511912 560996 511964
rect 580172 511912 580224 511964
rect 42708 509872 42760 509924
rect 57704 509872 57756 509924
rect 302884 487160 302936 487212
rect 520924 487160 520976 487212
rect 158720 480020 158772 480072
rect 158996 480020 159048 480072
rect 187792 480020 187844 480072
rect 188068 480020 188120 480072
rect 248420 480020 248472 480072
rect 248788 480020 248840 480072
rect 161496 479816 161548 479868
rect 162032 479816 162084 479868
rect 223596 479816 223648 479868
rect 223764 479816 223816 479868
rect 295356 479816 295408 479868
rect 295984 479816 296036 479868
rect 50988 478932 51040 478984
rect 84384 478932 84436 478984
rect 140780 478932 140832 478984
rect 197728 478932 197780 478984
rect 52092 478864 52144 478916
rect 99380 478864 99432 478916
rect 109500 478864 109552 478916
rect 207112 478864 207164 478916
rect 54576 478796 54628 478848
rect 63684 478796 63736 478848
rect 68284 478796 68336 478848
rect 91836 478796 91888 478848
rect 149980 478796 150032 478848
rect 212540 478796 212592 478848
rect 236276 478796 236328 478848
rect 357440 478796 357492 478848
rect 50896 478728 50948 478780
rect 73160 478728 73212 478780
rect 156144 478728 156196 478780
rect 213920 478728 213972 478780
rect 56416 478660 56468 478712
rect 81716 478660 81768 478712
rect 149520 478660 149572 478712
rect 205640 478660 205692 478712
rect 50068 478592 50120 478644
rect 77300 478592 77352 478644
rect 153476 478592 153528 478644
rect 208492 478592 208544 478644
rect 59176 478524 59228 478576
rect 91008 478524 91060 478576
rect 152188 478524 152240 478576
rect 204352 478524 204404 478576
rect 239404 478524 239456 478576
rect 356704 478524 356756 478576
rect 52828 478456 52880 478508
rect 74264 478456 74316 478508
rect 74356 478456 74408 478508
rect 105084 478456 105136 478508
rect 154856 478456 154908 478508
rect 205640 478456 205692 478508
rect 240232 478456 240284 478508
rect 358360 478456 358412 478508
rect 56324 478388 56376 478440
rect 89168 478388 89220 478440
rect 151268 478388 151320 478440
rect 200672 478388 200724 478440
rect 239864 478388 239916 478440
rect 358268 478388 358320 478440
rect 53472 478320 53524 478372
rect 73160 478320 73212 478372
rect 73896 478320 73948 478372
rect 110328 478320 110380 478372
rect 149152 478320 149204 478372
rect 197360 478320 197412 478372
rect 232780 478320 232832 478372
rect 366456 478320 366508 478372
rect 52000 478252 52052 478304
rect 100208 478252 100260 478304
rect 157064 478252 157116 478304
rect 200120 478252 200172 478304
rect 200212 478252 200264 478304
rect 217508 478252 217560 478304
rect 224408 478252 224460 478304
rect 362224 478252 362276 478304
rect 62764 478184 62816 478236
rect 116308 478184 116360 478236
rect 158352 478184 158404 478236
rect 201500 478184 201552 478236
rect 205456 478184 205508 478236
rect 221740 478184 221792 478236
rect 225696 478184 225748 478236
rect 363604 478184 363656 478236
rect 43812 478116 43864 478168
rect 102416 478116 102468 478168
rect 138940 478116 138992 478168
rect 185584 478116 185636 478168
rect 198464 478116 198516 478168
rect 217324 478116 217376 478168
rect 225328 478116 225380 478168
rect 373264 478116 373316 478168
rect 64144 478048 64196 478100
rect 72424 478048 72476 478100
rect 74080 478048 74132 478100
rect 95332 478048 95384 478100
rect 166264 478048 166316 478100
rect 204904 478048 204956 478100
rect 74172 477980 74224 478032
rect 94964 477980 95016 478032
rect 139400 477980 139452 478032
rect 169024 477980 169076 478032
rect 186136 477980 186188 478032
rect 186504 477980 186556 478032
rect 186964 477980 187016 478032
rect 198004 477980 198056 478032
rect 73988 477912 74040 477964
rect 91376 477912 91428 477964
rect 71320 477844 71372 477896
rect 84844 477844 84896 477896
rect 195336 477572 195388 477624
rect 199384 477572 199436 477624
rect 73804 477504 73856 477556
rect 74356 477504 74408 477556
rect 194876 477504 194928 477556
rect 196992 477504 197044 477556
rect 209412 477504 209464 477556
rect 210332 477504 210384 477556
rect 212080 477504 212132 477556
rect 215944 477504 215996 477556
rect 217416 477504 217468 477556
rect 219716 477504 219768 477556
rect 219992 477504 220044 477556
rect 222660 477504 222712 477556
rect 283012 477436 283064 477488
rect 359832 477436 359884 477488
rect 294420 477368 294472 477420
rect 375196 477368 375248 477420
rect 275928 477300 275980 477352
rect 377312 477300 377364 477352
rect 254768 477232 254820 477284
rect 356796 477232 356848 477284
rect 267556 477164 267608 477216
rect 371056 477164 371108 477216
rect 255688 477096 255740 477148
rect 361028 477096 361080 477148
rect 269764 477028 269816 477080
rect 377956 477028 378008 477080
rect 167644 476960 167696 477012
rect 214564 476960 214616 477012
rect 260564 476960 260616 477012
rect 369492 476960 369544 477012
rect 163228 476892 163280 476944
rect 210240 476892 210292 476944
rect 256608 476892 256660 476944
rect 368112 476892 368164 476944
rect 60556 476824 60608 476876
rect 133144 476824 133196 476876
rect 164056 476824 164108 476876
rect 214656 476824 214708 476876
rect 242900 476824 242952 476876
rect 363788 476824 363840 476876
rect 14464 476756 14516 476808
rect 378140 476756 378192 476808
rect 70400 476076 70452 476128
rect 70860 476076 70912 476128
rect 85580 476076 85632 476128
rect 85764 476076 85816 476128
rect 51908 476008 51960 476060
rect 98460 476008 98512 476060
rect 48044 475940 48096 475992
rect 97172 475940 97224 475992
rect 178132 475940 178184 475992
rect 203524 475940 203576 475992
rect 49056 475872 49108 475924
rect 98000 475872 98052 475924
rect 186504 475872 186556 475924
rect 212080 475872 212132 475924
rect 283840 475872 283892 475924
rect 359924 475872 359976 475924
rect 59820 475804 59872 475856
rect 119620 475804 119672 475856
rect 165436 475804 165488 475856
rect 211804 475804 211856 475856
rect 294880 475804 294932 475856
rect 379152 475804 379204 475856
rect 48136 475736 48188 475788
rect 111708 475736 111760 475788
rect 160100 475736 160152 475788
rect 210424 475736 210476 475788
rect 272432 475736 272484 475788
rect 367008 475736 367060 475788
rect 47860 475668 47912 475720
rect 112076 475668 112128 475720
rect 137652 475668 137704 475720
rect 198096 475668 198148 475720
rect 271512 475668 271564 475720
rect 371792 475668 371844 475720
rect 46388 475600 46440 475652
rect 111248 475600 111300 475652
rect 138572 475600 138624 475652
rect 200396 475600 200448 475652
rect 270224 475600 270276 475652
rect 376484 475600 376536 475652
rect 48964 475532 49016 475584
rect 115204 475532 115256 475584
rect 138112 475532 138164 475584
rect 200304 475532 200356 475584
rect 260932 475532 260984 475584
rect 374920 475532 374972 475584
rect 46756 475464 46808 475516
rect 115664 475464 115716 475516
rect 135904 475464 135956 475516
rect 197820 475464 197872 475516
rect 209964 475464 210016 475516
rect 210148 475464 210200 475516
rect 211252 475464 211304 475516
rect 246396 475464 246448 475516
rect 365168 475464 365220 475516
rect 49148 475396 49200 475448
rect 120080 475396 120132 475448
rect 122840 475396 122892 475448
rect 123668 475396 123720 475448
rect 136732 475396 136784 475448
rect 199660 475396 199712 475448
rect 60740 475328 60792 475380
rect 61108 475328 61160 475380
rect 62120 475328 62172 475380
rect 62948 475328 63000 475380
rect 63040 475328 63092 475380
rect 134984 475328 135036 475380
rect 139400 475328 139452 475380
rect 140044 475328 140096 475380
rect 140872 475328 140924 475380
rect 141700 475328 141752 475380
rect 54760 475260 54812 475312
rect 96712 475260 96764 475312
rect 100852 475260 100904 475312
rect 101588 475260 101640 475312
rect 103612 475260 103664 475312
rect 103796 475260 103848 475312
rect 104992 475260 105044 475312
rect 105636 475260 105688 475312
rect 106372 475260 106424 475312
rect 106556 475260 106608 475312
rect 113272 475260 113324 475312
rect 113548 475260 113600 475312
rect 122932 475260 122984 475312
rect 123300 475260 123352 475312
rect 124220 475260 124272 475312
rect 124956 475260 125008 475312
rect 125600 475260 125652 475312
rect 126336 475260 126388 475312
rect 140780 475260 140832 475312
rect 141332 475260 141384 475312
rect 58808 475192 58860 475244
rect 96252 475192 96304 475244
rect 103520 475192 103572 475244
rect 104348 475192 104400 475244
rect 106280 475192 106332 475244
rect 106924 475192 106976 475244
rect 135444 475192 135496 475244
rect 143632 475260 143684 475312
rect 144460 475260 144512 475312
rect 146300 475260 146352 475312
rect 146668 475260 146720 475312
rect 165620 475260 165672 475312
rect 166356 475260 166408 475312
rect 168380 475260 168432 475312
rect 169116 475260 169168 475312
rect 172520 475260 172572 475312
rect 173532 475260 173584 475312
rect 173900 475260 173952 475312
rect 174268 475260 174320 475312
rect 175280 475260 175332 475312
rect 176108 475260 176160 475312
rect 205732 475328 205784 475380
rect 206468 475328 206520 475380
rect 207204 475328 207256 475380
rect 207756 475328 207808 475380
rect 209780 475328 209832 475380
rect 210516 475328 210568 475380
rect 238116 475396 238168 475448
rect 362408 475396 362460 475448
rect 212724 475328 212776 475380
rect 213092 475328 213144 475380
rect 213920 475328 213972 475380
rect 214932 475328 214984 475380
rect 215392 475328 215444 475380
rect 216220 475328 216272 475380
rect 218060 475328 218112 475380
rect 218796 475328 218848 475380
rect 219440 475328 219492 475380
rect 220084 475328 220136 475380
rect 223580 475328 223632 475380
rect 224500 475328 224552 475380
rect 226340 475328 226392 475380
rect 226708 475328 226760 475380
rect 227720 475328 227772 475380
rect 228548 475328 228600 475380
rect 229100 475328 229152 475380
rect 229468 475328 229520 475380
rect 240140 475328 240192 475380
rect 240876 475328 240928 475380
rect 244280 475328 244332 475380
rect 244740 475328 244792 475380
rect 247132 475328 247184 475380
rect 247500 475328 247552 475380
rect 203708 475260 203760 475312
rect 209504 475260 209556 475312
rect 211252 475260 211304 475312
rect 212540 475260 212592 475312
rect 213460 475260 213512 475312
rect 215300 475260 215352 475312
rect 215668 475260 215720 475312
rect 244372 475260 244424 475312
rect 244556 475260 244608 475312
rect 247040 475260 247092 475312
rect 247868 475260 247920 475312
rect 198188 475192 198240 475244
rect 210332 475192 210384 475244
rect 220820 475192 220872 475244
rect 221004 475192 221056 475244
rect 242072 475192 242124 475244
rect 369124 475328 369176 475380
rect 248512 475260 248564 475312
rect 249156 475260 249208 475312
rect 262220 475260 262272 475312
rect 262404 475260 262456 475312
rect 263600 475260 263652 475312
rect 264244 475260 264296 475312
rect 264980 475260 265032 475312
rect 265900 475260 265952 475312
rect 292580 475260 292632 475312
rect 293316 475260 293368 475312
rect 296720 475260 296772 475312
rect 297732 475260 297784 475312
rect 59728 475124 59780 475176
rect 97540 475124 97592 475176
rect 142160 475124 142212 475176
rect 142620 475124 142672 475176
rect 57336 475056 57388 475108
rect 63040 475056 63092 475108
rect 66260 475056 66312 475108
rect 66812 475056 66864 475108
rect 67824 475056 67876 475108
rect 68652 475056 68704 475108
rect 71780 475056 71832 475108
rect 72608 475056 72660 475108
rect 74540 475056 74592 475108
rect 75276 475056 75328 475108
rect 78772 475056 78824 475108
rect 79692 475056 79744 475108
rect 92572 475056 92624 475108
rect 93308 475056 93360 475108
rect 67640 474988 67692 475040
rect 67916 474988 67968 475040
rect 210332 474988 210384 475040
rect 297088 474580 297140 474632
rect 362776 474580 362828 474632
rect 282552 474512 282604 474564
rect 375104 474512 375156 474564
rect 272892 474444 272944 474496
rect 369676 474444 369728 474496
rect 282092 474376 282144 474428
rect 379980 474376 380032 474428
rect 265256 474308 265308 474360
rect 369584 474308 369636 474360
rect 254400 474240 254452 474292
rect 358452 474240 358504 474292
rect 265348 474172 265400 474224
rect 372160 474172 372212 474224
rect 205916 474104 205968 474156
rect 217324 474104 217376 474156
rect 260104 474104 260156 474156
rect 368204 474104 368256 474156
rect 176016 474036 176068 474088
rect 206560 474036 206612 474088
rect 246028 474036 246080 474088
rect 369216 474036 369268 474088
rect 57888 473968 57940 474020
rect 114284 473968 114336 474020
rect 159640 473968 159692 474020
rect 216036 473968 216088 474020
rect 237196 473968 237248 474020
rect 366732 473968 366784 474020
rect 48228 473288 48280 473340
rect 117872 473288 117924 473340
rect 46572 473220 46624 473272
rect 116492 473220 116544 473272
rect 49240 473152 49292 473204
rect 119160 473152 119212 473204
rect 284760 473152 284812 473204
rect 360016 473152 360068 473204
rect 45468 473084 45520 473136
rect 118240 473084 118292 473136
rect 295984 473084 296036 473136
rect 372620 473084 372672 473136
rect 53564 473016 53616 473068
rect 131948 473016 132000 473068
rect 274180 473016 274232 473068
rect 362868 473016 362920 473068
rect 57060 472948 57112 473000
rect 136364 472948 136416 473000
rect 192116 472948 192168 473000
rect 192668 472948 192720 473000
rect 261852 472948 261904 473000
rect 372252 472948 372304 473000
rect 50160 472880 50212 472932
rect 131488 472880 131540 472932
rect 182272 472880 182324 472932
rect 183100 472880 183152 472932
rect 242440 472880 242492 472932
rect 360936 472880 360988 472932
rect 48872 472812 48924 472864
rect 129740 472812 129792 472864
rect 245568 472812 245620 472864
rect 370688 472812 370740 472864
rect 47768 472744 47820 472796
rect 131028 472744 131080 472796
rect 234988 472744 235040 472796
rect 364984 472744 365036 472796
rect 46296 472676 46348 472728
rect 130568 472676 130620 472728
rect 172428 472676 172480 472728
rect 210608 472676 210660 472728
rect 238944 472676 238996 472728
rect 378784 472676 378836 472728
rect 46112 472608 46164 472660
rect 143816 472608 143868 472660
rect 147772 472608 147824 472660
rect 218704 472608 218756 472660
rect 227536 472608 227588 472660
rect 371884 472608 371936 472660
rect 46664 472540 46716 472592
rect 116952 472540 117004 472592
rect 50436 472472 50488 472524
rect 116032 472472 116084 472524
rect 58624 472404 58676 472456
rect 118700 472404 118752 472456
rect 258080 472064 258132 472116
rect 258908 472064 258960 472116
rect 280252 471928 280304 471980
rect 280436 471928 280488 471980
rect 292212 471928 292264 471980
rect 368296 471928 368348 471980
rect 269304 471860 269356 471912
rect 356888 471860 356940 471912
rect 263784 471792 263836 471844
rect 365352 471792 365404 471844
rect 258356 471724 258408 471776
rect 362592 471724 362644 471776
rect 273720 471656 273772 471708
rect 378048 471656 378100 471708
rect 270684 471588 270736 471640
rect 377680 471588 377732 471640
rect 252192 471520 252244 471572
rect 361212 471520 361264 471572
rect 198924 471452 198976 471504
rect 199108 471452 199160 471504
rect 263140 471452 263192 471504
rect 375012 471452 375064 471504
rect 180340 471384 180392 471436
rect 209228 471384 209280 471436
rect 237656 471384 237708 471436
rect 367744 471384 367796 471436
rect 57244 471316 57296 471368
rect 129280 471316 129332 471368
rect 162032 471316 162084 471368
rect 211896 471316 211948 471368
rect 246856 471316 246908 471368
rect 378876 471316 378928 471368
rect 61936 471248 61988 471300
rect 81532 471180 81584 471232
rect 82268 471180 82320 471232
rect 82820 471180 82872 471232
rect 83004 471180 83056 471232
rect 85672 471180 85724 471232
rect 86316 471180 86368 471232
rect 189172 471180 189224 471232
rect 189724 471180 189776 471232
rect 192024 471180 192076 471232
rect 192852 471180 192904 471232
rect 193220 471180 193272 471232
rect 193772 471180 193824 471232
rect 196716 471248 196768 471300
rect 196900 471248 196952 471300
rect 197360 471248 197412 471300
rect 197636 471248 197688 471300
rect 198740 471248 198792 471300
rect 199476 471248 199528 471300
rect 201500 471248 201552 471300
rect 201684 471248 201736 471300
rect 203064 471248 203116 471300
rect 203892 471248 203944 471300
rect 204352 471248 204404 471300
rect 205180 471248 205232 471300
rect 199200 471180 199252 471232
rect 202880 471180 202932 471232
rect 203156 471180 203208 471232
rect 204996 471180 205048 471232
rect 217692 471248 217744 471300
rect 227904 471248 227956 471300
rect 362316 471248 362368 471300
rect 277400 471180 277452 471232
rect 277860 471180 277912 471232
rect 278780 471180 278832 471232
rect 279148 471180 279200 471232
rect 287060 471180 287112 471232
rect 287980 471180 288032 471232
rect 191840 471112 191892 471164
rect 192392 471112 192444 471164
rect 193312 471112 193364 471164
rect 194140 471112 194192 471164
rect 287428 471112 287480 471164
rect 361304 471180 361356 471232
rect 82820 471044 82872 471096
rect 83556 471044 83608 471096
rect 55680 470500 55732 470552
rect 128360 470500 128412 470552
rect 54392 470432 54444 470484
rect 127072 470432 127124 470484
rect 57152 470364 57204 470416
rect 132776 470364 132828 470416
rect 275192 470364 275244 470416
rect 359464 470364 359516 470416
rect 43904 470296 43956 470348
rect 122840 470296 122892 470348
rect 187700 470296 187752 470348
rect 188436 470296 188488 470348
rect 274732 470296 274784 470348
rect 364156 470296 364208 470348
rect 42432 470228 42484 470280
rect 122932 470228 122984 470280
rect 286048 470228 286100 470280
rect 376760 470228 376812 470280
rect 43720 470160 43772 470212
rect 124404 470160 124456 470212
rect 265072 470160 265124 470212
rect 362684 470160 362736 470212
rect 42340 470092 42392 470144
rect 123024 470092 123076 470144
rect 256884 470092 256936 470144
rect 366824 470092 366876 470144
rect 51540 470024 51592 470076
rect 133972 470024 134024 470076
rect 244464 470024 244516 470076
rect 371976 470024 372028 470076
rect 48780 469956 48832 470008
rect 133420 469956 133472 470008
rect 236000 469956 236052 470008
rect 365076 469956 365128 470008
rect 46204 469888 46256 469940
rect 132868 469888 132920 469940
rect 178132 469888 178184 469940
rect 214840 469888 214892 469940
rect 227812 469888 227864 469940
rect 358176 469888 358228 469940
rect 43444 469820 43496 469872
rect 132132 469820 132184 469872
rect 158812 469820 158864 469872
rect 207664 469820 207716 469872
rect 229284 469820 229336 469872
rect 374644 469820 374696 469872
rect 58532 469752 58584 469804
rect 127164 469752 127216 469804
rect 58440 469684 58492 469736
rect 126980 469684 127032 469736
rect 280896 469140 280948 469192
rect 364064 469140 364116 469192
rect 264980 469072 265032 469124
rect 358544 469072 358596 469124
rect 42156 469004 42208 469056
rect 62212 469004 62264 469056
rect 273260 469004 273312 469056
rect 372436 469004 372488 469056
rect 47952 468936 48004 468988
rect 73896 468936 73948 468988
rect 270500 468936 270552 468988
rect 373172 468936 373224 468988
rect 42524 468868 42576 468920
rect 73988 468868 74040 468920
rect 259460 468868 259512 468920
rect 370872 468868 370924 468920
rect 41328 468800 41380 468852
rect 74080 468800 74132 468852
rect 256792 468800 256844 468852
rect 370964 468800 371016 468852
rect 39856 468732 39908 468784
rect 74172 468732 74224 468784
rect 175372 468732 175424 468784
rect 207848 468732 207900 468784
rect 251272 468732 251324 468784
rect 368020 468732 368072 468784
rect 43628 468664 43680 468716
rect 103704 468664 103756 468716
rect 169024 468664 169076 468716
rect 205916 468664 205968 468716
rect 244372 468664 244424 468716
rect 366548 468664 366600 468716
rect 45376 468596 45428 468648
rect 106464 468596 106516 468648
rect 165712 468596 165764 468648
rect 218796 468596 218848 468648
rect 241520 468596 241572 468648
rect 367836 468596 367888 468648
rect 45284 468528 45336 468580
rect 106372 468528 106424 468580
rect 139492 468528 139544 468580
rect 207480 468528 207532 468580
rect 227720 468528 227772 468580
rect 360844 468528 360896 468580
rect 60832 468460 60884 468512
rect 214196 468460 214248 468512
rect 226432 468460 226484 468512
rect 376024 468460 376076 468512
rect 291476 468392 291528 468444
rect 371700 468392 371752 468444
rect 88524 468120 88576 468172
rect 89260 468120 89312 468172
rect 88432 467984 88484 468036
rect 88708 467984 88760 468036
rect 274640 467712 274692 467764
rect 358728 467712 358780 467764
rect 290188 467644 290240 467696
rect 376668 467644 376720 467696
rect 285772 467576 285824 467628
rect 286692 467576 286744 467628
rect 290556 467576 290608 467628
rect 379244 467576 379296 467628
rect 266452 467508 266504 467560
rect 359648 467508 359700 467560
rect 267924 467440 267976 467492
rect 361396 467440 361448 467492
rect 256700 467372 256752 467424
rect 365444 467372 365496 467424
rect 262312 467304 262364 467356
rect 378968 467304 379020 467356
rect 57796 467236 57848 467288
rect 113272 467236 113324 467288
rect 175280 467236 175332 467288
rect 205088 467236 205140 467288
rect 242992 467236 243044 467288
rect 373356 467236 373408 467288
rect 45192 467168 45244 467220
rect 106280 467168 106332 467220
rect 160192 467168 160244 467220
rect 202144 467168 202196 467220
rect 229192 467168 229244 467220
rect 363696 467168 363748 467220
rect 59360 467100 59412 467152
rect 179512 467100 179564 467152
rect 186412 467100 186464 467152
rect 203708 467100 203760 467152
rect 207296 467100 207348 467152
rect 217784 467100 217836 467152
rect 223672 467100 223724 467152
rect 370504 467100 370556 467152
rect 50620 466352 50672 466404
rect 83004 466352 83056 466404
rect 189172 466352 189224 466404
rect 206284 466352 206336 466404
rect 49424 466284 49476 466336
rect 82912 466284 82964 466336
rect 183652 466284 183704 466336
rect 200764 466284 200816 466336
rect 298192 466284 298244 466336
rect 357072 466284 357124 466336
rect 56508 466216 56560 466268
rect 103612 466216 103664 466268
rect 183744 466216 183796 466268
rect 205180 466216 205232 466268
rect 298284 466216 298336 466268
rect 369860 466216 369912 466268
rect 51816 466148 51868 466200
rect 99472 466148 99524 466200
rect 182456 466148 182508 466200
rect 209320 466148 209372 466200
rect 299480 466148 299532 466200
rect 373816 466148 373868 466200
rect 53196 466080 53248 466132
rect 100944 466080 100996 466132
rect 189264 466080 189316 466132
rect 216404 466080 216456 466132
rect 289820 466080 289872 466132
rect 365536 466080 365588 466132
rect 53104 466012 53156 466064
rect 100852 466012 100904 466064
rect 174084 466012 174136 466064
rect 210792 466012 210844 466064
rect 288624 466012 288676 466064
rect 368388 466012 368440 466064
rect 50252 465944 50304 465996
rect 98184 465944 98236 465996
rect 139400 465944 139452 465996
rect 197084 465944 197136 465996
rect 288532 465944 288584 465996
rect 376576 465944 376628 465996
rect 58716 465876 58768 465928
rect 110604 465876 110656 465928
rect 140964 465876 141016 465928
rect 200580 465876 200632 465928
rect 249984 465876 250036 465928
rect 366640 465876 366692 465928
rect 45008 465808 45060 465860
rect 105084 465808 105136 465860
rect 140780 465808 140832 465860
rect 203156 465808 203208 465860
rect 251180 465808 251232 465860
rect 369308 465808 369360 465860
rect 45100 465740 45152 465792
rect 104992 465740 105044 465792
rect 140872 465740 140924 465792
rect 204444 465740 204496 465792
rect 240232 465740 240284 465792
rect 373448 465740 373500 465792
rect 43536 465672 43588 465724
rect 103520 465672 103572 465724
rect 125784 465672 125836 465724
rect 201592 465672 201644 465724
rect 226340 465672 226392 465724
rect 370596 465672 370648 465724
rect 52276 465604 52328 465656
rect 82820 465604 82872 465656
rect 192024 465604 192076 465656
rect 199568 465604 199620 465656
rect 44732 465536 44784 465588
rect 65064 465536 65116 465588
rect 44824 465468 44876 465520
rect 64972 465468 65024 465520
rect 190644 465468 190696 465520
rect 203892 465604 203944 465656
rect 192668 465400 192720 465452
rect 201040 465400 201092 465452
rect 288440 464924 288492 464976
rect 357256 464924 357308 464976
rect 292672 464856 292724 464908
rect 365628 464856 365680 464908
rect 292764 464788 292816 464840
rect 366272 464788 366324 464840
rect 292580 464720 292632 464772
rect 369032 464720 369084 464772
rect 284392 464652 284444 464704
rect 362040 464652 362092 464704
rect 285680 464584 285732 464636
rect 363512 464584 363564 464636
rect 291200 464516 291252 464568
rect 370412 464516 370464 464568
rect 293960 464448 294012 464500
rect 376852 464448 376904 464500
rect 57428 464380 57480 464432
rect 114744 464380 114796 464432
rect 285864 464380 285916 464432
rect 375380 464380 375432 464432
rect 42248 464312 42300 464364
rect 102324 464312 102376 464364
rect 285772 464312 285824 464364
rect 379336 464312 379388 464364
rect 56048 463632 56100 463684
rect 86960 463632 87012 463684
rect 176844 463632 176896 463684
rect 200856 463632 200908 463684
rect 287152 463632 287204 463684
rect 360752 463632 360804 463684
rect 49332 463564 49384 463616
rect 81624 463564 81676 463616
rect 193404 463564 193456 463616
rect 217600 463564 217652 463616
rect 277492 463564 277544 463616
rect 357164 463564 357216 463616
rect 56232 463496 56284 463548
rect 88616 463496 88668 463548
rect 180984 463496 181036 463548
rect 206652 463496 206704 463548
rect 276204 463496 276256 463548
rect 361488 463496 361540 463548
rect 54944 463428 54996 463480
rect 87144 463428 87196 463480
rect 178040 463428 178092 463480
rect 216128 463428 216180 463480
rect 276112 463428 276164 463480
rect 364892 463428 364944 463480
rect 53288 463360 53340 463412
rect 85672 463360 85724 463412
rect 169760 463360 169812 463412
rect 209136 463360 209188 463412
rect 280252 463360 280304 463412
rect 370320 463360 370372 463412
rect 55128 463292 55180 463344
rect 88524 463292 88576 463344
rect 161572 463292 161624 463344
rect 204996 463292 205048 463344
rect 277584 463292 277636 463344
rect 368940 463292 368992 463344
rect 55036 463224 55088 463276
rect 88432 463224 88484 463276
rect 161480 463224 161532 463276
rect 210700 463224 210752 463276
rect 267832 463224 267884 463276
rect 359556 463224 359608 463276
rect 56140 463156 56192 463208
rect 89812 463156 89864 463208
rect 142344 463156 142396 463208
rect 200488 463156 200540 463208
rect 278964 463156 279016 463208
rect 374460 463156 374512 463208
rect 57612 463088 57664 463140
rect 113364 463088 113416 463140
rect 142252 463088 142304 463140
rect 208584 463088 208636 463140
rect 249892 463088 249944 463140
rect 365260 463088 365312 463140
rect 53380 463020 53432 463072
rect 87052 463020 87104 463072
rect 107752 463020 107804 463072
rect 201868 463020 201920 463072
rect 249800 463020 249852 463072
rect 372068 463020 372120 463072
rect 53012 462952 53064 463004
rect 100760 462952 100812 463004
rect 109132 462952 109184 463004
rect 205640 462952 205692 463004
rect 240140 462952 240192 463004
rect 362500 462952 362552 463004
rect 54852 462884 54904 462936
rect 85580 462884 85632 462936
rect 189080 462884 189132 462936
rect 212264 462884 212316 462936
rect 284300 462884 284352 462936
rect 357808 462884 357860 462936
rect 47584 462816 47636 462868
rect 64880 462816 64932 462868
rect 182364 462816 182416 462868
rect 202328 462816 202380 462868
rect 47676 462748 47728 462800
rect 63684 462748 63736 462800
rect 193312 462748 193364 462800
rect 213092 462748 213144 462800
rect 133144 462272 133196 462324
rect 178316 462272 178368 462324
rect 185584 462136 185636 462188
rect 203248 462136 203300 462188
rect 190552 462068 190604 462120
rect 208952 462068 209004 462120
rect 282920 462068 282972 462120
rect 358084 462068 358136 462120
rect 176752 462000 176804 462052
rect 202236 462000 202288 462052
rect 296720 462000 296772 462052
rect 374000 462000 374052 462052
rect 184940 461932 184992 461984
rect 213276 461932 213328 461984
rect 278872 461932 278924 461984
rect 357992 461932 358044 461984
rect 182272 461864 182324 461916
rect 212172 461864 212224 461916
rect 277400 461864 277452 461916
rect 366180 461864 366232 461916
rect 180892 461796 180944 461848
rect 213368 461796 213420 461848
rect 253940 461796 253992 461848
rect 363972 461796 364024 461848
rect 179512 461728 179564 461780
rect 212908 461728 212960 461780
rect 260840 461728 260892 461780
rect 376392 461728 376444 461780
rect 57704 461660 57756 461712
rect 111892 461660 111944 461712
rect 158720 461660 158772 461712
rect 206468 461660 206520 461712
rect 252560 461660 252612 461712
rect 373632 461660 373684 461712
rect 52184 461592 52236 461644
rect 71044 461592 71096 461644
rect 107660 461592 107712 461644
rect 198280 461592 198332 461644
rect 252652 461592 252704 461644
rect 376208 461592 376260 461644
rect 498200 461116 498252 461168
rect 517704 461116 517756 461168
rect 339776 461048 339828 461100
rect 356980 461048 357032 461100
rect 178316 460980 178368 461032
rect 201960 460980 202012 461032
rect 338304 460980 338356 461032
rect 362960 460980 363012 461032
rect 190920 460912 190972 460964
rect 207020 460912 207072 460964
rect 212908 460912 212960 460964
rect 339776 460912 339828 460964
rect 351000 460912 351052 460964
rect 360200 460912 360252 460964
rect 499856 460980 499908 461032
rect 517612 460980 517664 461032
rect 498200 460912 498252 460964
rect 510896 460912 510948 460964
rect 517520 460912 517572 460964
rect 50712 460844 50764 460896
rect 80060 460844 80112 460896
rect 287060 460844 287112 460896
rect 367652 460844 367704 460896
rect 53748 460776 53800 460828
rect 78772 460776 78824 460828
rect 179420 460776 179472 460828
rect 218980 460776 219032 460828
rect 262220 460776 262272 460828
rect 361120 460776 361172 460828
rect 53656 460708 53708 460760
rect 66352 460708 66404 460760
rect 258172 460708 258224 460760
rect 363880 460708 363932 460760
rect 43260 460640 43312 460692
rect 60740 460640 60792 460692
rect 183560 460640 183612 460692
rect 203800 460640 203852 460692
rect 267740 460640 267792 460692
rect 373724 460640 373776 460692
rect 43352 460572 43404 460624
rect 62120 460572 62172 460624
rect 187792 460572 187844 460624
rect 209412 460572 209464 460624
rect 248604 460572 248656 460624
rect 367928 460572 367980 460624
rect 49516 460504 49568 460556
rect 70400 460504 70452 460556
rect 180800 460504 180852 460556
rect 205272 460504 205324 460556
rect 248420 460504 248472 460556
rect 370780 460504 370832 460556
rect 39948 460436 40000 460488
rect 66260 460436 66312 460488
rect 193220 460436 193272 460488
rect 219164 460436 219216 460488
rect 248512 460436 248564 460488
rect 373540 460436 373592 460488
rect 44916 460368 44968 460420
rect 73804 460368 73856 460420
rect 168472 460368 168524 460420
rect 206376 460368 206428 460420
rect 244280 460368 244332 460420
rect 369400 460368 369452 460420
rect 49608 460300 49660 460352
rect 78864 460300 78916 460352
rect 165620 460300 165672 460352
rect 203616 460300 203668 460352
rect 247224 460300 247276 460352
rect 376116 460300 376168 460352
rect 50528 460232 50580 460284
rect 92572 460232 92624 460284
rect 247132 460232 247184 460284
rect 376300 460232 376352 460284
rect 44088 460164 44140 460216
rect 71780 460164 71832 460216
rect 72424 460164 72476 460216
rect 199016 460164 199068 460216
rect 237380 460164 237432 460216
rect 374736 460164 374788 460216
rect 59268 460096 59320 460148
rect 67732 460096 67784 460148
rect 59912 460028 59964 460080
rect 68284 460028 68336 460080
rect 194600 459620 194652 459672
rect 199476 459620 199528 459672
rect 215760 459620 215812 459672
rect 220912 459620 220964 459672
rect 218612 459552 218664 459604
rect 221004 459552 221056 459604
rect 187700 459484 187752 459536
rect 200948 459484 201000 459536
rect 191840 459416 191892 459468
rect 205364 459416 205416 459468
rect 295340 459416 295392 459468
rect 357900 459416 357952 459468
rect 190460 459348 190512 459400
rect 208032 459348 208084 459400
rect 298100 459348 298152 459400
rect 364248 459348 364300 459400
rect 58900 459280 58952 459332
rect 92480 459280 92532 459332
rect 182180 459280 182232 459332
rect 207940 459280 207992 459332
rect 281540 459280 281592 459332
rect 359740 459280 359792 459332
rect 55956 459212 56008 459264
rect 89904 459212 89956 459264
rect 173992 459212 174044 459264
rect 206744 459212 206796 459264
rect 280160 459212 280212 459264
rect 362132 459212 362184 459264
rect 57520 459144 57572 459196
rect 111984 459144 112036 459196
rect 176660 459144 176712 459196
rect 210884 459144 210936 459196
rect 276020 459144 276072 459196
rect 367560 459144 367612 459196
rect 54668 459076 54720 459128
rect 117504 459076 117556 459128
rect 173900 459076 173952 459128
rect 216220 459076 216272 459128
rect 271880 459076 271932 459128
rect 364800 459076 364852 459128
rect 51724 459008 51776 459060
rect 121460 459008 121512 459060
rect 125600 459008 125652 459060
rect 197544 459008 197596 459060
rect 263600 459008 263652 459060
rect 366916 459008 366968 459060
rect 55772 458940 55824 458992
rect 130016 458940 130068 458992
rect 136640 458940 136692 458992
rect 199108 458940 199160 458992
rect 258080 458940 258132 458992
rect 372344 458940 372396 458992
rect 54484 458872 54536 458924
rect 134064 458872 134116 458924
rect 142160 458872 142212 458924
rect 211344 458872 211396 458924
rect 242900 458872 242952 458924
rect 374828 458872 374880 458924
rect 52920 458804 52972 458856
rect 99564 458804 99616 458856
rect 109316 458804 109368 458856
rect 197636 458804 197688 458856
rect 247040 458804 247092 458856
rect 379060 458804 379112 458856
rect 191932 458736 191984 458788
rect 202420 458736 202472 458788
rect 199016 458328 199068 458380
rect 46020 458260 46072 458312
rect 358820 458260 358872 458312
rect 516600 458260 516652 458312
rect 207388 458192 207440 458244
rect 208124 458192 208176 458244
rect 204352 457444 204404 457496
rect 217876 457444 217928 457496
rect 50712 456084 50764 456136
rect 50988 456084 51040 456136
rect 356612 456084 356664 456136
rect 356980 456084 357032 456136
rect 519544 454656 519596 454708
rect 580264 454656 580316 454708
rect 54392 414196 54444 414248
rect 55588 414196 55640 414248
rect 205824 413924 205876 413976
rect 207296 413924 207348 413976
rect 208124 413244 208176 413296
rect 216956 413244 217008 413296
rect 46020 412564 46072 412616
rect 56968 412564 57020 412616
rect 54392 411884 54444 411936
rect 58440 411884 58492 411936
rect 199660 411884 199712 411936
rect 205824 411884 205876 411936
rect 363512 411884 363564 411936
rect 377036 411884 377088 411936
rect 2964 411204 3016 411256
rect 14464 411204 14516 411256
rect 57060 410796 57112 410848
rect 58440 410796 58492 410848
rect 198096 410524 198148 410576
rect 199292 410524 199344 410576
rect 362040 410524 362092 410576
rect 377220 410524 377272 410576
rect 44640 409844 44692 409896
rect 57060 409844 57112 409896
rect 53564 409776 53616 409828
rect 56876 409776 56928 409828
rect 205732 409096 205784 409148
rect 216680 409096 216732 409148
rect 360016 409096 360068 409148
rect 377220 409096 377272 409148
rect 47492 408484 47544 408536
rect 57060 408484 57112 408536
rect 373908 407804 373960 407856
rect 376852 407804 376904 407856
rect 207296 407736 207348 407788
rect 216680 407736 216732 407788
rect 357808 407736 357860 407788
rect 377128 407736 377180 407788
rect 47400 407124 47452 407176
rect 56968 407124 57020 407176
rect 359924 406376 359976 406428
rect 377220 406376 377272 406428
rect 53564 405696 53616 405748
rect 57060 405696 57112 405748
rect 375932 405628 375984 405680
rect 376760 405628 376812 405680
rect 377680 405628 377732 405680
rect 378600 405628 378652 405680
rect 358084 404948 358136 405000
rect 377588 404948 377640 405000
rect 51632 404336 51684 404388
rect 57060 404336 57112 404388
rect 51724 404268 51776 404320
rect 53840 404268 53892 404320
rect 359832 403588 359884 403640
rect 377680 403588 377732 403640
rect 52368 402976 52420 403028
rect 56968 402976 57020 403028
rect 199660 393932 199712 393984
rect 214196 393932 214248 393984
rect 198188 393388 198240 393440
rect 198372 393320 198424 393372
rect 200580 393320 200632 393372
rect 200580 393184 200632 393236
rect 199568 391212 199620 391264
rect 211528 391212 211580 391264
rect 377404 388696 377456 388748
rect 377772 388696 377824 388748
rect 216772 388560 216824 388612
rect 216956 388560 217008 388612
rect 520924 388424 520976 388476
rect 580356 388424 580408 388476
rect 46112 384956 46164 385008
rect 56968 384956 57020 385008
rect 209504 384956 209556 385008
rect 216680 384956 216732 385008
rect 359740 384956 359792 385008
rect 376944 384956 376996 385008
rect 56968 383596 57020 383648
rect 57152 383596 57204 383648
rect 57244 383596 57296 383648
rect 57336 383596 57388 383648
rect 207020 383596 207072 383648
rect 216680 383596 216732 383648
rect 360200 383596 360252 383648
rect 376944 383596 376996 383648
rect 57152 383460 57204 383512
rect 57244 383460 57296 383512
rect 359648 383528 359700 383580
rect 376852 383528 376904 383580
rect 216864 383460 216916 383512
rect 217324 383460 217376 383512
rect 212264 383324 212316 383376
rect 216864 383324 216916 383376
rect 358084 382236 358136 382288
rect 360200 382236 360252 382288
rect 42708 382168 42760 382220
rect 56876 382168 56928 382220
rect 57244 382168 57296 382220
rect 212632 379788 212684 379840
rect 213460 379788 213512 379840
rect 51724 379516 51776 379568
rect 53840 379516 53892 379568
rect 218060 378768 218112 378820
rect 218336 378768 218388 378820
rect 57152 378564 57204 378616
rect 57336 378564 57388 378616
rect 53564 375368 53616 375420
rect 53748 375300 53800 375352
rect 197176 375300 197228 375352
rect 198188 375300 198240 375352
rect 217232 375300 217284 375352
rect 217784 375300 217836 375352
rect 51632 375028 51684 375080
rect 217232 375028 217284 375080
rect 53748 374960 53800 375012
rect 217324 374960 217376 375012
rect 375196 374960 375248 375012
rect 380900 374960 380952 375012
rect 56508 374892 56560 374944
rect 60740 374892 60792 374944
rect 200212 374756 200264 374808
rect 304264 374756 304316 374808
rect 200672 374688 200724 374740
rect 305000 374688 305052 374740
rect 375380 374688 375432 374740
rect 201684 374620 201736 374672
rect 311808 374620 311860 374672
rect 377404 374620 377456 374672
rect 377772 374620 377824 374672
rect 404176 374620 404228 374672
rect 165988 374552 166040 374604
rect 200488 374552 200540 374604
rect 201776 374552 201828 374604
rect 320916 374552 320968 374604
rect 371056 374552 371108 374604
rect 407764 374552 407816 374604
rect 158536 374484 158588 374536
rect 204444 374484 204496 374536
rect 215944 374484 215996 374536
rect 220912 374484 220964 374536
rect 373724 374484 373776 374536
rect 410708 374484 410760 374536
rect 156512 374416 156564 374468
rect 203156 374416 203208 374468
rect 208492 374416 208544 374468
rect 210240 374416 210292 374468
rect 221556 374416 221608 374468
rect 380900 374416 380952 374468
rect 425060 374416 425112 374468
rect 163412 374348 163464 374400
rect 211344 374348 211396 374400
rect 240692 374348 240744 374400
rect 244280 374348 244332 374400
rect 378048 374348 378100 374400
rect 443092 374348 443144 374400
rect 160928 374280 160980 374332
rect 208584 374280 208636 374332
rect 211712 374280 211764 374332
rect 221648 374280 221700 374332
rect 240784 374280 240836 374332
rect 247592 374280 247644 374332
rect 367008 374280 367060 374332
rect 436008 374280 436060 374332
rect 146208 374212 146260 374264
rect 207480 374212 207532 374264
rect 208400 374212 208452 374264
rect 218060 374212 218112 374264
rect 219348 374212 219400 374264
rect 265256 374212 265308 374264
rect 369676 374212 369728 374264
rect 438492 374212 438544 374264
rect 143540 374144 143592 374196
rect 205916 374144 205968 374196
rect 217600 374144 217652 374196
rect 270500 374144 270552 374196
rect 372436 374144 372488 374196
rect 440332 374144 440384 374196
rect 56968 374076 57020 374128
rect 105452 374076 105504 374128
rect 148968 374076 149020 374128
rect 197084 374076 197136 374128
rect 199476 374076 199528 374128
rect 283012 374076 283064 374128
rect 364800 374076 364852 374128
rect 433616 374076 433668 374128
rect 54484 374008 54536 374060
rect 116032 374008 116084 374060
rect 140964 374008 141016 374060
rect 203248 374008 203300 374060
rect 209964 374008 210016 374060
rect 211712 374008 211764 374060
rect 218060 374008 218112 374060
rect 219072 374008 219124 374060
rect 240692 374008 240744 374060
rect 240876 374008 240928 374060
rect 244740 374008 244792 374060
rect 250628 374008 250680 374060
rect 253480 374008 253532 374060
rect 364156 374008 364208 374060
rect 451004 374008 451056 374060
rect 44640 373940 44692 373992
rect 217048 373940 217100 373992
rect 377956 373940 378008 373992
rect 421012 373940 421064 373992
rect 47400 373872 47452 373924
rect 216864 373872 216916 373924
rect 376484 373872 376536 373924
rect 423036 373872 423088 373924
rect 47768 373804 47820 373856
rect 96068 373804 96120 373856
rect 139216 373804 139268 373856
rect 200396 373804 200448 373856
rect 215392 373804 215444 373856
rect 219348 373804 219400 373856
rect 372620 373804 372672 373856
rect 373724 373804 373776 373856
rect 426900 373804 426952 373856
rect 57336 373736 57388 373788
rect 118332 373736 118384 373788
rect 136456 373736 136508 373788
rect 200304 373736 200356 373788
rect 361396 373736 361448 373788
rect 416044 373736 416096 373788
rect 43444 373668 43496 373720
rect 103520 373668 103572 373720
rect 133696 373668 133748 373720
rect 199292 373668 199344 373720
rect 371792 373668 371844 373720
rect 430580 373668 430632 373720
rect 51540 373600 51592 373652
rect 113548 373600 113600 373652
rect 131028 373600 131080 373652
rect 199108 373600 199160 373652
rect 204260 373600 204312 373652
rect 219256 373600 219308 373652
rect 377312 373600 377364 373652
rect 455420 373600 455472 373652
rect 46204 373532 46256 373584
rect 107844 373532 107896 373584
rect 124128 373532 124180 373584
rect 197820 373532 197872 373584
rect 362868 373532 362920 373584
rect 445852 373532 445904 373584
rect 58440 373464 58492 373516
rect 125692 373464 125744 373516
rect 128912 373464 128964 373516
rect 205824 373464 205876 373516
rect 209688 373464 209740 373516
rect 214196 373464 214248 373516
rect 215300 373464 215352 373516
rect 263692 373464 263744 373516
rect 358728 373464 358780 373516
rect 447692 373464 447744 373516
rect 48780 373396 48832 373448
rect 110420 373396 110472 373448
rect 121368 373396 121420 373448
rect 200580 373396 200632 373448
rect 367560 373396 367612 373448
rect 458180 373396 458232 373448
rect 50160 373328 50212 373380
rect 98276 373328 98328 373380
rect 99380 373328 99432 373380
rect 204260 373328 204312 373380
rect 262772 373328 262824 373380
rect 269212 373328 269264 373380
rect 359464 373328 359516 373380
rect 452844 373328 452896 373380
rect 46296 373260 46348 373312
rect 93676 373260 93728 373312
rect 95056 373260 95108 373312
rect 213460 373260 213512 373312
rect 219808 373260 219860 373312
rect 220728 373260 220780 373312
rect 364064 373260 364116 373312
rect 485780 373260 485832 373312
rect 57060 373192 57112 373244
rect 100852 373192 100904 373244
rect 151728 373192 151780 373244
rect 197728 373192 197780 373244
rect 213920 373192 213972 373244
rect 261300 373192 261352 373244
rect 367652 373192 367704 373244
rect 376760 373192 376812 373244
rect 48872 373124 48924 373176
rect 88340 373124 88392 373176
rect 154120 373124 154172 373176
rect 198372 373124 198424 373176
rect 207204 373124 207256 373176
rect 213552 373124 213604 373176
rect 242900 373124 242952 373176
rect 55772 373056 55824 373108
rect 90180 373056 90232 373108
rect 214104 373056 214156 373108
rect 217784 373056 217836 373108
rect 220728 373056 220780 373108
rect 253940 373056 253992 373108
rect 212908 372988 212960 373040
rect 255412 372988 255464 373040
rect 212632 372920 212684 372972
rect 256700 372920 256752 372972
rect 214012 372852 214064 372904
rect 217048 372784 217100 372836
rect 217692 372784 217744 372836
rect 217784 372784 217836 372836
rect 224132 372784 224184 372836
rect 224316 372852 224368 372904
rect 259644 372852 259696 372904
rect 259460 372784 259512 372836
rect 210148 372716 210200 372768
rect 210332 372716 210384 372768
rect 212540 372716 212592 372768
rect 258080 372716 258132 372768
rect 203064 372648 203116 372700
rect 216312 372648 216364 372700
rect 51632 372580 51684 372632
rect 54392 372580 54444 372632
rect 56968 372580 57020 372632
rect 58532 372580 58584 372632
rect 95976 372580 96028 372632
rect 212908 372580 212960 372632
rect 215300 372580 215352 372632
rect 215668 372580 215720 372632
rect 219256 372648 219308 372700
rect 236092 372648 236144 372700
rect 369676 372648 369728 372700
rect 373724 372648 373776 372700
rect 376760 372648 376812 372700
rect 378048 372648 378100 372700
rect 408500 372648 408552 372700
rect 236000 372580 236052 372632
rect 372528 372580 372580 372632
rect 374000 372580 374052 372632
rect 375196 372580 375248 372632
rect 379152 372580 379204 372632
rect 379336 372580 379388 372632
rect 426440 372580 426492 372632
rect 89352 372512 89404 372564
rect 209872 372512 209924 372564
rect 210332 372512 210384 372564
rect 211712 372512 211764 372564
rect 213736 372512 213788 372564
rect 214472 372512 214524 372564
rect 219532 372512 219584 372564
rect 273260 372512 273312 372564
rect 305000 372512 305052 372564
rect 313280 372512 313332 372564
rect 369860 372512 369912 372564
rect 437480 372512 437532 372564
rect 92388 372444 92440 372496
rect 90088 372376 90140 372428
rect 77208 372308 77260 372360
rect 99380 372308 99432 372360
rect 304264 372444 304316 372496
rect 310520 372444 310572 372496
rect 375196 372444 375248 372496
rect 433340 372444 433392 372496
rect 220728 372376 220780 372428
rect 248420 372376 248472 372428
rect 211160 372308 211212 372360
rect 221004 372308 221056 372360
rect 221924 372308 221976 372360
rect 209780 372240 209832 372292
rect 220084 372240 220136 372292
rect 221556 372172 221608 372224
rect 240876 372172 240928 372224
rect 86592 372104 86644 372156
rect 210148 372104 210200 372156
rect 215760 372104 215812 372156
rect 245660 372104 245712 372156
rect 210332 372036 210384 372088
rect 219532 372036 219584 372088
rect 220728 372036 220780 372088
rect 47676 371968 47728 372020
rect 78496 371968 78548 372020
rect 213460 371968 213512 372020
rect 219624 371968 219676 372020
rect 251180 372036 251232 372088
rect 368388 372036 368440 372088
rect 376760 372036 376812 372088
rect 221648 371968 221700 372020
rect 240784 371968 240836 372020
rect 357256 371968 357308 372020
rect 379520 371968 379572 372020
rect 379980 371968 380032 372020
rect 396080 371968 396132 372020
rect 44732 371900 44784 371952
rect 48872 371900 48924 371952
rect 108856 371900 108908 371952
rect 204168 371900 204220 371952
rect 217048 371900 217100 371952
rect 262864 371900 262916 371952
rect 360752 371900 360804 371952
rect 376484 371900 376536 371952
rect 379428 371900 379480 371952
rect 404360 371900 404412 371952
rect 47584 371832 47636 371884
rect 79968 371832 80020 371884
rect 85488 371832 85540 371884
rect 106188 371832 106240 371884
rect 114008 371832 114060 371884
rect 214472 371832 214524 371884
rect 215024 371832 215076 371884
rect 88064 371764 88116 371816
rect 211712 371764 211764 371816
rect 93584 371696 93636 371748
rect 220912 371832 220964 371884
rect 250628 371832 250680 371884
rect 275376 371832 275428 371884
rect 356980 371832 357032 371884
rect 375196 371832 375248 371884
rect 400220 371832 400272 371884
rect 517888 371832 517940 371884
rect 580448 371832 580500 371884
rect 222108 371764 222160 371816
rect 241520 371764 241572 371816
rect 92204 371628 92256 371680
rect 211252 371628 211304 371680
rect 213460 371628 213512 371680
rect 215300 371560 215352 371612
rect 215576 371560 215628 371612
rect 240416 371560 240468 371612
rect 241428 371560 241480 371612
rect 276296 371764 276348 371816
rect 357256 371764 357308 371816
rect 372988 371764 373040 371816
rect 398840 371764 398892 371816
rect 273260 371696 273312 371748
rect 305000 371696 305052 371748
rect 371056 371696 371108 371748
rect 397460 371696 397512 371748
rect 278688 371628 278740 371680
rect 357440 371628 357492 371680
rect 379520 371628 379572 371680
rect 379888 371628 379940 371680
rect 409880 371628 409932 371680
rect 371148 371560 371200 371612
rect 48872 371492 48924 371544
rect 81900 371492 81952 371544
rect 82452 371492 82504 371544
rect 85120 371492 85172 371544
rect 210240 371492 210292 371544
rect 215116 371492 215168 371544
rect 221924 371492 221976 371544
rect 223120 371492 223172 371544
rect 237380 371492 237432 371544
rect 238116 371492 238168 371544
rect 371056 371492 371108 371544
rect 376576 371560 376628 371612
rect 380992 371560 381044 371612
rect 411260 371560 411312 371612
rect 401600 371492 401652 371544
rect 79968 371424 80020 371476
rect 209596 371424 209648 371476
rect 239312 371424 239364 371476
rect 372988 371424 373040 371476
rect 376484 371424 376536 371476
rect 407120 371424 407172 371476
rect 78496 371356 78548 371408
rect 208216 371356 208268 371408
rect 237380 371356 237432 371408
rect 241428 371356 241480 371408
rect 375196 371356 375248 371408
rect 376760 371356 376812 371408
rect 377956 371356 378008 371408
rect 411260 371356 411312 371408
rect 439872 371356 439924 371408
rect 516600 371356 516652 371408
rect 44824 371220 44876 371272
rect 46296 371220 46348 371272
rect 80520 371288 80572 371340
rect 215300 371288 215352 371340
rect 219900 371288 219952 371340
rect 220084 371288 220136 371340
rect 249800 371288 249852 371340
rect 342904 371288 342956 371340
rect 343456 371288 343508 371340
rect 363052 371288 363104 371340
rect 503536 371288 503588 371340
rect 517888 371288 517940 371340
rect 82452 371220 82504 371272
rect 220820 371220 220872 371272
rect 222108 371220 222160 371272
rect 223120 371220 223172 371272
rect 251180 371220 251232 371272
rect 343088 371220 343140 371272
rect 360200 371220 360252 371272
rect 503168 371220 503220 371272
rect 517796 371220 517848 371272
rect 580264 371220 580316 371272
rect 43352 371152 43404 371204
rect 183192 371152 183244 371204
rect 201040 371152 201092 371204
rect 201500 371152 201552 371204
rect 317420 371152 317472 371204
rect 375104 371152 375156 371204
rect 376576 371152 376628 371204
rect 376760 371152 376812 371204
rect 402980 371152 403032 371204
rect 54576 371084 54628 371136
rect 182824 371084 182876 371136
rect 198832 371084 198884 371136
rect 302240 371084 302292 371136
rect 357992 371084 358044 371136
rect 473360 371084 473412 371136
rect 197360 371016 197412 371068
rect 295340 371016 295392 371068
rect 357164 371016 357216 371068
rect 465080 371016 465132 371068
rect 102784 370948 102836 371000
rect 215484 370948 215536 371000
rect 217508 370948 217560 371000
rect 307760 370948 307812 371000
rect 366180 370948 366232 371000
rect 467840 370948 467892 371000
rect 198924 370880 198976 370932
rect 300860 370880 300912 370932
rect 368940 370880 368992 370932
rect 470600 370880 470652 370932
rect 197452 370812 197504 370864
rect 292580 370812 292632 370864
rect 361488 370812 361540 370864
rect 462320 370812 462372 370864
rect 196716 370744 196768 370796
rect 289820 370744 289872 370796
rect 364892 370744 364944 370796
rect 460940 370744 460992 370796
rect 196808 370676 196860 370728
rect 287244 370676 287296 370728
rect 359556 370676 359608 370728
rect 413192 370676 413244 370728
rect 196624 370608 196676 370660
rect 285680 370608 285732 370660
rect 373816 370608 373868 370660
rect 375932 370608 375984 370660
rect 376760 370608 376812 370660
rect 379244 370608 379296 370660
rect 415400 370608 415452 370660
rect 199384 370540 199436 370592
rect 280160 370540 280212 370592
rect 369032 370540 369084 370592
rect 374000 370540 374052 370592
rect 422300 370540 422352 370592
rect 102048 370472 102100 370524
rect 209504 370472 209556 370524
rect 213920 370472 213972 370524
rect 217416 370472 217468 370524
rect 298100 370472 298152 370524
rect 360016 370472 360068 370524
rect 518992 370472 519044 370524
rect 196992 370404 197044 370456
rect 277768 370404 277820 370456
rect 376668 370404 376720 370456
rect 379796 370404 379848 370456
rect 414020 370404 414072 370456
rect 198740 370336 198792 370388
rect 273260 370336 273312 370388
rect 376576 370336 376628 370388
rect 396080 370336 396132 370388
rect 77024 370268 77076 370320
rect 203064 370268 203116 370320
rect 212908 370268 212960 370320
rect 213460 370268 213512 370320
rect 215668 370268 215720 370320
rect 217140 370268 217192 370320
rect 362132 370268 362184 370320
rect 483020 370268 483072 370320
rect 359464 369860 359516 369912
rect 360016 369860 360068 369912
rect 83832 369792 83884 369844
rect 207204 369792 207256 369844
rect 216404 369792 216456 369844
rect 247040 369792 247092 369844
rect 373908 369792 373960 369844
rect 376944 369792 376996 369844
rect 378048 369792 378100 369844
rect 202880 369724 202932 369776
rect 325884 369724 325936 369776
rect 374460 369724 374512 369776
rect 477500 369724 477552 369776
rect 202972 369656 203024 369708
rect 322940 369656 322992 369708
rect 356888 369656 356940 369708
rect 418160 369656 418212 369708
rect 205364 369588 205416 369640
rect 264980 369588 265032 369640
rect 373172 369588 373224 369640
rect 427820 369588 427872 369640
rect 54576 369520 54628 369572
rect 56508 369520 56560 369572
rect 211528 369520 211580 369572
rect 267740 369520 267792 369572
rect 370412 369520 370464 369572
rect 202420 369452 202472 369504
rect 263600 369452 263652 369504
rect 201132 369384 201184 369436
rect 260840 369384 260892 369436
rect 378600 369520 378652 369572
rect 425060 369520 425112 369572
rect 378048 369452 378100 369504
rect 423680 369452 423732 369504
rect 374552 369384 374604 369436
rect 416780 369384 416832 369436
rect 203892 369316 203944 369368
rect 258172 369316 258224 369368
rect 371700 369316 371752 369368
rect 375932 369316 375984 369368
rect 418252 369316 418304 369368
rect 100116 369248 100168 369300
rect 214012 369248 214064 369300
rect 214380 369248 214432 369300
rect 219164 369248 219216 369300
rect 273352 369248 273404 369300
rect 365628 369248 365680 369300
rect 377128 369248 377180 369300
rect 419540 369248 419592 369300
rect 99288 369180 99340 369232
rect 211620 369180 211672 369232
rect 212540 369180 212592 369232
rect 366272 369180 366324 369232
rect 371792 369180 371844 369232
rect 420920 369180 420972 369232
rect 97724 369112 97776 369164
rect 210240 369112 210292 369164
rect 212632 369112 212684 369164
rect 359556 369112 359608 369164
rect 360108 369112 360160 369164
rect 519084 369112 519136 369164
rect 206284 369044 206336 369096
rect 249892 369044 249944 369096
rect 368296 369044 368348 369096
rect 376668 369044 376720 369096
rect 418344 369044 418396 369096
rect 106188 368976 106240 369028
rect 208400 368976 208452 369028
rect 213092 368976 213144 369028
rect 276020 368976 276072 369028
rect 361304 368976 361356 369028
rect 378692 368976 378744 369028
rect 405740 368976 405792 369028
rect 208032 368908 208084 368960
rect 252560 368908 252612 368960
rect 370320 368908 370372 368960
rect 480260 368908 480312 368960
rect 208860 368840 208912 368892
rect 255320 368840 255372 368892
rect 101036 368772 101088 368824
rect 214104 368772 214156 368824
rect 214472 368772 214524 368824
rect 54484 368636 54536 368688
rect 55864 368636 55916 368688
rect 215300 368432 215352 368484
rect 216588 368432 216640 368484
rect 219716 368432 219768 368484
rect 266360 368432 266412 368484
rect 365536 368092 365588 368144
rect 379336 368092 379388 368144
rect 412640 368092 412692 368144
rect 357900 368024 357952 368076
rect 368388 368024 368440 368076
rect 427912 368024 427964 368076
rect 357072 367956 357124 368008
rect 375104 367956 375156 368008
rect 436100 367956 436152 368008
rect 362776 367888 362828 367940
rect 370412 367888 370464 367940
rect 431960 367888 432012 367940
rect 364248 367820 364300 367872
rect 368296 367820 368348 367872
rect 434720 367820 434772 367872
rect 107568 367752 107620 367804
rect 215300 367752 215352 367804
rect 359004 367752 359056 367804
rect 359924 367752 359976 367804
rect 519176 367752 519228 367804
rect 199384 366324 199436 366376
rect 199752 366324 199804 366376
rect 359004 366324 359056 366376
rect 201040 364284 201092 364336
rect 343088 364284 343140 364336
rect 199476 362176 199528 362228
rect 359096 362176 359148 362228
rect 359464 362176 359516 362228
rect 208400 360136 208452 360188
rect 209688 360136 209740 360188
rect 359188 360136 359240 360188
rect 199752 359456 199804 359508
rect 208400 359456 208452 359508
rect 359280 359456 359332 359508
rect 359832 359456 359884 359508
rect 519268 359456 519320 359508
rect 3332 358708 3384 358760
rect 18604 358708 18656 358760
rect 359464 358096 359516 358148
rect 519360 358096 519412 358148
rect 199568 358028 199620 358080
rect 359280 358028 359332 358080
rect 182824 356668 182876 356720
rect 202880 356668 202932 356720
rect 342904 356668 342956 356720
rect 191380 355988 191432 356040
rect 206928 356056 206980 356108
rect 215944 356056 215996 356108
rect 357348 355988 357400 356040
rect 362960 355988 363012 356040
rect 179788 355920 179840 355972
rect 195888 355920 195940 355972
rect 500868 355444 500920 355496
rect 517612 355444 517664 355496
rect 340052 355376 340104 355428
rect 356612 355376 356664 355428
rect 498844 355376 498896 355428
rect 517704 355376 517756 355428
rect 351736 355308 351788 355360
rect 358084 355308 358136 355360
rect 195888 355172 195940 355224
rect 197360 355172 197412 355224
rect 356612 354968 356664 355020
rect 356888 354968 356940 355020
rect 338120 354764 338172 354816
rect 357348 354764 357400 354816
rect 510896 354764 510948 354816
rect 517520 354764 517572 354816
rect 178592 354696 178644 354748
rect 197728 354696 197780 354748
rect 201960 354696 202012 354748
rect 199660 353948 199712 354000
rect 359556 353948 359608 354000
rect 373172 353948 373224 354000
rect 381084 353948 381136 354000
rect 217876 353404 217928 353456
rect 220820 353404 220872 353456
rect 55864 353336 55916 353388
rect 60740 353336 60792 353388
rect 218612 353336 218664 353388
rect 220912 353336 220964 353388
rect 378600 353336 378652 353388
rect 380900 353336 380952 353388
rect 58624 353268 58676 353320
rect 62120 353268 62172 353320
rect 219164 353268 219216 353320
rect 221004 353268 221056 353320
rect 359188 353268 359240 353320
rect 359556 353268 359608 353320
rect 379244 353268 379296 353320
rect 380992 353268 381044 353320
rect 54392 352520 54444 352572
rect 59452 352520 59504 352572
rect 56876 351908 56928 351960
rect 59360 351908 59412 351960
rect 58532 350548 58584 350600
rect 59728 350548 59780 350600
rect 47860 298052 47912 298104
rect 57520 298052 57572 298104
rect 520188 284316 520240 284368
rect 580264 284316 580316 284368
rect 519084 282888 519136 282940
rect 580356 282888 580408 282940
rect 200948 280100 201000 280152
rect 216680 280100 216732 280152
rect 55680 278672 55732 278724
rect 58716 278672 58768 278724
rect 206744 278672 206796 278724
rect 216680 278672 216732 278724
rect 361212 278672 361264 278724
rect 376760 278672 376812 278724
rect 215944 278264 215996 278316
rect 216956 278264 217008 278316
rect 358084 277992 358136 278044
rect 376852 277992 376904 278044
rect 378600 270444 378652 270496
rect 379612 270444 379664 270496
rect 51448 269764 51500 269816
rect 54484 269764 54536 269816
rect 55220 269764 55272 269816
rect 373172 269764 373224 269816
rect 374460 269764 374512 269816
rect 45192 269696 45244 269748
rect 148508 269696 148560 269748
rect 46204 269628 46256 269680
rect 59820 269628 59872 269680
rect 60096 269628 60148 269680
rect 51540 269560 51592 269612
rect 51724 269560 51776 269612
rect 52920 269560 52972 269612
rect 110972 269560 111024 269612
rect 43536 269492 43588 269544
rect 133420 269492 133472 269544
rect 379612 269492 379664 269544
rect 425244 269492 425296 269544
rect 44916 269424 44968 269476
rect 135904 269424 135956 269476
rect 363972 269424 364024 269476
rect 416044 269424 416096 269476
rect 45008 269356 45060 269408
rect 138480 269356 138532 269408
rect 374460 269356 374512 269408
rect 433340 269356 433392 269408
rect 45100 269288 45152 269340
rect 140872 269288 140924 269340
rect 210792 269288 210844 269340
rect 250720 269288 250772 269340
rect 371700 269288 371752 269340
rect 372528 269288 372580 269340
rect 434352 269288 434404 269340
rect 45376 269220 45428 269272
rect 143540 269220 143592 269272
rect 205272 269220 205324 269272
rect 283472 269220 283524 269272
rect 370964 269220 371016 269272
rect 436008 269220 436060 269272
rect 45284 269152 45336 269204
rect 145932 269152 145984 269204
rect 206652 269152 206704 269204
rect 288256 269152 288308 269204
rect 372528 269152 372580 269204
rect 374000 269152 374052 269204
rect 374460 269152 374512 269204
rect 375012 269152 375064 269204
rect 468484 269152 468536 269204
rect 45468 269016 45520 269068
rect 50344 269016 50396 269068
rect 51724 269016 51776 269068
rect 91284 269084 91336 269136
rect 207940 269084 207992 269136
rect 291016 269084 291068 269136
rect 365352 269084 365404 269136
rect 470968 269084 471020 269136
rect 196624 269016 196676 269068
rect 197176 269016 197228 269068
rect 213552 269016 213604 269068
rect 215392 269016 215444 269068
rect 373080 269016 373132 269068
rect 373724 269016 373776 269068
rect 379520 269016 379572 269068
rect 379796 269016 379848 269068
rect 62120 268948 62172 269000
rect 211620 268948 211672 269000
rect 216956 268948 217008 269000
rect 46480 268880 46532 268932
rect 54668 268880 54720 268932
rect 213460 268880 213512 268932
rect 236000 268880 236052 268932
rect 212172 268812 212224 268864
rect 298468 268812 298520 268864
rect 374460 268812 374512 268864
rect 422852 268812 422904 268864
rect 209320 268744 209372 268796
rect 295892 268744 295944 268796
rect 368112 268744 368164 268796
rect 430948 268744 431000 268796
rect 60096 268676 60148 268728
rect 94504 268676 94556 268728
rect 202328 268676 202380 268728
rect 293408 268676 293460 268728
rect 361028 268676 361080 268728
rect 425980 268676 426032 268728
rect 58532 268608 58584 268660
rect 93584 268608 93636 268660
rect 203800 268608 203852 268660
rect 300860 268608 300912 268660
rect 356796 268608 356848 268660
rect 421012 268608 421064 268660
rect 48044 268540 48096 268592
rect 90732 268540 90784 268592
rect 205180 268540 205232 268592
rect 305920 268540 305972 268592
rect 366916 268540 366968 268592
rect 475844 268540 475896 268592
rect 51908 268472 51960 268524
rect 98460 268472 98512 268524
rect 200764 268472 200816 268524
rect 303436 268472 303488 268524
rect 369584 268472 369636 268524
rect 478420 268472 478472 268524
rect 49056 268404 49108 268456
rect 96068 268404 96120 268456
rect 209504 268404 209556 268456
rect 214472 268404 214524 268456
rect 214932 268404 214984 268456
rect 323308 268404 323360 268456
rect 372160 268404 372212 268456
rect 480904 268404 480956 268456
rect 51540 268336 51592 268388
rect 53748 268336 53800 268388
rect 55220 268336 55272 268388
rect 100760 268336 100812 268388
rect 198004 268336 198056 268388
rect 318432 268336 318484 268388
rect 362684 268336 362736 268388
rect 483388 268336 483440 268388
rect 48136 268200 48188 268252
rect 77116 268200 77168 268252
rect 373724 268200 373776 268252
rect 429752 268200 429804 268252
rect 54208 268132 54260 268184
rect 54484 268132 54536 268184
rect 66260 268132 66312 268184
rect 95884 268132 95936 268184
rect 373172 268132 373224 268184
rect 432236 268132 432288 268184
rect 46388 268064 46440 268116
rect 76012 268064 76064 268116
rect 79324 268064 79376 268116
rect 106372 268064 106424 268116
rect 396724 268064 396776 268116
rect 415400 268064 415452 268116
rect 48964 267996 49016 268048
rect 83096 267996 83148 268048
rect 395344 267996 395396 268048
rect 416964 267996 417016 268048
rect 54300 267928 54352 267980
rect 54668 267928 54720 267980
rect 96988 267928 97040 267980
rect 236000 267928 236052 267980
rect 247040 267928 247092 267980
rect 373816 267928 373868 267980
rect 374276 267928 374328 267980
rect 402980 267928 403032 267980
rect 58716 267860 58768 267912
rect 59820 267860 59872 267912
rect 102692 267860 102744 267912
rect 106924 267860 106976 267912
rect 119068 267860 119120 267912
rect 215392 267860 215444 267912
rect 243084 267860 243136 267912
rect 379520 267860 379572 267912
rect 414388 267860 414440 267912
rect 54208 267792 54260 267844
rect 99380 267792 99432 267844
rect 112352 267792 112404 267844
rect 197912 267792 197964 267844
rect 201592 267792 201644 267844
rect 217968 267792 218020 267844
rect 258080 267792 258132 267844
rect 427084 267792 427136 267844
rect 434720 267792 434772 267844
rect 51448 267724 51500 267776
rect 51724 267724 51776 267776
rect 98000 267724 98052 267776
rect 111248 267724 111300 267776
rect 196624 267724 196676 267776
rect 214472 267724 214524 267776
rect 261668 267724 261720 267776
rect 425704 267724 425756 267776
rect 428556 267724 428608 267776
rect 43628 267656 43680 267708
rect 128360 267656 128412 267708
rect 158536 267656 158588 267708
rect 205640 267656 205692 267708
rect 247040 267656 247092 267708
rect 255320 267656 255372 267708
rect 372252 267656 372304 267708
rect 460940 267656 460992 267708
rect 42248 267588 42300 267640
rect 125600 267588 125652 267640
rect 150992 267588 151044 267640
rect 198096 267588 198148 267640
rect 209228 267588 209280 267640
rect 280160 267588 280212 267640
rect 369492 267588 369544 267640
rect 452660 267588 452712 267640
rect 43812 267520 43864 267572
rect 120080 267520 120132 267572
rect 203524 267520 203576 267572
rect 267832 267520 267884 267572
rect 370412 267520 370464 267572
rect 373172 267520 373224 267572
rect 376392 267520 376444 267572
rect 458180 267520 458232 267572
rect 42340 267452 42392 267504
rect 50988 267452 51040 267504
rect 55864 267452 55916 267504
rect 129740 267452 129792 267504
rect 163504 267452 163556 267504
rect 197636 267452 197688 267504
rect 200856 267452 200908 267504
rect 264980 267452 265032 267504
rect 368204 267452 368256 267504
rect 449900 267452 449952 267504
rect 53104 267384 53156 267436
rect 117320 267384 117372 267436
rect 155960 267384 156012 267436
rect 201868 267384 201920 267436
rect 202236 267384 202288 267436
rect 263600 267384 263652 267436
rect 374920 267384 374972 267436
rect 455788 267384 455840 267436
rect 53196 267316 53248 267368
rect 115940 267316 115992 267368
rect 160928 267316 160980 267368
rect 207112 267316 207164 267368
rect 214840 267316 214892 267368
rect 273260 267316 273312 267368
rect 49148 267248 49200 267300
rect 52920 267248 52972 267300
rect 53012 267248 53064 267300
rect 113548 267248 113600 267300
rect 218980 267248 219032 267300
rect 276020 267248 276072 267300
rect 343456 267248 343508 267300
rect 360200 267316 360252 267368
rect 363880 267316 363932 267368
rect 443000 267316 443052 267368
rect 52000 267180 52052 267232
rect 107660 267180 107712 267232
rect 216128 267180 216180 267232
rect 270500 267180 270552 267232
rect 278136 267180 278188 267232
rect 357716 267248 357768 267300
rect 362592 267248 362644 267300
rect 440240 267248 440292 267300
rect 356612 267180 356664 267232
rect 357256 267180 357308 267232
rect 370872 267180 370924 267232
rect 447140 267180 447192 267232
rect 503168 267180 503220 267232
rect 517796 267180 517848 267232
rect 51816 267112 51868 267164
rect 104900 267112 104952 267164
rect 205088 267112 205140 267164
rect 258264 267112 258316 267164
rect 279148 267112 279200 267164
rect 358820 267112 358872 267164
rect 372344 267112 372396 267164
rect 445760 267112 445812 267164
rect 52092 267044 52144 267096
rect 103520 267044 103572 267096
rect 198280 267044 198332 267096
rect 202880 267044 202932 267096
rect 210884 267044 210936 267096
rect 260840 267044 260892 267096
rect 277032 267044 277084 267096
rect 356612 267044 356664 267096
rect 366824 267044 366876 267096
rect 437480 267044 437532 267096
rect 503536 267044 503588 267096
rect 517888 267044 517940 267096
rect 50252 266976 50304 267028
rect 100760 266976 100812 267028
rect 183284 266976 183336 267028
rect 200120 266976 200172 267028
rect 201040 266976 201092 267028
rect 215024 266976 215076 267028
rect 273260 266976 273312 267028
rect 275928 266976 275980 267028
rect 356980 266976 357032 267028
rect 365444 266976 365496 267028
rect 433340 266976 433392 267028
rect 440056 266976 440108 267028
rect 516600 266976 516652 267028
rect 54760 266908 54812 266960
rect 88340 266908 88392 266960
rect 206560 266908 206612 266960
rect 255320 266908 255372 266960
rect 358452 266908 358504 266960
rect 418160 266908 418212 266960
rect 48044 266840 48096 266892
rect 78680 266840 78732 266892
rect 207848 266840 207900 266892
rect 252560 266840 252612 266892
rect 376208 266840 376260 266892
rect 412916 266840 412968 266892
rect 47768 266772 47820 266824
rect 77300 266772 77352 266824
rect 216220 266772 216272 266824
rect 247040 266772 247092 266824
rect 373632 266772 373684 266824
rect 409880 266772 409932 266824
rect 213368 266704 213420 266756
rect 285680 266704 285732 266756
rect 47676 266500 47728 266552
rect 48044 266500 48096 266552
rect 50344 266364 50396 266416
rect 50988 266364 51040 266416
rect 80060 266364 80112 266416
rect 104900 266364 104952 266416
rect 183468 266364 183520 266416
rect 197452 266364 197504 266416
rect 198280 266364 198332 266416
rect 343456 266364 343508 266416
rect 357072 266432 357124 266484
rect 363052 266432 363104 266484
rect 356796 266364 356848 266416
rect 356980 266364 357032 266416
rect 421564 266364 421616 266416
rect 437480 266364 437532 266416
rect 517796 266364 517848 266416
rect 517980 266364 518032 266416
rect 55772 266296 55824 266348
rect 56876 266296 56928 266348
rect 57980 266296 58032 266348
rect 58624 266296 58676 266348
rect 92388 266296 92440 266348
rect 109960 266296 110012 266348
rect 196808 266296 196860 266348
rect 216220 266296 216272 266348
rect 262220 266296 262272 266348
rect 379980 266296 380032 266348
rect 396080 266296 396132 266348
rect 54576 266228 54628 266280
rect 55864 266228 55916 266280
rect 117320 266228 117372 266280
rect 213736 266228 213788 266280
rect 247040 266228 247092 266280
rect 379244 266228 379296 266280
rect 411260 266228 411312 266280
rect 51908 266160 51960 266212
rect 57980 266160 58032 266212
rect 216956 266160 217008 266212
rect 219164 266160 219216 266212
rect 251272 266160 251324 266212
rect 373908 266160 373960 266212
rect 376484 266160 376536 266212
rect 407120 266160 407172 266212
rect 62212 266092 62264 266144
rect 92480 266092 92532 266144
rect 219256 266092 219308 266144
rect 219624 266092 219676 266144
rect 251180 266092 251232 266144
rect 378048 266092 378100 266144
rect 408500 266092 408552 266144
rect 54484 266024 54536 266076
rect 84200 266024 84252 266076
rect 215668 266024 215720 266076
rect 245660 266024 245712 266076
rect 379888 266024 379940 266076
rect 409880 266024 409932 266076
rect 57980 265956 58032 266008
rect 89720 265956 89772 266008
rect 196716 265956 196768 266008
rect 197544 265956 197596 266008
rect 215116 265956 215168 266008
rect 216128 265956 216180 266008
rect 217968 265956 218020 266008
rect 219900 265956 219952 266008
rect 249800 265956 249852 266008
rect 375196 265956 375248 266008
rect 400220 265956 400272 266008
rect 54576 265888 54628 265940
rect 85580 265888 85632 265940
rect 219164 265888 219216 265940
rect 219532 265888 219584 265940
rect 248512 265888 248564 265940
rect 370228 265888 370280 265940
rect 372988 265888 373040 265940
rect 398840 265888 398892 265940
rect 50436 265684 50488 265736
rect 52000 265820 52052 265872
rect 85396 265820 85448 265872
rect 218612 265820 218664 265872
rect 219900 265820 219952 265872
rect 252560 265820 252612 265872
rect 379704 265820 379756 265872
rect 404360 265820 404412 265872
rect 55864 265752 55916 265804
rect 88340 265752 88392 265804
rect 217140 265752 217192 265804
rect 218980 265752 219032 265804
rect 263600 265752 263652 265804
rect 371056 265752 371108 265804
rect 372436 265752 372488 265804
rect 398196 265752 398248 265804
rect 53104 265684 53156 265736
rect 86960 265684 87012 265736
rect 88248 265684 88300 265736
rect 113732 265684 113784 265736
rect 215484 265684 215536 265736
rect 216220 265684 216272 265736
rect 219348 265684 219400 265736
rect 219624 265684 219676 265736
rect 265164 265684 265216 265736
rect 376576 265684 376628 265736
rect 403164 265684 403216 265736
rect 59728 265616 59780 265668
rect 107660 265616 107712 265668
rect 114376 265616 114428 265668
rect 196716 265616 196768 265668
rect 216588 265616 216640 265668
rect 218612 265616 218664 265668
rect 266360 265616 266412 265668
rect 371148 265616 371200 265668
rect 372344 265616 372396 265668
rect 401692 265616 401744 265668
rect 216128 265548 216180 265600
rect 244280 265548 244332 265600
rect 377956 265548 378008 265600
rect 411352 265548 411404 265600
rect 375288 265412 375340 265464
rect 376576 265412 376628 265464
rect 376392 265276 376444 265328
rect 374092 265208 374144 265260
rect 379980 265208 380032 265260
rect 375932 265140 375984 265192
rect 213644 265072 213696 265124
rect 215668 265072 215720 265124
rect 214380 265004 214432 265056
rect 230388 265004 230440 265056
rect 378508 265004 378560 265056
rect 379704 265004 379756 265056
rect 47952 264936 48004 264988
rect 214288 264936 214340 264988
rect 215760 264936 215812 264988
rect 233148 264936 233200 264988
rect 376852 264936 376904 264988
rect 378048 264936 378100 264988
rect 378600 264936 378652 264988
rect 379888 264936 379940 264988
rect 390560 265004 390612 265056
rect 391940 264936 391992 264988
rect 51632 264868 51684 264920
rect 88248 264868 88300 264920
rect 212172 264868 212224 264920
rect 273168 264868 273220 264920
rect 388444 264868 388496 264920
rect 420920 264868 420972 264920
rect 43720 264800 43772 264852
rect 59728 264800 59780 264852
rect 211712 264800 211764 264852
rect 270500 264800 270552 264852
rect 389180 264800 389232 264852
rect 419540 264800 419592 264852
rect 49240 264732 49292 264784
rect 62212 264732 62264 264784
rect 219808 264732 219860 264784
rect 253940 264732 253992 264784
rect 378692 264732 378744 264784
rect 405740 264732 405792 264784
rect 48228 264664 48280 264716
rect 57980 264664 58032 264716
rect 230388 264664 230440 264716
rect 259552 264664 259604 264716
rect 390560 264664 390612 264716
rect 418252 264664 418304 264716
rect 46756 264596 46808 264648
rect 54484 264596 54536 264648
rect 233148 264596 233200 264648
rect 259460 264596 259512 264648
rect 391940 264596 391992 264648
rect 418160 264596 418212 264648
rect 46664 264528 46716 264580
rect 53104 264528 53156 264580
rect 215116 264528 215168 264580
rect 219072 264528 219124 264580
rect 244372 264528 244424 264580
rect 46572 264460 46624 264512
rect 54576 264460 54628 264512
rect 210240 264256 210292 264308
rect 217140 264256 217192 264308
rect 256700 264256 256752 264308
rect 57796 264188 57848 264240
rect 80060 264188 80112 264240
rect 213552 264188 213604 264240
rect 269120 264188 269172 264240
rect 379336 264188 379388 264240
rect 413008 264188 413060 264240
rect 210332 263644 210384 263696
rect 213552 263644 213604 263696
rect 211712 263576 211764 263628
rect 212080 263576 212132 263628
rect 376484 263576 376536 263628
rect 378692 263576 378744 263628
rect 379336 263576 379388 263628
rect 379888 263576 379940 263628
rect 42432 263508 42484 263560
rect 57244 263508 57296 263560
rect 57796 263508 57848 263560
rect 375104 263508 375156 263560
rect 436100 263508 436152 263560
rect 214380 262964 214432 263016
rect 378968 262828 379020 262880
rect 426440 262828 426492 262880
rect 214472 262692 214524 262744
rect 369676 262148 369728 262200
rect 378968 262148 379020 262200
rect 220820 251132 220872 251184
rect 221372 251132 221424 251184
rect 266452 251132 266504 251184
rect 369768 251132 369820 251184
rect 370412 251132 370464 251184
rect 374552 251132 374604 251184
rect 395344 251132 395396 251184
rect 197360 251064 197412 251116
rect 197636 251064 197688 251116
rect 368388 251064 368440 251116
rect 370964 251064 371016 251116
rect 379152 251064 379204 251116
rect 379428 251064 379480 251116
rect 396724 251064 396776 251116
rect 368296 250996 368348 251048
rect 370872 250996 370924 251048
rect 500040 250656 500092 250708
rect 517612 250656 517664 250708
rect 204168 250588 204220 250640
rect 58716 250520 58768 250572
rect 79324 250520 79376 250572
rect 85856 250520 85908 250572
rect 106924 250520 106976 250572
rect 179788 250520 179840 250572
rect 197636 250520 197688 250572
rect 58624 250452 58676 250504
rect 106280 250452 106332 250504
rect 179328 250452 179380 250504
rect 197544 250452 197596 250504
rect 203524 250452 203576 250504
rect 215944 250452 215996 250504
rect 340052 250588 340104 250640
rect 356888 250588 356940 250640
rect 370412 250588 370464 250640
rect 421564 250588 421616 250640
rect 219072 250520 219124 250572
rect 236000 250520 236052 250572
rect 338488 250520 338540 250572
rect 357624 250520 357676 250572
rect 370964 250520 371016 250572
rect 425704 250520 425756 250572
rect 499028 250520 499080 250572
rect 517704 250520 517756 250572
rect 219532 250452 219584 250504
rect 267740 250452 267792 250504
rect 351736 250452 351788 250504
rect 358084 250452 358136 250504
rect 370872 250452 370924 250504
rect 427084 250452 427136 250504
rect 517612 250248 517664 250300
rect 518072 250248 518124 250300
rect 510896 249908 510948 249960
rect 517520 249908 517572 249960
rect 190920 249772 190972 249824
rect 203524 249772 203576 249824
rect 218520 249772 218572 249824
rect 221372 249772 221424 249824
rect 43904 249704 43956 249756
rect 58716 249704 58768 249756
rect 56968 248956 57020 249008
rect 62120 248956 62172 249008
rect 3056 202784 3108 202836
rect 42064 202784 42116 202836
rect 520188 182180 520240 182232
rect 580264 182180 580316 182232
rect 519544 182112 519596 182164
rect 580356 182112 580408 182164
rect 368020 175176 368072 175228
rect 376852 175176 376904 175228
rect 43996 173816 44048 173868
rect 57796 173816 57848 173868
rect 203524 173816 203576 173868
rect 204168 173816 204220 173868
rect 216680 173816 216732 173868
rect 366732 173816 366784 173868
rect 377128 173816 377180 173868
rect 206468 173748 206520 173800
rect 217048 173748 217100 173800
rect 198004 173136 198056 173188
rect 204168 173136 204220 173188
rect 358084 173136 358136 173188
rect 376852 173136 376904 173188
rect 54392 165520 54444 165572
rect 56508 165520 56560 165572
rect 50620 164636 50672 164688
rect 96068 164636 96120 164688
rect 55680 164568 55732 164620
rect 56508 164568 56560 164620
rect 115756 164568 115808 164620
rect 59176 164500 59228 164552
rect 140872 164500 140924 164552
rect 55956 164432 56008 164484
rect 138480 164432 138532 164484
rect 42524 164364 42576 164416
rect 143540 164364 143592 164416
rect 373448 164364 373500 164416
rect 425980 164364 426032 164416
rect 39856 164296 39908 164348
rect 163320 164296 163372 164348
rect 210700 164296 210752 164348
rect 261024 164296 261076 164348
rect 369400 164296 369452 164348
rect 451004 164296 451056 164348
rect 41328 164228 41380 164280
rect 165896 164228 165948 164280
rect 203616 164228 203668 164280
rect 288256 164228 288308 164280
rect 365260 164228 365312 164280
rect 480904 164228 480956 164280
rect 357532 164160 357584 164212
rect 360200 164160 360252 164212
rect 374920 164160 374972 164212
rect 375748 164160 375800 164212
rect 375932 164160 375984 164212
rect 393964 164160 394016 164212
rect 356704 164092 356756 164144
rect 418436 164092 418488 164144
rect 52276 164024 52328 164076
rect 101036 164024 101088 164076
rect 358268 164024 358320 164076
rect 421012 164024 421064 164076
rect 49424 163956 49476 164008
rect 98460 163956 98512 164008
rect 367836 163956 367888 164008
rect 430948 163956 431000 164008
rect 50896 163888 50948 163940
rect 103520 163888 103572 163940
rect 211988 163888 212040 163940
rect 265900 163888 265952 163940
rect 358360 163888 358412 163940
rect 423496 163888 423548 163940
rect 52184 163820 52236 163872
rect 105912 163820 105964 163872
rect 110788 163820 110840 163872
rect 111156 163820 111208 163872
rect 196624 163820 196676 163872
rect 204904 163820 204956 163872
rect 285956 163820 286008 163872
rect 362500 163820 362552 163872
rect 428188 163820 428240 163872
rect 438860 163820 438912 163872
rect 516600 163820 516652 163872
rect 47952 163752 48004 163804
rect 52276 163752 52328 163804
rect 59912 163752 59964 163804
rect 145932 163752 145984 163804
rect 213184 163752 213236 163804
rect 303436 163752 303488 163804
rect 373540 163752 373592 163804
rect 475844 163752 475896 163804
rect 50804 163684 50856 163736
rect 108212 163684 108264 163736
rect 110512 163684 110564 163736
rect 196808 163684 196860 163736
rect 206376 163684 206428 163736
rect 298468 163684 298520 163736
rect 370780 163684 370832 163736
rect 473452 163684 473504 163736
rect 59084 163616 59136 163668
rect 148508 163616 148560 163668
rect 207756 163616 207808 163668
rect 300860 163616 300912 163668
rect 367928 163616 367980 163668
rect 470968 163616 471020 163668
rect 510528 163616 510580 163668
rect 517520 163616 517572 163668
rect 58900 163548 58952 163600
rect 150900 163548 150952 163600
rect 209136 163548 209188 163600
rect 305920 163548 305972 163600
rect 372068 163548 372120 163600
rect 478420 163548 478472 163600
rect 60004 163480 60056 163532
rect 153384 163480 153436 163532
rect 214748 163480 214800 163532
rect 313372 163480 313424 163532
rect 366640 163480 366692 163532
rect 483388 163480 483440 163532
rect 218612 163412 218664 163464
rect 219716 163412 219768 163464
rect 220452 163412 220504 163464
rect 373172 163140 373224 163192
rect 374184 163140 374236 163192
rect 375288 163140 375340 163192
rect 53196 163004 53248 163056
rect 113456 163004 113508 163056
rect 123024 163004 123076 163056
rect 373724 163004 373776 163056
rect 374920 163004 374972 163056
rect 429752 163004 429804 163056
rect 52276 162936 52328 162988
rect 114376 162936 114428 162988
rect 217140 162936 217192 162988
rect 236644 162936 236696 162988
rect 375288 162936 375340 162988
rect 431960 162936 432012 162988
rect 55772 162868 55824 162920
rect 118056 162868 118108 162920
rect 197452 162868 197504 162920
rect 200120 162868 200172 162920
rect 220452 162868 220504 162920
rect 267556 162868 267608 162920
rect 375748 162868 375800 162920
rect 436928 162868 436980 162920
rect 50528 162800 50580 162852
rect 155960 162800 156012 162852
rect 210608 162800 210660 162852
rect 320916 162800 320968 162852
rect 356704 162800 356756 162852
rect 357072 162800 357124 162852
rect 365168 162800 365220 162852
rect 458364 162800 458416 162852
rect 517612 162800 517664 162852
rect 517888 162800 517940 162852
rect 56140 162732 56192 162784
rect 135996 162732 136048 162784
rect 214564 162732 214616 162784
rect 293224 162732 293276 162784
rect 369216 162732 369268 162784
rect 455788 162732 455840 162784
rect 517520 162732 517572 162784
rect 517980 162732 518032 162784
rect 55128 162664 55180 162716
rect 133420 162664 133472 162716
rect 211804 162664 211856 162716
rect 280804 162664 280856 162716
rect 370688 162664 370740 162716
rect 453396 162664 453448 162716
rect 56324 162596 56376 162648
rect 130844 162596 130896 162648
rect 218796 162596 218848 162648
rect 283748 162596 283800 162648
rect 366548 162596 366600 162648
rect 448244 162596 448296 162648
rect 55036 162528 55088 162580
rect 128360 162528 128412 162580
rect 204996 162528 205048 162580
rect 263692 162528 263744 162580
rect 360936 162528 360988 162580
rect 435916 162528 435968 162580
rect 54944 162460 54996 162512
rect 122748 162460 122800 162512
rect 123024 162460 123076 162512
rect 196716 162460 196768 162512
rect 214656 162460 214708 162512
rect 273444 162460 273496 162512
rect 371976 162460 372028 162512
rect 445852 162460 445904 162512
rect 56232 162392 56284 162444
rect 125876 162392 125928 162444
rect 210424 162392 210476 162444
rect 268292 162392 268344 162444
rect 363788 162392 363840 162444
rect 438492 162392 438544 162444
rect 53380 162324 53432 162376
rect 120724 162324 120776 162376
rect 183468 162324 183520 162376
rect 197360 162324 197412 162376
rect 218888 162324 218940 162376
rect 276112 162324 276164 162376
rect 373356 162324 373408 162376
rect 443460 162324 443512 162376
rect 53288 162256 53340 162308
rect 116032 162256 116084 162308
rect 202144 162256 202196 162308
rect 256148 162256 256200 162308
rect 343456 162256 343508 162308
rect 356704 162256 356756 162308
rect 374828 162256 374880 162308
rect 440884 162256 440936 162308
rect 503260 162256 503312 162308
rect 517520 162256 517572 162308
rect 56048 162188 56100 162240
rect 118332 162188 118384 162240
rect 183192 162188 183244 162240
rect 197452 162188 197504 162240
rect 211896 162188 211948 162240
rect 258356 162188 258408 162240
rect 369124 162188 369176 162240
rect 433524 162188 433576 162240
rect 100024 162120 100076 162172
rect 100760 162120 100812 162172
rect 112812 162120 112864 162172
rect 113088 162120 113140 162172
rect 197820 162120 197872 162172
rect 209044 162120 209096 162172
rect 253572 162120 253624 162172
rect 343364 162120 343416 162172
rect 357532 162120 357584 162172
rect 362408 162120 362460 162172
rect 410616 162120 410668 162172
rect 415308 162120 415360 162172
rect 418252 162120 418304 162172
rect 503628 162120 503680 162172
rect 517612 162120 517664 162172
rect 53472 162052 53524 162104
rect 110972 162052 111024 162104
rect 210516 162052 210568 162104
rect 250628 162052 250680 162104
rect 367744 162052 367796 162104
rect 408316 162052 408368 162104
rect 49332 161984 49384 162036
rect 90732 161984 90784 162036
rect 216036 161984 216088 162036
rect 248236 161984 248288 162036
rect 374736 161984 374788 162036
rect 413560 161984 413612 162036
rect 56416 161916 56468 161968
rect 88340 161916 88392 161968
rect 378784 161916 378836 161968
rect 416044 161916 416096 161968
rect 54852 161848 54904 161900
rect 113180 161848 113232 161900
rect 428740 161508 428792 161560
rect 435732 161508 435784 161560
rect 98644 161440 98696 161492
rect 103796 161440 103848 161492
rect 56876 161372 56928 161424
rect 115940 161372 115992 161424
rect 219532 161372 219584 161424
rect 267740 161372 267792 161424
rect 379980 161372 380032 161424
rect 426440 161372 426492 161424
rect 58624 161304 58676 161356
rect 106372 161304 106424 161356
rect 218520 161304 218572 161356
rect 266360 161304 266412 161356
rect 379704 161304 379756 161356
rect 425060 161304 425112 161356
rect 54208 161236 54260 161288
rect 55036 161236 55088 161288
rect 99380 161236 99432 161288
rect 214288 161236 214340 161288
rect 260840 161236 260892 161288
rect 219624 161168 219676 161220
rect 264980 161168 265032 161220
rect 218980 161100 219032 161152
rect 219348 161100 219400 161152
rect 263600 161100 263652 161152
rect 217876 161032 217928 161084
rect 258080 161032 258132 161084
rect 52920 160964 52972 161016
rect 57796 160964 57848 161016
rect 95240 160964 95292 161016
rect 54300 160896 54352 160948
rect 59084 160896 59136 160948
rect 96620 160896 96672 160948
rect 51448 160828 51500 160880
rect 55128 160828 55180 160880
rect 98000 160828 98052 160880
rect 373816 160828 373868 160880
rect 374736 160828 374788 160880
rect 430580 160828 430632 160880
rect 60004 160760 60056 160812
rect 106280 160760 106332 160812
rect 371700 160760 371752 160812
rect 373632 160760 373684 160812
rect 433340 160760 433392 160812
rect 47860 160692 47912 160744
rect 59360 160692 59412 160744
rect 118700 160692 118752 160744
rect 213276 160692 213328 160744
rect 273260 160692 273312 160744
rect 370412 160692 370464 160744
rect 374552 160692 374604 160744
rect 437388 160692 437440 160744
rect 58716 160556 58768 160608
rect 60004 160556 60056 160608
rect 212172 160420 212224 160472
rect 213276 160420 213328 160472
rect 58624 160080 58676 160132
rect 59176 160080 59228 160132
rect 214288 160080 214340 160132
rect 214748 160080 214800 160132
rect 218244 160080 218296 160132
rect 218520 160080 218572 160132
rect 379796 160080 379848 160132
rect 379980 160080 380032 160132
rect 214840 160012 214892 160064
rect 259552 160012 259604 160064
rect 376300 160012 376352 160064
rect 420920 160012 420972 160064
rect 216404 159944 216456 159996
rect 259460 159944 259512 159996
rect 377680 159944 377732 159996
rect 419540 159944 419592 159996
rect 215760 159536 215812 159588
rect 216404 159536 216456 159588
rect 376392 159400 376444 159452
rect 379612 159400 379664 159452
rect 418160 159400 418212 159452
rect 370872 159332 370924 159384
rect 372252 159332 372304 159384
rect 428740 159332 428792 159384
rect 376668 158720 376720 158772
rect 377680 158720 377732 158772
rect 217140 156612 217192 156664
rect 217876 156612 217928 156664
rect 215024 148996 215076 149048
rect 274732 148996 274784 149048
rect 380808 148996 380860 149048
rect 429200 148996 429252 149048
rect 213368 148928 213420 148980
rect 240140 148928 240192 148980
rect 379888 148928 379940 148980
rect 412732 148928 412784 148980
rect 214932 148860 214984 148912
rect 241520 148860 241572 148912
rect 373724 148860 373776 148912
rect 375012 148860 375064 148912
rect 400220 148860 400272 148912
rect 215668 148792 215720 148844
rect 238760 148792 238812 148844
rect 48044 148656 48096 148708
rect 52092 148656 52144 148708
rect 78680 148656 78732 148708
rect 46480 148588 46532 148640
rect 53380 148588 53432 148640
rect 80060 148588 80112 148640
rect 49148 148520 49200 148572
rect 53288 148520 53340 148572
rect 81440 148520 81492 148572
rect 372344 148520 372396 148572
rect 375012 148520 375064 148572
rect 401600 148520 401652 148572
rect 54760 148452 54812 148504
rect 110788 148452 110840 148504
rect 370228 148452 370280 148504
rect 371976 148452 372028 148504
rect 398840 148452 398892 148504
rect 54944 148384 54996 148436
rect 113180 148384 113232 148436
rect 370320 148384 370372 148436
rect 52184 148316 52236 148368
rect 110512 148316 110564 148368
rect 213460 148316 213512 148368
rect 215944 148316 215996 148368
rect 271880 148316 271932 148368
rect 380256 148384 380308 148436
rect 423680 148384 423732 148436
rect 376392 148316 376444 148368
rect 377680 148248 377732 148300
rect 380256 148248 380308 148300
rect 434720 148316 434772 148368
rect 213184 147636 213236 147688
rect 215024 147636 215076 147688
rect 374368 147636 374420 147688
rect 376392 147636 376444 147688
rect 379428 147636 379480 147688
rect 379888 147636 379940 147688
rect 59728 147568 59780 147620
rect 107660 147568 107712 147620
rect 379336 147568 379388 147620
rect 426532 147568 426584 147620
rect 57060 147500 57112 147552
rect 104900 147500 104952 147552
rect 378968 147364 379020 147416
rect 379336 147364 379388 147416
rect 213460 146276 213512 146328
rect 47768 146208 47820 146260
rect 51816 146208 51868 146260
rect 56232 146208 56284 146260
rect 57980 146208 58032 146260
rect 58900 146208 58952 146260
rect 59820 146208 59872 146260
rect 102140 146208 102192 146260
rect 179052 146208 179104 146260
rect 197544 146208 197596 146260
rect 219072 146208 219124 146260
rect 255320 146208 255372 146260
rect 274824 146208 274876 146260
rect 356796 146208 356848 146260
rect 376208 146208 376260 146260
rect 376852 146208 376904 146260
rect 377956 146208 378008 146260
rect 411260 146208 411312 146260
rect 53104 146140 53156 146192
rect 86960 146140 87012 146192
rect 179696 146140 179748 146192
rect 197636 146140 197688 146192
rect 236644 146140 236696 146192
rect 256700 146140 256752 146192
rect 276020 146140 276072 146192
rect 356612 146140 356664 146192
rect 375840 146140 375892 146192
rect 379060 146140 379112 146192
rect 379244 146140 379296 146192
rect 411352 146140 411404 146192
rect 500224 146140 500276 146192
rect 518072 146140 518124 146192
rect 518256 146140 518308 146192
rect 56968 146072 57020 146124
rect 58992 146072 59044 146124
rect 59452 146072 59504 146124
rect 88432 146072 88484 146124
rect 219808 146072 219860 146124
rect 253940 146072 253992 146124
rect 338488 146072 338540 146124
rect 357624 146072 357676 146124
rect 378600 146072 378652 146124
rect 409880 146072 409932 146124
rect 498660 146072 498712 146124
rect 517704 146072 517756 146124
rect 57980 146004 58032 146056
rect 89812 146004 89864 146056
rect 219900 146004 219952 146056
rect 252560 146004 252612 146056
rect 340236 146004 340288 146056
rect 356888 146004 356940 146056
rect 376852 146004 376904 146056
rect 408500 146004 408552 146056
rect 54852 145936 54904 145988
rect 85580 145936 85632 145988
rect 219256 145936 219308 145988
rect 251180 145936 251232 145988
rect 376484 145936 376536 145988
rect 405740 145936 405792 145988
rect 58716 145868 58768 145920
rect 84292 145868 84344 145920
rect 217968 145868 218020 145920
rect 249800 145868 249852 145920
rect 374276 145868 374328 145920
rect 403072 145868 403124 145920
rect 56508 145800 56560 145852
rect 84200 145800 84252 145852
rect 219164 145800 219216 145852
rect 248420 145800 248472 145852
rect 376576 145800 376628 145852
rect 402980 145800 403032 145852
rect 48964 145732 49016 145784
rect 54392 145732 54444 145784
rect 82820 145732 82872 145784
rect 215116 145732 215168 145784
rect 244372 145732 244424 145784
rect 375196 145732 375248 145784
rect 378508 145732 378560 145784
rect 404360 145732 404412 145784
rect 58992 145664 59044 145716
rect 91192 145664 91244 145716
rect 216128 145664 216180 145716
rect 244280 145664 244332 145716
rect 375288 145664 375340 145716
rect 397460 145664 397512 145716
rect 57060 145596 57112 145648
rect 91100 145596 91152 145648
rect 216588 145596 216640 145648
rect 247040 145596 247092 145648
rect 280068 145596 280120 145648
rect 356612 145596 356664 145648
rect 358820 145596 358872 145648
rect 378048 145596 378100 145648
rect 378600 145596 378652 145648
rect 378784 145596 378836 145648
rect 407212 145596 407264 145648
rect 517704 145596 517756 145648
rect 580356 145596 580408 145648
rect 46204 145528 46256 145580
rect 59820 145528 59872 145580
rect 93860 145528 93912 145580
rect 191748 145528 191800 145580
rect 198004 145528 198056 145580
rect 204904 145528 204956 145580
rect 214656 145528 214708 145580
rect 245660 145528 245712 145580
rect 351644 145528 351696 145580
rect 358084 145528 358136 145580
rect 358728 145528 358780 145580
rect 510528 145528 510580 145580
rect 518256 145528 518308 145580
rect 580264 145528 580316 145580
rect 51816 145460 51868 145512
rect 77300 145460 77352 145512
rect 215392 145460 215444 145512
rect 242900 145460 242952 145512
rect 378876 145460 378928 145512
rect 396080 145460 396132 145512
rect 48136 145392 48188 145444
rect 54576 145392 54628 145444
rect 75920 145392 75972 145444
rect 218612 145392 218664 145444
rect 236092 145392 236144 145444
rect 376116 145392 376168 145444
rect 376576 145392 376628 145444
rect 379060 145392 379112 145444
rect 396172 145392 396224 145444
rect 46388 145324 46440 145376
rect 54668 145324 54720 145376
rect 76012 145324 76064 145376
rect 216220 145324 216272 145376
rect 218980 145324 219032 145376
rect 236000 145324 236052 145376
rect 378968 145324 379020 145376
rect 393964 145324 394016 145376
rect 56140 145256 56192 145308
rect 59452 145256 59504 145308
rect 217140 145120 217192 145172
rect 251272 145256 251324 145308
rect 218520 145052 218572 145104
rect 219072 145052 219124 145104
rect 215392 144984 215444 145036
rect 216220 144984 216272 145036
rect 218796 144984 218848 145036
rect 219900 144984 219952 145036
rect 215852 144916 215904 144968
rect 216128 144916 216180 144968
rect 217048 144916 217100 144968
rect 217968 144916 218020 144968
rect 218888 144916 218940 144968
rect 219256 144916 219308 144968
rect 54484 144848 54536 144900
rect 55956 144848 56008 144900
rect 56508 144848 56560 144900
rect 209596 144848 209648 144900
rect 214564 144848 214616 144900
rect 372436 144848 372488 144900
rect 375104 144916 375156 144968
rect 375288 144916 375340 144968
rect 373908 144848 373960 144900
rect 378784 144848 378836 144900
rect 52000 144780 52052 144832
rect 58716 144780 58768 144832
rect 213736 144780 213788 144832
rect 216036 144780 216088 144832
rect 216588 144780 216640 144832
rect 374092 144780 374144 144832
rect 378876 144780 378928 144832
rect 51908 144712 51960 144764
rect 57060 144712 57112 144764
rect 213644 144712 213696 144764
rect 214656 144712 214708 144764
rect 50344 144644 50396 144696
rect 55864 144644 55916 144696
rect 56416 144644 56468 144696
rect 213552 144644 213604 144696
rect 216128 144644 216180 144696
rect 216312 144644 216364 144696
rect 374276 144644 374328 144696
rect 375196 144644 375248 144696
rect 49240 144576 49292 144628
rect 58624 144576 58676 144628
rect 212080 144576 212132 144628
rect 215024 144576 215076 144628
rect 520188 79976 520240 80028
rect 580448 79976 580500 80028
rect 207664 70320 207716 70372
rect 216680 70320 216732 70372
rect 365076 70320 365128 70372
rect 376944 70320 376996 70372
rect 46848 68960 46900 69012
rect 56876 68960 56928 69012
rect 358084 68416 358136 68468
rect 358728 68416 358780 68468
rect 376944 68280 376996 68332
rect 204904 67600 204956 67652
rect 216680 67600 216732 67652
rect 218796 61072 218848 61124
rect 219072 61072 219124 61124
rect 379060 59712 379112 59764
rect 397092 59712 397144 59764
rect 218612 59644 218664 59696
rect 237104 59644 237156 59696
rect 378876 59644 378928 59696
rect 396080 59644 396132 59696
rect 54576 59576 54628 59628
rect 77116 59576 77168 59628
rect 218520 59576 218572 59628
rect 255872 59576 255924 59628
rect 378968 59576 379020 59628
rect 418160 59576 418212 59628
rect 54392 59508 54444 59560
rect 83096 59508 83148 59560
rect 217876 59508 217928 59560
rect 256976 59508 257028 59560
rect 375932 59508 375984 59560
rect 416964 59508 417016 59560
rect 55036 59440 55088 59492
rect 99472 59440 99524 59492
rect 219348 59440 219400 59492
rect 263876 59440 263928 59492
rect 377680 59440 377732 59492
rect 423956 59440 424008 59492
rect 49516 59372 49568 59424
rect 113548 59372 113600 59424
rect 214748 59372 214800 59424
rect 261760 59372 261812 59424
rect 362224 59372 362276 59424
rect 418436 59372 418488 59424
rect 55956 59304 56008 59356
rect 84200 59304 84252 59356
rect 217968 59304 218020 59356
rect 358084 59304 358136 59356
rect 59820 59236 59872 59288
rect 94504 59236 94556 59288
rect 375196 59236 375248 59288
rect 403072 59236 403124 59288
rect 57796 59168 57848 59220
rect 95884 59168 95936 59220
rect 214840 59168 214892 59220
rect 260656 59168 260708 59220
rect 379612 59168 379664 59220
rect 419448 59168 419500 59220
rect 59084 59100 59136 59152
rect 96988 59100 97040 59152
rect 215760 59100 215812 59152
rect 262772 59100 262824 59152
rect 279240 59100 279292 59152
rect 356612 59100 356664 59152
rect 376668 59100 376720 59152
rect 420644 59100 420696 59152
rect 58900 59032 58952 59084
rect 102784 59032 102836 59084
rect 205548 59032 205600 59084
rect 290924 59032 290976 59084
rect 376300 59032 376352 59084
rect 421748 59032 421800 59084
rect 56048 58964 56100 59016
rect 101772 58964 101824 59016
rect 208952 58964 209004 59016
rect 298468 58964 298520 59016
rect 379704 58964 379756 59016
rect 425244 58964 425296 59016
rect 55864 58896 55916 58948
rect 103888 58896 103940 58948
rect 215208 58896 215260 58948
rect 313372 58896 313424 58948
rect 373264 58896 373316 58948
rect 423496 58896 423548 58948
rect 54760 58828 54812 58880
rect 111156 58828 111208 58880
rect 206836 58828 206888 58880
rect 305920 58828 305972 58880
rect 363604 58828 363656 58880
rect 425980 58828 426032 58880
rect 42616 58760 42668 58812
rect 115940 58760 115992 58812
rect 201408 58760 201460 58812
rect 318432 58760 318484 58812
rect 366456 58760 366508 58812
rect 465908 58760 465960 58812
rect 50068 58692 50120 58744
rect 148508 58692 148560 58744
rect 202788 58692 202840 58744
rect 325884 58692 325936 58744
rect 358636 58692 358688 58744
rect 485964 58692 486016 58744
rect 53564 58624 53616 58676
rect 150900 58624 150952 58676
rect 219256 58624 219308 58676
rect 428188 58624 428240 58676
rect 216404 58556 216456 58608
rect 259460 58556 259512 58608
rect 376116 58556 376168 58608
rect 404176 58556 404228 58608
rect 57888 57876 57940 57928
rect 204904 57876 204956 57928
rect 210976 57876 211028 57928
rect 323308 57876 323360 57928
rect 343180 57876 343232 57928
rect 357532 57876 357584 57928
rect 364984 57876 365036 57928
rect 478420 57876 478472 57928
rect 503352 57876 503404 57928
rect 517612 57876 517664 57928
rect 52368 57808 52420 57860
rect 145564 57808 145616 57860
rect 183284 57808 183336 57860
rect 197452 57808 197504 57860
rect 212356 57808 212408 57860
rect 315764 57808 315816 57860
rect 343456 57808 343508 57860
rect 356704 57808 356756 57860
rect 360844 57808 360896 57860
rect 443460 57808 443512 57860
rect 503260 57808 503312 57860
rect 517520 57808 517572 57860
rect 44088 57740 44140 57792
rect 123484 57740 123536 57792
rect 183468 57740 183520 57792
rect 197360 57740 197412 57792
rect 218704 57740 218756 57792
rect 320916 57740 320968 57792
rect 358176 57740 358228 57792
rect 440884 57740 440936 57792
rect 52828 57672 52880 57724
rect 130844 57672 130896 57724
rect 208308 57672 208360 57724
rect 308496 57672 308548 57724
rect 363696 57672 363748 57724
rect 445852 57672 445904 57724
rect 54944 57604 54996 57656
rect 57244 57536 57296 57588
rect 57888 57536 57940 57588
rect 58072 57604 58124 57656
rect 133236 57604 133288 57656
rect 216496 57604 216548 57656
rect 310980 57604 311032 57656
rect 374644 57604 374696 57656
rect 451004 57604 451056 57656
rect 112076 57536 112128 57588
rect 213828 57536 213880 57588
rect 303436 57536 303488 57588
rect 362316 57536 362368 57588
rect 438492 57536 438544 57588
rect 39948 57468 40000 57520
rect 90732 57468 90784 57520
rect 211068 57468 211120 57520
rect 295892 57468 295944 57520
rect 371884 57468 371936 57520
rect 435916 57468 435968 57520
rect 55128 57400 55180 57452
rect 98092 57400 98144 57452
rect 218336 57400 218388 57452
rect 300860 57400 300912 57452
rect 370596 57400 370648 57452
rect 433524 57400 433576 57452
rect 53656 57332 53708 57384
rect 88340 57332 88392 57384
rect 212448 57332 212500 57384
rect 293316 57332 293368 57384
rect 376024 57332 376076 57384
rect 430948 57332 431000 57384
rect 55496 57264 55548 57316
rect 58072 57264 58124 57316
rect 59268 57264 59320 57316
rect 93676 57264 93728 57316
rect 215300 57264 215352 57316
rect 287612 57264 287664 57316
rect 370504 57264 370556 57316
rect 416044 57264 416096 57316
rect 51816 57196 51868 57248
rect 78220 57196 78272 57248
rect 218796 57196 218848 57248
rect 265900 57196 265952 57248
rect 379152 57196 379204 57248
rect 415492 57196 415544 57248
rect 54668 57128 54720 57180
rect 76012 57128 76064 57180
rect 58716 56516 58768 56568
rect 85396 56516 85448 56568
rect 214932 56516 214984 56568
rect 241612 56516 241664 56568
rect 375012 56516 375064 56568
rect 401692 56516 401744 56568
rect 53196 56448 53248 56500
rect 113180 56448 113232 56500
rect 215668 56448 215720 56500
rect 239220 56448 239272 56500
rect 374552 56448 374604 56500
rect 438308 56448 438360 56500
rect 59912 56380 59964 56432
rect 108028 56380 108080 56432
rect 218980 56380 219032 56432
rect 236000 56380 236052 56432
rect 372252 56380 372304 56432
rect 435732 56380 435784 56432
rect 59176 56312 59228 56364
rect 107384 56312 107436 56364
rect 215024 56312 215076 56364
rect 271236 56312 271288 56364
rect 376392 56312 376444 56364
rect 433340 56312 433392 56364
rect 60004 56244 60056 56296
rect 106372 56244 106424 56296
rect 219532 56244 219584 56296
rect 268476 56244 268528 56296
rect 379336 56244 379388 56296
rect 427636 56244 427688 56296
rect 57060 56176 57112 56228
rect 92112 56176 92164 56228
rect 218244 56176 218296 56228
rect 266360 56176 266412 56228
rect 379796 56176 379848 56228
rect 426440 56176 426492 56228
rect 56140 56108 56192 56160
rect 88708 56108 88760 56160
rect 219072 56108 219124 56160
rect 253388 56108 253440 56160
rect 379980 56108 380032 56160
rect 414572 56108 414624 56160
rect 54852 56040 54904 56092
rect 86500 56040 86552 56092
rect 218888 56040 218940 56092
rect 251180 56040 251232 56092
rect 379428 56040 379480 56092
rect 412640 56040 412692 56092
rect 53288 55972 53340 56024
rect 81808 55972 81860 56024
rect 219164 55972 219216 56024
rect 248604 55972 248656 56024
rect 376208 55972 376260 56024
rect 408684 55972 408736 56024
rect 52092 55904 52144 55956
rect 79508 55904 79560 55956
rect 215852 55904 215904 55956
rect 245292 55904 245344 55956
rect 379244 55904 379296 55956
rect 411260 55904 411312 55956
rect 49608 55836 49660 55888
rect 157432 55836 157484 55888
rect 213460 55836 213512 55888
rect 275468 55836 275520 55888
rect 371976 55836 372028 55888
rect 399484 55836 399536 55888
rect 219992 55768 220044 55820
rect 408316 55768 408368 55820
rect 213184 55700 213236 55752
rect 273260 55700 273312 55752
rect 55772 55156 55824 55208
rect 117320 55156 117372 55208
rect 216220 55156 216272 55208
rect 242900 55156 242952 55208
rect 375748 55156 375800 55208
rect 436100 55156 436152 55208
rect 52276 55088 52328 55140
rect 113272 55088 113324 55140
rect 215944 55088 215996 55140
rect 271880 55088 271932 55140
rect 375104 55088 375156 55140
rect 397460 55088 397512 55140
rect 55680 55020 55732 55072
rect 114560 55020 114612 55072
rect 216128 55020 216180 55072
rect 269120 55020 269172 55072
rect 374184 55020 374236 55072
rect 431960 55020 432012 55072
rect 52184 54952 52236 55004
rect 109040 54952 109092 55004
rect 219716 54952 219768 55004
rect 266452 54952 266504 55004
rect 374736 54952 374788 55004
rect 430580 54952 430632 55004
rect 53104 54884 53156 54936
rect 86960 54884 87012 54936
rect 219624 54884 219676 54936
rect 264980 54884 265032 54936
rect 374920 54884 374972 54936
rect 429200 54884 429252 54936
rect 58624 54816 58676 54868
rect 92480 54816 92532 54868
rect 219808 54816 219860 54868
rect 253940 54816 253992 54868
rect 377956 54816 378008 54868
rect 411352 54816 411404 54868
rect 56232 54748 56284 54800
rect 89720 54748 89772 54800
rect 217140 54748 217192 54800
rect 251364 54748 251416 54800
rect 378048 54748 378100 54800
rect 409880 54748 409932 54800
rect 58992 54680 59044 54732
rect 91192 54680 91244 54732
rect 217048 54680 217100 54732
rect 249800 54680 249852 54732
rect 376484 54680 376536 54732
rect 405832 54680 405884 54732
rect 53380 54612 53432 54664
rect 80060 54612 80112 54664
rect 216036 54612 216088 54664
rect 247040 54612 247092 54664
rect 375288 54612 375340 54664
rect 404360 54612 404412 54664
rect 214656 54544 214708 54596
rect 245660 54544 245712 54596
rect 378784 54544 378836 54596
rect 407212 54544 407264 54596
rect 215116 54476 215168 54528
rect 244372 54476 244424 54528
rect 373724 54476 373776 54528
rect 400220 54476 400272 54528
rect 213276 54408 213328 54460
rect 273352 54408 273404 54460
rect 373632 54408 373684 54460
rect 433432 54408 433484 54460
rect 213368 54340 213420 54392
rect 240140 54340 240192 54392
rect 214564 54272 214616 54324
rect 237380 54272 237432 54324
rect 2780 20340 2832 20392
rect 4804 20340 4856 20392
rect 572 3408 624 3460
rect 57244 3408 57296 3460
rect 125876 3408 125928 3460
rect 366364 3408 366416 3460
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 639606 3464 684247
rect 3424 639600 3476 639606
rect 3424 639542 3476 639548
rect 3514 632088 3570 632097
rect 3514 632023 3570 632032
rect 3422 580000 3478 580009
rect 3422 579935 3478 579944
rect 3436 561134 3464 579935
rect 3424 561128 3476 561134
rect 3424 561070 3476 561076
rect 3424 559564 3476 559570
rect 3424 559506 3476 559512
rect 2964 411256 3016 411262
rect 2964 411198 3016 411204
rect 2976 410553 3004 411198
rect 2962 410544 3018 410553
rect 2962 410479 3018 410488
rect 3332 358760 3384 358766
rect 3332 358702 3384 358708
rect 3344 358465 3372 358702
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3056 202836 3108 202842
rect 3056 202778 3108 202784
rect 3068 201929 3096 202778
rect 3054 201920 3110 201929
rect 3054 201855 3110 201864
rect 3436 58585 3464 559506
rect 3528 555490 3556 632023
rect 18604 630760 18656 630766
rect 18604 630702 18656 630708
rect 4804 556844 4856 556850
rect 4804 556786 4856 556792
rect 3516 555484 3568 555490
rect 3516 555426 3568 555432
rect 3516 553444 3568 553450
rect 3516 553386 3568 553392
rect 3528 97617 3556 553386
rect 3608 540116 3660 540122
rect 3608 540058 3660 540064
rect 3620 514865 3648 540058
rect 3606 514856 3662 514865
rect 3606 514791 3662 514800
rect 3606 475416 3662 475425
rect 3606 475351 3662 475360
rect 3620 462641 3648 475351
rect 3606 462632 3662 462641
rect 3606 462567 3662 462576
rect 3514 97608 3570 97617
rect 3514 97543 3570 97552
rect 3422 58576 3478 58585
rect 3422 58511 3478 58520
rect 4816 20398 4844 556786
rect 14464 476808 14516 476814
rect 14464 476750 14516 476756
rect 14476 411262 14504 476750
rect 14464 411256 14516 411262
rect 14464 411198 14516 411204
rect 18616 358766 18644 630702
rect 40052 549234 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 57888 700324 57940 700330
rect 57888 700266 57940 700272
rect 42062 632088 42118 632097
rect 42062 632023 42118 632032
rect 40040 549228 40092 549234
rect 40040 549170 40092 549176
rect 41328 468852 41380 468858
rect 41328 468794 41380 468800
rect 39856 468784 39908 468790
rect 39856 468726 39908 468732
rect 18604 358760 18656 358766
rect 18604 358702 18656 358708
rect 39868 164354 39896 468726
rect 39948 460488 40000 460494
rect 39948 460430 40000 460436
rect 39856 164348 39908 164354
rect 39856 164290 39908 164296
rect 39960 57526 39988 460430
rect 41340 164286 41368 468794
rect 42076 202842 42104 632023
rect 54852 625320 54904 625326
rect 54852 625262 54904 625268
rect 54864 559774 54892 625262
rect 55128 625252 55180 625258
rect 55128 625194 55180 625200
rect 55036 622668 55088 622674
rect 55036 622610 55088 622616
rect 54944 622600 54996 622606
rect 54944 622542 54996 622548
rect 54852 559768 54904 559774
rect 54852 559710 54904 559716
rect 54956 543250 54984 622542
rect 55048 543590 55076 622610
rect 55140 543658 55168 625194
rect 56508 625184 56560 625190
rect 56508 625126 56560 625132
rect 56324 622532 56376 622538
rect 56324 622474 56376 622480
rect 55128 543652 55180 543658
rect 55128 543594 55180 543600
rect 55036 543584 55088 543590
rect 55036 543526 55088 543532
rect 54944 543244 54996 543250
rect 54944 543186 54996 543192
rect 56336 543182 56364 622474
rect 56416 622464 56468 622470
rect 56416 622406 56468 622412
rect 56428 543318 56456 622406
rect 56520 543386 56548 625126
rect 57796 623892 57848 623898
rect 57796 623834 57848 623840
rect 57702 620664 57758 620673
rect 57702 620599 57758 620608
rect 57518 614408 57574 614417
rect 57518 614343 57574 614352
rect 57426 589928 57482 589937
rect 57426 589863 57482 589872
rect 57334 586392 57390 586401
rect 57334 586327 57390 586336
rect 57058 577688 57114 577697
rect 57058 577623 57114 577632
rect 57072 559910 57100 577623
rect 57150 574968 57206 574977
rect 57150 574903 57206 574912
rect 57164 560250 57192 574903
rect 57348 572354 57376 586327
rect 57336 572348 57388 572354
rect 57336 572290 57388 572296
rect 57334 571568 57390 571577
rect 57334 571503 57390 571512
rect 57242 565448 57298 565457
rect 57242 565383 57298 565392
rect 57152 560244 57204 560250
rect 57152 560186 57204 560192
rect 57060 559904 57112 559910
rect 57060 559846 57112 559852
rect 57256 545834 57284 565383
rect 57348 557054 57376 571503
rect 57440 558890 57468 589863
rect 57532 583778 57560 614343
rect 57610 593464 57666 593473
rect 57610 593399 57666 593408
rect 57520 583772 57572 583778
rect 57520 583714 57572 583720
rect 57518 583672 57574 583681
rect 57518 583607 57574 583616
rect 57428 558884 57480 558890
rect 57428 558826 57480 558832
rect 57336 557048 57388 557054
rect 57336 556990 57388 556996
rect 57532 551478 57560 583607
rect 57520 551472 57572 551478
rect 57520 551414 57572 551420
rect 57624 547398 57652 593399
rect 57716 552770 57744 620599
rect 57704 552764 57756 552770
rect 57704 552706 57756 552712
rect 57612 547392 57664 547398
rect 57612 547334 57664 547340
rect 57244 545828 57296 545834
rect 57244 545770 57296 545776
rect 57808 543522 57836 623834
rect 57900 599593 57928 700266
rect 104912 636886 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 170324 702434 170352 703520
rect 169772 702406 170352 702434
rect 137836 683188 137888 683194
rect 137836 683130 137888 683136
rect 104900 636880 104952 636886
rect 104900 636822 104952 636828
rect 100576 625796 100628 625802
rect 100576 625738 100628 625744
rect 124680 625796 124732 625802
rect 124680 625738 124732 625744
rect 83188 625592 83240 625598
rect 83188 625534 83240 625540
rect 77392 625184 77444 625190
rect 77392 625126 77444 625132
rect 59360 623960 59412 623966
rect 59360 623902 59412 623908
rect 59266 617808 59322 617817
rect 59266 617743 59322 617752
rect 59082 611688 59138 611697
rect 59082 611623 59138 611632
rect 58898 608288 58954 608297
rect 58898 608223 58954 608232
rect 57886 599584 57942 599593
rect 57886 599519 57942 599528
rect 57886 596048 57942 596057
rect 57886 595983 57942 595992
rect 57900 561202 57928 595983
rect 58624 583772 58676 583778
rect 58624 583714 58676 583720
rect 58530 568848 58586 568857
rect 58530 568783 58586 568792
rect 57888 561196 57940 561202
rect 57888 561138 57940 561144
rect 57796 543516 57848 543522
rect 57796 543458 57848 543464
rect 56508 543380 56560 543386
rect 56508 543322 56560 543328
rect 56416 543312 56468 543318
rect 56416 543254 56468 543260
rect 56324 543176 56376 543182
rect 56324 543118 56376 543124
rect 57900 509969 57928 561138
rect 58544 554130 58572 568783
rect 58532 554124 58584 554130
rect 58532 554066 58584 554072
rect 58636 543046 58664 583714
rect 58806 581088 58862 581097
rect 58806 581023 58862 581032
rect 58716 572348 58768 572354
rect 58716 572290 58768 572296
rect 58728 543454 58756 572290
rect 58716 543448 58768 543454
rect 58716 543390 58768 543396
rect 58820 543114 58848 581023
rect 58912 558210 58940 608223
rect 58990 602168 59046 602177
rect 58990 602103 59046 602112
rect 58900 558204 58952 558210
rect 58900 558146 58952 558152
rect 59004 551410 59032 602103
rect 59096 559842 59124 611623
rect 59174 605568 59230 605577
rect 59174 605503 59230 605512
rect 59084 559836 59136 559842
rect 59084 559778 59136 559784
rect 58992 551404 59044 551410
rect 58992 551346 59044 551352
rect 59188 548554 59216 605503
rect 59280 555626 59308 617743
rect 59268 555620 59320 555626
rect 59268 555562 59320 555568
rect 59176 548548 59228 548554
rect 59176 548490 59228 548496
rect 59372 547874 59400 623902
rect 69020 623824 69072 623830
rect 69020 623766 69072 623772
rect 69032 623084 69060 623766
rect 77404 623084 77432 625126
rect 80612 623892 80664 623898
rect 80612 623834 80664 623840
rect 80624 623084 80652 623834
rect 83200 623084 83228 625534
rect 88984 625320 89036 625326
rect 88984 625262 89036 625268
rect 86408 623892 86460 623898
rect 86408 623834 86460 623840
rect 86420 623084 86448 623834
rect 88996 623084 89024 625262
rect 92204 625252 92256 625258
rect 92204 625194 92256 625200
rect 94780 625252 94832 625258
rect 94780 625194 94832 625200
rect 92216 623084 92244 625194
rect 94792 623084 94820 625194
rect 98000 623960 98052 623966
rect 98000 623902 98052 623908
rect 98012 623084 98040 623902
rect 100588 623084 100616 625738
rect 115388 625728 115440 625734
rect 115388 625670 115440 625676
rect 124588 625728 124640 625734
rect 124588 625670 124640 625676
rect 112168 625660 112220 625666
rect 112168 625602 112220 625608
rect 109592 625524 109644 625530
rect 109592 625466 109644 625472
rect 106372 625456 106424 625462
rect 106372 625398 106424 625404
rect 103796 625388 103848 625394
rect 103796 625330 103848 625336
rect 103808 623084 103836 625330
rect 106384 623084 106412 625398
rect 109604 623084 109632 625466
rect 112180 623084 112208 625602
rect 115400 623084 115428 625670
rect 124496 625660 124548 625666
rect 124496 625602 124548 625608
rect 122840 625524 122892 625530
rect 122840 625466 122892 625472
rect 120908 625456 120960 625462
rect 120908 625398 120960 625404
rect 62960 622674 63250 622690
rect 62948 622668 63250 622674
rect 63000 622662 63250 622668
rect 62948 622610 63000 622616
rect 65524 622600 65576 622606
rect 65576 622548 65826 622554
rect 65524 622542 65826 622548
rect 65536 622526 65826 622542
rect 71240 622538 71622 622554
rect 71228 622532 71622 622538
rect 71280 622526 71622 622532
rect 71228 622474 71280 622480
rect 74632 622464 74684 622470
rect 59464 622390 60030 622418
rect 74684 622412 74842 622418
rect 74632 622406 74842 622412
rect 74644 622390 74842 622406
rect 117990 622402 118280 622418
rect 117990 622396 118292 622402
rect 117990 622390 118240 622396
rect 59464 552906 59492 622390
rect 120566 622390 120764 622418
rect 118240 622338 118292 622344
rect 59542 562788 59598 562797
rect 59542 562723 59598 562732
rect 59452 552900 59504 552906
rect 59452 552842 59504 552848
rect 59556 550050 59584 562723
rect 62120 560244 62172 560250
rect 62120 560186 62172 560192
rect 60030 560102 60320 560130
rect 60292 558754 60320 560102
rect 60740 558884 60792 558890
rect 60740 558826 60792 558832
rect 60280 558748 60332 558754
rect 60280 558690 60332 558696
rect 60752 557534 60780 558826
rect 62132 557534 62160 560186
rect 106280 560176 106332 560182
rect 62606 560102 62896 560130
rect 62764 558748 62816 558754
rect 62764 558690 62816 558696
rect 60752 557506 60964 557534
rect 62132 557506 62436 557534
rect 59544 550044 59596 550050
rect 59544 549986 59596 549992
rect 59372 547846 60320 547874
rect 58808 543108 58860 543114
rect 58808 543050 58860 543056
rect 58624 543040 58676 543046
rect 58624 542982 58676 542988
rect 60292 539963 60320 547846
rect 60936 539963 60964 557506
rect 61660 543720 61712 543726
rect 61660 543662 61712 543668
rect 61672 539963 61700 543662
rect 62408 539963 62436 557506
rect 62776 547262 62804 558690
rect 62868 558346 62896 560102
rect 65076 560102 65182 560130
rect 68402 560102 68784 560130
rect 70978 560102 71360 560130
rect 63500 559632 63552 559638
rect 63500 559574 63552 559580
rect 62856 558340 62908 558346
rect 62856 558282 62908 558288
rect 62764 547256 62816 547262
rect 62764 547198 62816 547204
rect 63132 547188 63184 547194
rect 63132 547130 63184 547136
rect 63144 539963 63172 547130
rect 63512 543930 63540 559574
rect 65076 557598 65104 560102
rect 67732 559904 67784 559910
rect 67732 559846 67784 559852
rect 67640 559700 67692 559706
rect 67640 559642 67692 559648
rect 64144 557592 64196 557598
rect 64144 557534 64196 557540
rect 65064 557592 65116 557598
rect 65064 557534 65116 557540
rect 63776 556912 63828 556918
rect 63776 556854 63828 556860
rect 63500 543924 63552 543930
rect 63500 543866 63552 543872
rect 63788 539963 63816 556854
rect 64156 543726 64184 557534
rect 64880 555552 64932 555558
rect 64880 555494 64932 555500
rect 64512 543924 64564 543930
rect 64892 543912 64920 555494
rect 66720 554056 66772 554062
rect 66720 553998 66772 554004
rect 65984 551336 66036 551342
rect 65984 551278 66036 551284
rect 64892 543884 65288 543912
rect 64512 543866 64564 543872
rect 64144 543720 64196 543726
rect 64144 543662 64196 543668
rect 64524 539963 64552 543866
rect 65260 539963 65288 543884
rect 65996 539963 66024 551278
rect 66732 539963 66760 553998
rect 67652 543912 67680 559642
rect 67744 557534 67772 559846
rect 68756 558482 68784 560102
rect 68744 558476 68796 558482
rect 68744 558418 68796 558424
rect 71044 558476 71096 558482
rect 71044 558418 71096 558424
rect 67744 557506 68876 557534
rect 67652 543884 68140 543912
rect 67364 543652 67416 543658
rect 67364 543594 67416 543600
rect 67376 539963 67404 543594
rect 68112 539963 68140 543884
rect 68848 539963 68876 557506
rect 69020 552696 69072 552702
rect 69020 552638 69072 552644
rect 69032 543912 69060 552638
rect 69112 549976 69164 549982
rect 69112 549918 69164 549924
rect 69124 544066 69152 549918
rect 70952 549908 71004 549914
rect 70952 549850 71004 549856
rect 69112 544060 69164 544066
rect 69112 544002 69164 544008
rect 70308 544060 70360 544066
rect 70308 544002 70360 544008
rect 69032 543884 69612 543912
rect 69584 539963 69612 543884
rect 70320 539963 70348 544002
rect 70964 539963 70992 549850
rect 71056 544406 71084 558418
rect 71332 558278 71360 560102
rect 73816 560102 74198 560130
rect 76774 560102 77064 560130
rect 71320 558272 71372 558278
rect 71320 558214 71372 558220
rect 73816 557938 73844 560102
rect 77036 558414 77064 560102
rect 79888 560102 79994 560130
rect 82570 560102 82768 560130
rect 85790 560102 86080 560130
rect 88366 560102 88656 560130
rect 78680 559768 78732 559774
rect 78680 559710 78732 559716
rect 77024 558408 77076 558414
rect 77024 558350 77076 558356
rect 74540 558204 74592 558210
rect 74540 558146 74592 558152
rect 71780 557932 71832 557938
rect 71780 557874 71832 557880
rect 73804 557932 73856 557938
rect 73804 557874 73856 557880
rect 71792 557534 71820 557874
rect 71792 557506 72464 557534
rect 71688 545760 71740 545766
rect 71688 545702 71740 545708
rect 71044 544400 71096 544406
rect 71044 544342 71096 544348
rect 71700 539963 71728 545702
rect 72436 539963 72464 557506
rect 73252 554192 73304 554198
rect 73252 554134 73304 554140
rect 73264 540138 73292 554134
rect 73804 543176 73856 543182
rect 73804 543118 73856 543124
rect 73188 540110 73292 540138
rect 73188 539920 73216 540110
rect 73816 539963 73844 543118
rect 74552 539963 74580 558146
rect 75920 552900 75972 552906
rect 75920 552842 75972 552848
rect 75276 552832 75328 552838
rect 75276 552774 75328 552780
rect 75288 539963 75316 552774
rect 75932 543946 75960 552842
rect 77392 552764 77444 552770
rect 77392 552706 77444 552712
rect 76748 548616 76800 548622
rect 76748 548558 76800 548564
rect 75932 543918 76052 543946
rect 76024 539963 76052 543918
rect 76760 539963 76788 548558
rect 77404 539963 77432 552706
rect 78692 543930 78720 559710
rect 79888 558210 79916 560102
rect 82740 558482 82768 560102
rect 82912 559836 82964 559842
rect 82912 559778 82964 559784
rect 82728 558476 82780 558482
rect 82728 558418 82780 558424
rect 80704 558340 80756 558346
rect 80704 558282 80756 558288
rect 79876 558204 79928 558210
rect 79876 558146 79928 558152
rect 78864 556980 78916 556986
rect 78864 556922 78916 556928
rect 78680 543924 78732 543930
rect 78680 543866 78732 543872
rect 78128 543176 78180 543182
rect 78128 543118 78180 543124
rect 78140 539963 78168 543118
rect 78876 539963 78904 556922
rect 80060 552764 80112 552770
rect 80060 552706 80112 552712
rect 80072 543946 80100 552706
rect 80716 550118 80744 558282
rect 82924 557534 82952 559778
rect 85580 559768 85632 559774
rect 85580 559710 85632 559716
rect 82924 557506 83228 557534
rect 81716 557048 81768 557054
rect 81716 556990 81768 556996
rect 80980 551540 81032 551546
rect 80980 551482 81032 551488
rect 80704 550112 80756 550118
rect 80704 550054 80756 550060
rect 79600 543924 79652 543930
rect 80072 543918 80376 543946
rect 79600 543866 79652 543872
rect 79612 539963 79640 543866
rect 80348 539963 80376 543918
rect 80992 539963 81020 551482
rect 81728 539963 81756 556990
rect 82452 545896 82504 545902
rect 82452 545838 82504 545844
rect 82464 539963 82492 545838
rect 83200 539963 83228 557506
rect 84568 547324 84620 547330
rect 84568 547266 84620 547272
rect 83924 543380 83976 543386
rect 83924 543322 83976 543328
rect 83936 539963 83964 543322
rect 84580 539963 84608 547266
rect 85592 543946 85620 559710
rect 85672 558408 85724 558414
rect 85672 558350 85724 558356
rect 85684 557534 85712 558350
rect 86052 558346 86080 560102
rect 86960 559904 87012 559910
rect 86960 559846 87012 559852
rect 86040 558340 86092 558346
rect 86040 558282 86092 558288
rect 85684 557506 86816 557534
rect 85592 543918 86080 543946
rect 85304 543380 85356 543386
rect 85304 543322 85356 543328
rect 85316 539963 85344 543322
rect 86052 539963 86080 543918
rect 86788 539963 86816 557506
rect 86972 543946 87000 559846
rect 87052 559836 87104 559842
rect 87052 559778 87104 559784
rect 87064 557534 87092 559778
rect 87064 557506 88196 557534
rect 86972 543918 87460 543946
rect 87432 539963 87460 543918
rect 88168 539963 88196 557506
rect 88628 552906 88656 560102
rect 91112 560102 91586 560130
rect 94162 560102 94544 560130
rect 88984 558476 89036 558482
rect 88984 558418 89036 558424
rect 88616 552900 88668 552906
rect 88616 552842 88668 552848
rect 88432 548684 88484 548690
rect 88432 548626 88484 548632
rect 88444 543930 88472 548626
rect 88432 543924 88484 543930
rect 88432 543866 88484 543872
rect 88996 543726 89024 558418
rect 89812 551472 89864 551478
rect 89812 551414 89864 551420
rect 89824 543930 89852 551414
rect 89628 543924 89680 543930
rect 89628 543866 89680 543872
rect 89812 543924 89864 543930
rect 89812 543866 89864 543872
rect 91008 543924 91060 543930
rect 91008 543866 91060 543872
rect 88984 543720 89036 543726
rect 88984 543662 89036 543668
rect 88892 543584 88944 543590
rect 88892 543526 88944 543532
rect 88904 539963 88932 543526
rect 89640 539963 89668 543866
rect 90364 543720 90416 543726
rect 90364 543662 90416 543668
rect 90376 539963 90404 543662
rect 91020 539963 91048 543866
rect 91112 543658 91140 560102
rect 93860 559972 93912 559978
rect 93860 559914 93912 559920
rect 92572 555620 92624 555626
rect 92572 555562 92624 555568
rect 91744 547392 91796 547398
rect 91744 547334 91796 547340
rect 91100 543652 91152 543658
rect 91100 543594 91152 543600
rect 91756 539963 91784 547334
rect 92584 540138 92612 555562
rect 93872 547874 93900 559914
rect 94516 558414 94544 560102
rect 97000 560102 97382 560130
rect 98092 560108 98144 560114
rect 96804 560040 96856 560046
rect 96804 559982 96856 559988
rect 94504 558408 94556 558414
rect 94504 558350 94556 558356
rect 93952 558272 94004 558278
rect 93952 558214 94004 558220
rect 93964 551478 93992 558214
rect 93952 551472 94004 551478
rect 93952 551414 94004 551420
rect 96816 547874 96844 559982
rect 97000 552838 97028 560102
rect 99958 560102 100248 560130
rect 98092 560050 98144 560056
rect 98104 557534 98132 560050
rect 100220 558278 100248 560102
rect 102888 560102 103178 560130
rect 104912 560102 105754 560130
rect 106280 560118 106332 560124
rect 102888 558822 102916 560102
rect 100760 558816 100812 558822
rect 100760 558758 100812 558764
rect 102876 558816 102928 558822
rect 102876 558758 102928 558764
rect 100208 558272 100260 558278
rect 100208 558214 100260 558220
rect 98104 557506 98224 557534
rect 96988 552832 97040 552838
rect 96988 552774 97040 552780
rect 93872 547846 93992 547874
rect 96816 547846 97488 547874
rect 93216 543516 93268 543522
rect 93216 543458 93268 543464
rect 92508 540110 92612 540138
rect 92508 539920 92536 540110
rect 93228 539963 93256 543458
rect 93964 539963 93992 547846
rect 94596 544468 94648 544474
rect 94596 544410 94648 544416
rect 94608 539963 94636 544410
rect 96804 543652 96856 543658
rect 96804 543594 96856 543600
rect 96068 543584 96120 543590
rect 96068 543526 96120 543532
rect 95332 543448 95384 543454
rect 95332 543390 95384 543396
rect 95344 539963 95372 543390
rect 96080 539963 96108 543526
rect 96816 539963 96844 543594
rect 97460 539963 97488 547846
rect 98196 539963 98224 557506
rect 100392 555620 100444 555626
rect 100392 555562 100444 555568
rect 99656 543312 99708 543318
rect 99656 543254 99708 543260
rect 98920 543244 98972 543250
rect 98920 543186 98972 543192
rect 98932 539963 98960 543186
rect 99668 539963 99696 543254
rect 100404 539963 100432 555562
rect 100772 543930 100800 558758
rect 104164 558408 104216 558414
rect 104164 558350 104216 558356
rect 103520 552900 103572 552906
rect 103520 552842 103572 552848
rect 102508 551404 102560 551410
rect 102508 551346 102560 551352
rect 101036 550044 101088 550050
rect 101036 549986 101088 549992
rect 100760 543924 100812 543930
rect 100760 543866 100812 543872
rect 101048 539963 101076 549986
rect 101772 543924 101824 543930
rect 101772 543866 101824 543872
rect 101784 539963 101812 543866
rect 102520 539963 102548 551346
rect 103244 545828 103296 545834
rect 103244 545770 103296 545776
rect 103256 539963 103284 545770
rect 103532 543946 103560 552842
rect 104176 544066 104204 558350
rect 104912 548690 104940 560102
rect 104900 548684 104952 548690
rect 104900 548626 104952 548632
rect 105360 547256 105412 547262
rect 105360 547198 105412 547204
rect 104164 544060 104216 544066
rect 104164 544002 104216 544008
rect 103532 543918 104664 543946
rect 103980 543244 104032 543250
rect 103980 543186 104032 543192
rect 103992 539963 104020 543186
rect 104636 539963 104664 543918
rect 105372 539963 105400 547198
rect 106292 543930 106320 560118
rect 108592 560102 108974 560130
rect 110524 560102 111550 560130
rect 114664 560102 114770 560130
rect 117346 560102 117452 560130
rect 108304 558340 108356 558346
rect 108304 558282 108356 558288
rect 106924 552900 106976 552906
rect 106924 552842 106976 552848
rect 106280 543924 106332 543930
rect 106280 543866 106332 543872
rect 106096 543720 106148 543726
rect 106096 543662 106148 543668
rect 106108 539963 106136 543662
rect 106936 543590 106964 552842
rect 108212 548548 108264 548554
rect 108212 548490 108264 548496
rect 107568 543924 107620 543930
rect 107568 543866 107620 543872
rect 106924 543584 106976 543590
rect 106924 543526 106976 543532
rect 106832 543312 106884 543318
rect 106832 543254 106884 543260
rect 106844 539963 106872 543254
rect 107580 539963 107608 543866
rect 108224 539963 108252 548490
rect 108316 543726 108344 558282
rect 108592 554198 108620 560102
rect 108580 554192 108632 554198
rect 108580 554134 108632 554140
rect 110420 554124 110472 554130
rect 110420 554066 110472 554072
rect 109684 550112 109736 550118
rect 109684 550054 109736 550060
rect 108948 544400 109000 544406
rect 108948 544342 109000 544348
rect 108304 543720 108356 543726
rect 108304 543662 108356 543668
rect 108960 539963 108988 544342
rect 109696 539963 109724 550054
rect 110432 543946 110460 554066
rect 110524 547194 110552 560102
rect 112444 558408 112496 558414
rect 112444 558350 112496 558356
rect 111892 558340 111944 558346
rect 111892 558282 111944 558288
rect 111904 547874 111932 558282
rect 112456 548622 112484 558350
rect 114560 558204 114612 558210
rect 114560 558146 114612 558152
rect 112444 548616 112496 548622
rect 112444 548558 112496 548564
rect 111904 547846 112576 547874
rect 110512 547188 110564 547194
rect 110512 547130 110564 547136
rect 110432 543918 111104 543946
rect 110420 543516 110472 543522
rect 110420 543458 110472 543464
rect 110432 539963 110460 543458
rect 111076 539963 111104 543918
rect 111800 543720 111852 543726
rect 111800 543662 111852 543668
rect 111812 539963 111840 543662
rect 112548 539963 112576 547846
rect 113272 544060 113324 544066
rect 113272 544002 113324 544008
rect 113284 539963 113312 544002
rect 114572 543930 114600 558146
rect 114664 552702 114692 560102
rect 116584 558816 116636 558822
rect 116584 558758 116636 558764
rect 115204 558272 115256 558278
rect 115204 558214 115256 558220
rect 114652 552696 114704 552702
rect 114652 552638 114704 552644
rect 114652 551472 114704 551478
rect 114652 551414 114704 551420
rect 114560 543924 114612 543930
rect 114560 543866 114612 543872
rect 114008 543448 114060 543454
rect 114008 543390 114060 543396
rect 114020 539963 114048 543390
rect 114664 539963 114692 551414
rect 115216 543726 115244 558214
rect 116596 545902 116624 558758
rect 117424 558414 117452 560102
rect 120184 560102 120566 560130
rect 120184 558822 120212 560102
rect 120172 558816 120224 558822
rect 120172 558758 120224 558764
rect 120736 558754 120764 622390
rect 120814 598360 120870 598369
rect 120814 598295 120870 598304
rect 119344 558748 119396 558754
rect 119344 558690 119396 558696
rect 120724 558748 120776 558754
rect 120724 558690 120776 558696
rect 117412 558408 117464 558414
rect 117412 558350 117464 558356
rect 118700 558272 118752 558278
rect 118700 558214 118752 558220
rect 116584 545896 116636 545902
rect 116584 545838 116636 545844
rect 115388 543924 115440 543930
rect 115388 543866 115440 543872
rect 115204 543720 115256 543726
rect 115204 543662 115256 543668
rect 115400 539963 115428 543866
rect 116124 543720 116176 543726
rect 116124 543662 116176 543668
rect 116136 539963 116164 543662
rect 118240 543584 118292 543590
rect 118240 543526 118292 543532
rect 116860 543108 116912 543114
rect 116860 543050 116912 543056
rect 116872 539963 116900 543050
rect 117596 543040 117648 543046
rect 117596 542982 117648 542988
rect 117608 539963 117636 542982
rect 118252 539963 118280 543526
rect 118712 543402 118740 558214
rect 119356 543522 119384 558690
rect 120828 552770 120856 598295
rect 120920 559910 120948 625398
rect 122288 625388 122340 625394
rect 122288 625330 122340 625336
rect 121644 625252 121696 625258
rect 121644 625194 121696 625200
rect 121552 622396 121604 622402
rect 121552 622338 121604 622344
rect 120998 576872 121054 576881
rect 120998 576807 121054 576816
rect 120908 559904 120960 559910
rect 120908 559846 120960 559852
rect 120816 552764 120868 552770
rect 120816 552706 120868 552712
rect 120264 550044 120316 550050
rect 120264 549986 120316 549992
rect 120276 543946 120304 549986
rect 121012 549982 121040 576807
rect 121458 571024 121514 571033
rect 121458 570959 121514 570968
rect 121090 564904 121146 564913
rect 121090 564839 121146 564848
rect 121000 549976 121052 549982
rect 121000 549918 121052 549924
rect 121104 544066 121132 564839
rect 121182 562184 121238 562193
rect 121182 562119 121238 562128
rect 121196 554062 121224 562119
rect 121472 556986 121500 570959
rect 121564 559842 121592 622338
rect 121552 559836 121604 559842
rect 121552 559778 121604 559784
rect 121460 556980 121512 556986
rect 121460 556922 121512 556928
rect 121184 554056 121236 554062
rect 121184 553998 121236 554004
rect 121460 552832 121512 552838
rect 121460 552774 121512 552780
rect 121092 544060 121144 544066
rect 121092 544002 121144 544008
rect 121472 543946 121500 552774
rect 121552 551472 121604 551478
rect 121552 551414 121604 551420
rect 121564 544066 121592 551414
rect 121656 547874 121684 625194
rect 121734 613864 121790 613873
rect 121734 613799 121790 613808
rect 121748 559774 121776 613799
rect 121918 611144 121974 611153
rect 121918 611079 121974 611088
rect 121826 601624 121882 601633
rect 121826 601559 121882 601568
rect 121736 559768 121788 559774
rect 121736 559710 121788 559716
rect 121840 549914 121868 601559
rect 121932 559706 121960 611079
rect 122194 586664 122250 586673
rect 122194 586599 122250 586608
rect 122102 583264 122158 583273
rect 122102 583199 122158 583208
rect 122010 580544 122066 580553
rect 122010 580479 122066 580488
rect 121920 559700 121972 559706
rect 121920 559642 121972 559648
rect 121828 549908 121880 549914
rect 121828 549850 121880 549856
rect 121656 547846 121960 547874
rect 121552 544060 121604 544066
rect 121552 544002 121604 544008
rect 120276 543918 121132 543946
rect 121472 543918 121868 543946
rect 119344 543516 119396 543522
rect 119344 543458 119396 543464
rect 120448 543516 120500 543522
rect 120448 543458 120500 543464
rect 118712 543374 119752 543402
rect 118976 543108 119028 543114
rect 118976 543050 119028 543056
rect 118988 539963 119016 543050
rect 119724 539963 119752 543374
rect 120460 539963 120488 543458
rect 121104 539963 121132 543918
rect 121840 539963 121868 543918
rect 121932 543386 121960 547846
rect 122024 547330 122052 580479
rect 122116 551546 122144 583199
rect 122208 555558 122236 586599
rect 122196 555552 122248 555558
rect 122196 555494 122248 555500
rect 122104 551540 122156 551546
rect 122104 551482 122156 551488
rect 122300 547874 122328 625330
rect 122852 560114 122880 625466
rect 124220 625320 124272 625326
rect 124220 625262 124272 625268
rect 122930 619984 122986 619993
rect 122930 619919 122986 619928
rect 122840 560108 122892 560114
rect 122840 560050 122892 560056
rect 122944 559638 122972 619919
rect 123114 617264 123170 617273
rect 123114 617199 123170 617208
rect 123022 607744 123078 607753
rect 123022 607679 123078 607688
rect 122932 559632 122984 559638
rect 122932 559574 122984 559580
rect 122840 557048 122892 557054
rect 122840 556990 122892 556996
rect 122208 547846 122328 547874
rect 122012 547324 122064 547330
rect 122012 547266 122064 547272
rect 121920 543380 121972 543386
rect 121920 543322 121972 543328
rect 122208 542978 122236 547846
rect 122656 547188 122708 547194
rect 122656 547130 122708 547136
rect 122564 544060 122616 544066
rect 122564 544002 122616 544008
rect 122196 542972 122248 542978
rect 122196 542914 122248 542920
rect 122576 539963 122604 544002
rect 122668 543522 122696 547130
rect 122852 543946 122880 556990
rect 122932 554192 122984 554198
rect 122932 554134 122984 554140
rect 122944 544048 122972 554134
rect 123036 545766 123064 607679
rect 123128 558346 123156 617199
rect 123206 605024 123262 605033
rect 123206 604959 123262 604968
rect 123116 558340 123168 558346
rect 123116 558282 123168 558288
rect 123220 551342 123248 604959
rect 123390 595504 123446 595513
rect 123390 595439 123446 595448
rect 123298 592784 123354 592793
rect 123298 592719 123354 592728
rect 123208 551336 123260 551342
rect 123208 551278 123260 551284
rect 123024 545760 123076 545766
rect 123024 545702 123076 545708
rect 123312 544474 123340 592719
rect 123404 552906 123432 595439
rect 124128 589416 124180 589422
rect 124126 589384 124128 589393
rect 124180 589384 124182 589393
rect 124126 589319 124182 589328
rect 123482 574424 123538 574433
rect 123482 574359 123538 574368
rect 123496 555626 123524 574359
rect 123574 568304 123630 568313
rect 123574 568239 123630 568248
rect 123588 556918 123616 568239
rect 123576 556912 123628 556918
rect 123576 556854 123628 556860
rect 123484 555620 123536 555626
rect 123484 555562 123536 555568
rect 123392 552900 123444 552906
rect 123392 552842 123444 552848
rect 123300 544468 123352 544474
rect 123300 544410 123352 544416
rect 122944 544020 124076 544048
rect 122852 543918 123340 543946
rect 122656 543516 122708 543522
rect 122656 543458 122708 543464
rect 123312 539963 123340 543918
rect 124048 539963 124076 544020
rect 124232 543930 124260 625262
rect 124312 623892 124364 623898
rect 124312 623834 124364 623840
rect 124220 543924 124272 543930
rect 124220 543866 124272 543872
rect 124324 543046 124352 623834
rect 124404 623824 124456 623830
rect 124404 623766 124456 623772
rect 124416 543454 124444 623766
rect 124508 560046 124536 625602
rect 124600 560182 124628 625670
rect 124588 560176 124640 560182
rect 124588 560118 124640 560124
rect 124496 560040 124548 560046
rect 124496 559982 124548 559988
rect 124692 559978 124720 625738
rect 137744 625728 137796 625734
rect 137744 625670 137796 625676
rect 125692 625592 125744 625598
rect 125692 625534 125744 625540
rect 135168 625592 135220 625598
rect 135168 625534 135220 625540
rect 125600 576904 125652 576910
rect 125600 576846 125652 576852
rect 124680 559972 124732 559978
rect 124680 559914 124732 559920
rect 124680 547324 124732 547330
rect 124680 547266 124732 547272
rect 124404 543448 124456 543454
rect 124404 543390 124456 543396
rect 124312 543040 124364 543046
rect 124312 542982 124364 542988
rect 124692 539963 124720 547266
rect 125612 543930 125640 576846
rect 125416 543924 125468 543930
rect 125416 543866 125468 543872
rect 125600 543924 125652 543930
rect 125600 543866 125652 543872
rect 125428 539963 125456 543866
rect 125704 543318 125732 625534
rect 134892 625388 134944 625394
rect 134892 625330 134944 625336
rect 133880 625184 133932 625190
rect 133880 625126 133932 625132
rect 133144 623892 133196 623898
rect 133144 623834 133196 623840
rect 126244 622736 126296 622742
rect 126244 622678 126296 622684
rect 126256 543590 126284 622678
rect 132500 607232 132552 607238
rect 132500 607174 132552 607180
rect 129740 558408 129792 558414
rect 129740 558350 129792 558356
rect 129004 552900 129056 552906
rect 129004 552842 129056 552848
rect 127624 545760 127676 545766
rect 127624 545702 127676 545708
rect 126888 543924 126940 543930
rect 126888 543866 126940 543872
rect 126244 543584 126296 543590
rect 126244 543526 126296 543532
rect 125692 543312 125744 543318
rect 125692 543254 125744 543260
rect 126152 543040 126204 543046
rect 126152 542982 126204 542988
rect 126164 539963 126192 542982
rect 126900 539963 126928 543866
rect 127636 539963 127664 545702
rect 128268 543244 128320 543250
rect 128268 543186 128320 543192
rect 128280 539963 128308 543186
rect 129016 539963 129044 552842
rect 129752 543930 129780 558350
rect 129832 554260 129884 554266
rect 129832 554202 129884 554208
rect 129740 543924 129792 543930
rect 129740 543866 129792 543872
rect 129844 540138 129872 554202
rect 131212 544400 131264 544406
rect 131212 544342 131264 544348
rect 130476 543924 130528 543930
rect 130476 543866 130528 543872
rect 129768 540110 129872 540138
rect 129768 539920 129796 540110
rect 130488 539963 130516 543866
rect 131224 539963 131252 544342
rect 132512 543946 132540 607174
rect 132592 558204 132644 558210
rect 132592 558146 132644 558152
rect 132604 557534 132632 558146
rect 132604 557506 132908 557534
rect 132512 543918 132632 543946
rect 131856 543584 131908 543590
rect 131856 543526 131908 543532
rect 131868 539963 131896 543526
rect 132604 539963 132632 543918
rect 132880 543402 132908 557506
rect 133156 543590 133184 623834
rect 133892 543946 133920 625126
rect 134616 589416 134668 589422
rect 134616 589358 134668 589364
rect 134524 589348 134576 589354
rect 134524 589290 134576 589296
rect 133972 558340 134024 558346
rect 133972 558282 134024 558288
rect 133984 557534 134012 558282
rect 133984 557506 134472 557534
rect 133892 543918 134104 543946
rect 133144 543584 133196 543590
rect 133144 543526 133196 543532
rect 132880 543374 133368 543402
rect 133340 539963 133368 543374
rect 134076 539963 134104 543918
rect 134444 542994 134472 557506
rect 134536 543114 134564 589290
rect 134628 560182 134656 589358
rect 134616 560176 134668 560182
rect 134616 560118 134668 560124
rect 134904 559774 134932 625330
rect 135076 622804 135128 622810
rect 135076 622746 135128 622752
rect 134984 622532 135036 622538
rect 134984 622474 135036 622480
rect 134892 559768 134944 559774
rect 134892 559710 134944 559716
rect 134996 543658 135024 622474
rect 134984 543652 135036 543658
rect 134984 543594 135036 543600
rect 135088 543454 135116 622746
rect 135180 543590 135208 625534
rect 136364 625524 136416 625530
rect 136364 625466 136416 625472
rect 135260 625252 135312 625258
rect 135260 625194 135312 625200
rect 135272 557534 135300 625194
rect 136376 559706 136404 625466
rect 136640 623824 136692 623830
rect 136640 623766 136692 623772
rect 136456 622668 136508 622674
rect 136456 622610 136508 622616
rect 136364 559700 136416 559706
rect 136364 559642 136416 559648
rect 135272 557506 136220 557534
rect 135444 543720 135496 543726
rect 135444 543662 135496 543668
rect 135168 543584 135220 543590
rect 135168 543526 135220 543532
rect 135076 543448 135128 543454
rect 135076 543390 135128 543396
rect 134524 543108 134576 543114
rect 134524 543050 134576 543056
rect 134444 542966 134748 542994
rect 134720 539963 134748 542966
rect 135456 539963 135484 543662
rect 136192 539963 136220 557506
rect 136468 543182 136496 622610
rect 136548 622600 136600 622606
rect 136548 622542 136600 622548
rect 136560 543522 136588 622542
rect 136652 543930 136680 623766
rect 137374 620664 137430 620673
rect 137374 620599 137430 620608
rect 136730 608288 136786 608297
rect 136730 608223 136786 608232
rect 136744 607238 136772 608223
rect 136732 607232 136784 607238
rect 136732 607174 136784 607180
rect 137282 594824 137338 594833
rect 137282 594759 137338 594768
rect 136730 589928 136786 589937
rect 136730 589863 136786 589872
rect 136744 589354 136772 589863
rect 136732 589348 136784 589354
rect 136732 589290 136784 589296
rect 136730 577688 136786 577697
rect 136730 577623 136786 577632
rect 136744 576910 136772 577623
rect 136732 576904 136784 576910
rect 136732 576846 136784 576852
rect 137296 561202 137324 594759
rect 137284 561196 137336 561202
rect 137284 561138 137336 561144
rect 136916 548548 136968 548554
rect 136916 548490 136968 548496
rect 136640 543924 136692 543930
rect 136640 543866 136692 543872
rect 136548 543516 136600 543522
rect 136548 543458 136600 543464
rect 136456 543176 136508 543182
rect 136456 543118 136508 543124
rect 136928 539963 136956 548490
rect 137388 543726 137416 620599
rect 137650 611688 137706 611697
rect 137650 611623 137706 611632
rect 137466 574968 137522 574977
rect 137466 574903 137522 574912
rect 137480 547194 137508 574903
rect 137558 571568 137614 571577
rect 137558 571503 137614 571512
rect 137468 547188 137520 547194
rect 137468 547130 137520 547136
rect 137572 543862 137600 571503
rect 137664 560250 137692 611623
rect 137652 560244 137704 560250
rect 137652 560186 137704 560192
rect 137756 559910 137784 625670
rect 137848 599593 137876 683130
rect 169772 635526 169800 702406
rect 235184 700398 235212 703520
rect 235172 700392 235224 700398
rect 235172 700334 235224 700340
rect 299492 641034 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 305644 700392 305696 700398
rect 305644 700334 305696 700340
rect 299480 641028 299532 641034
rect 299480 640970 299532 640976
rect 169760 635520 169812 635526
rect 169760 635462 169812 635468
rect 298100 633684 298152 633690
rect 298100 633626 298152 633632
rect 289820 633616 289872 633622
rect 289820 633558 289872 633564
rect 288440 633480 288492 633486
rect 288440 633422 288492 633428
rect 281078 632224 281134 632233
rect 281078 632159 281134 632168
rect 218704 630692 218756 630698
rect 218704 630634 218756 630640
rect 217784 629944 217836 629950
rect 217784 629886 217836 629892
rect 213920 625796 213972 625802
rect 213920 625738 213972 625744
rect 186504 625728 186556 625734
rect 186504 625670 186556 625676
rect 206468 625728 206520 625734
rect 206468 625670 206520 625676
rect 139308 625660 139360 625666
rect 139308 625602 139360 625608
rect 162860 625660 162912 625666
rect 162860 625602 162912 625608
rect 139124 625456 139176 625462
rect 139124 625398 139176 625404
rect 137928 622464 137980 622470
rect 137928 622406 137980 622412
rect 137834 599584 137890 599593
rect 137834 599519 137890 599528
rect 137940 596193 137968 622406
rect 139030 617808 139086 617817
rect 139030 617743 139086 617752
rect 138846 605568 138902 605577
rect 138846 605503 138902 605512
rect 137926 596184 137982 596193
rect 137926 596119 137982 596128
rect 137940 594833 137968 596119
rect 137926 594824 137982 594833
rect 137926 594759 137982 594768
rect 137926 593464 137982 593473
rect 137926 593399 137982 593408
rect 137834 583808 137890 583817
rect 137834 583743 137890 583752
rect 137744 559904 137796 559910
rect 137744 559846 137796 559852
rect 137848 555626 137876 583743
rect 137836 555620 137888 555626
rect 137836 555562 137888 555568
rect 137940 544474 137968 593399
rect 138754 587208 138810 587217
rect 138754 587143 138810 587152
rect 138662 581088 138718 581097
rect 138662 581023 138718 581032
rect 138570 568848 138626 568857
rect 138570 568783 138626 568792
rect 138478 565448 138534 565457
rect 138478 565383 138534 565392
rect 138492 552770 138520 565383
rect 138584 555558 138612 568783
rect 138572 555552 138624 555558
rect 138572 555494 138624 555500
rect 138480 552764 138532 552770
rect 138480 552706 138532 552712
rect 138676 552702 138704 581023
rect 138664 552696 138716 552702
rect 138664 552638 138716 552644
rect 138768 549982 138796 587143
rect 138860 559638 138888 605503
rect 138938 602168 138994 602177
rect 138938 602103 138994 602112
rect 138848 559632 138900 559638
rect 138848 559574 138900 559580
rect 138952 556918 138980 602103
rect 139044 559842 139072 617743
rect 139032 559836 139084 559842
rect 139032 559778 139084 559784
rect 139136 558958 139164 625398
rect 139214 614408 139270 614417
rect 139214 614343 139270 614352
rect 139124 558952 139176 558958
rect 139124 558894 139176 558900
rect 138940 556912 138992 556918
rect 138940 556854 138992 556860
rect 138756 549976 138808 549982
rect 138756 549918 138808 549924
rect 138296 545964 138348 545970
rect 138296 545906 138348 545912
rect 137928 544468 137980 544474
rect 137928 544410 137980 544416
rect 137652 543924 137704 543930
rect 137652 543866 137704 543872
rect 137560 543856 137612 543862
rect 137560 543798 137612 543804
rect 137376 543720 137428 543726
rect 137376 543662 137428 543668
rect 137664 539963 137692 543866
rect 138308 539963 138336 545906
rect 139032 545896 139084 545902
rect 139032 545838 139084 545844
rect 139044 539963 139072 545838
rect 139228 543318 139256 614343
rect 139320 543386 139348 625602
rect 160284 625592 160336 625598
rect 160284 625534 160336 625540
rect 139860 625184 139912 625190
rect 139860 625126 139912 625132
rect 157524 625184 157576 625190
rect 157524 625126 157576 625132
rect 139398 562796 139454 562805
rect 139398 562731 139454 562740
rect 139412 551342 139440 562731
rect 139400 551336 139452 551342
rect 139400 551278 139452 551284
rect 139872 546514 139900 625126
rect 140136 625116 140188 625122
rect 140136 625058 140188 625064
rect 140148 623098 140176 625058
rect 151268 623892 151320 623898
rect 151268 623834 151320 623840
rect 140070 623070 140176 623098
rect 151280 623098 151308 623834
rect 157536 623098 157564 625126
rect 151280 623070 151662 623098
rect 157458 623070 157564 623098
rect 160296 623098 160324 625534
rect 162872 623098 162900 625602
rect 166172 625524 166224 625530
rect 166172 625466 166224 625472
rect 166184 623098 166212 625466
rect 174452 625456 174504 625462
rect 174452 625398 174504 625404
rect 171876 625320 171928 625326
rect 171876 625262 171928 625268
rect 168748 623824 168800 623830
rect 168748 623766 168800 623772
rect 168760 623098 168788 623766
rect 171888 623098 171916 625262
rect 174464 623098 174492 625398
rect 180340 625388 180392 625394
rect 180340 625330 180392 625336
rect 180352 623098 180380 625330
rect 183652 625252 183704 625258
rect 183652 625194 183704 625200
rect 183664 623098 183692 625194
rect 160296 623070 160678 623098
rect 162872 623070 163254 623098
rect 166184 623070 166474 623098
rect 168760 623070 169050 623098
rect 171888 623070 172270 623098
rect 174464 623070 174846 623098
rect 180352 623070 180642 623098
rect 183664 623070 183862 623098
rect 186516 622962 186544 625670
rect 190000 625388 190052 625394
rect 190000 625330 190052 625336
rect 204444 625388 204496 625394
rect 204444 625330 204496 625336
rect 190012 623098 190040 625330
rect 192576 625252 192628 625258
rect 192576 625194 192628 625200
rect 201684 625252 201736 625258
rect 201684 625194 201736 625200
rect 192588 623098 192616 625194
rect 195704 625184 195756 625190
rect 195704 625126 195756 625132
rect 200856 625184 200908 625190
rect 200856 625126 200908 625132
rect 195716 623098 195744 625126
rect 189658 623070 190040 623098
rect 192234 623070 192616 623098
rect 195454 623070 195744 623098
rect 186438 622934 186544 622962
rect 145576 622810 145866 622826
rect 145564 622804 145866 622810
rect 145616 622798 145866 622804
rect 145564 622746 145616 622752
rect 177856 622736 177908 622742
rect 149086 622674 149192 622690
rect 177908 622684 178066 622690
rect 177856 622678 178066 622684
rect 149086 622668 149204 622674
rect 149086 622662 149152 622668
rect 177868 622662 178066 622678
rect 149152 622610 149204 622616
rect 154580 622600 154632 622606
rect 143000 622538 143290 622554
rect 154632 622548 154882 622554
rect 154580 622542 154882 622548
rect 142988 622532 143290 622538
rect 143040 622526 143290 622532
rect 154592 622526 154882 622542
rect 142988 622474 143040 622480
rect 198030 622402 198320 622418
rect 198030 622396 198332 622402
rect 198030 622390 198280 622396
rect 200606 622390 200712 622418
rect 198280 622338 198332 622344
rect 140780 560244 140832 560250
rect 140780 560186 140832 560192
rect 159836 560238 160034 560266
rect 165632 560238 165830 560266
rect 194612 560238 194810 560266
rect 140070 560102 140360 560130
rect 140332 558482 140360 560102
rect 140320 558476 140372 558482
rect 140320 558418 140372 558424
rect 140792 557534 140820 560186
rect 142646 560102 142936 560130
rect 142160 558952 142212 558958
rect 142160 558894 142212 558900
rect 140792 557506 141280 557534
rect 140504 547392 140556 547398
rect 140504 547334 140556 547340
rect 139860 546508 139912 546514
rect 139860 546450 139912 546456
rect 139768 543856 139820 543862
rect 139768 543798 139820 543804
rect 139308 543380 139360 543386
rect 139308 543322 139360 543328
rect 139216 543312 139268 543318
rect 139216 543254 139268 543260
rect 139780 539963 139808 543798
rect 140516 539963 140544 547334
rect 141252 539963 141280 557506
rect 141884 546508 141936 546514
rect 141884 546450 141936 546456
rect 141896 539963 141924 546450
rect 142172 543930 142200 558894
rect 142908 558550 142936 560102
rect 144932 560102 145222 560130
rect 147784 560102 148442 560130
rect 151018 560102 151400 560130
rect 142896 558544 142948 558550
rect 142896 558486 142948 558492
rect 144932 558278 144960 560102
rect 145104 559904 145156 559910
rect 145104 559846 145156 559852
rect 144920 558272 144972 558278
rect 144920 558214 144972 558220
rect 145116 557534 145144 559846
rect 147680 558680 147732 558686
rect 147680 558622 147732 558628
rect 145116 557506 145512 557534
rect 143540 556980 143592 556986
rect 143540 556922 143592 556928
rect 142620 550112 142672 550118
rect 142620 550054 142672 550060
rect 142160 543924 142212 543930
rect 142160 543866 142212 543872
rect 142632 539963 142660 550054
rect 143552 543930 143580 556922
rect 144092 551540 144144 551546
rect 144092 551482 144144 551488
rect 143356 543924 143408 543930
rect 143356 543866 143408 543872
rect 143540 543924 143592 543930
rect 143540 543866 143592 543872
rect 143368 539963 143396 543866
rect 144104 539963 144132 551482
rect 144736 543924 144788 543930
rect 144736 543866 144788 543872
rect 144748 539963 144776 543866
rect 145484 539963 145512 557506
rect 147692 547874 147720 558622
rect 147784 549914 147812 560102
rect 150624 559836 150676 559842
rect 150624 559778 150676 559784
rect 149060 555620 149112 555626
rect 149060 555562 149112 555568
rect 147772 549908 147824 549914
rect 147772 549850 147824 549856
rect 147692 547846 148364 547874
rect 147680 547188 147732 547194
rect 147680 547130 147732 547136
rect 146208 543720 146260 543726
rect 146208 543662 146260 543668
rect 146220 539963 146248 543662
rect 146944 543652 146996 543658
rect 146944 543594 146996 543600
rect 146956 539963 146984 543594
rect 147692 539963 147720 547130
rect 148336 539963 148364 547846
rect 149072 539963 149100 555562
rect 149796 544468 149848 544474
rect 149796 544410 149848 544416
rect 149808 539963 149836 544410
rect 150636 540138 150664 559778
rect 151372 558618 151400 560102
rect 153856 560102 154238 560130
rect 156432 560102 156814 560130
rect 151820 559768 151872 559774
rect 151820 559710 151872 559716
rect 151360 558612 151412 558618
rect 151360 558554 151412 558560
rect 151832 557534 151860 559710
rect 153856 558414 153884 560102
rect 154580 559836 154632 559842
rect 154580 559778 154632 559784
rect 153844 558408 153896 558414
rect 153844 558350 153896 558356
rect 151832 557506 151952 557534
rect 151268 543584 151320 543590
rect 151268 543526 151320 543532
rect 150560 540110 150664 540138
rect 150560 539920 150588 540110
rect 151280 539963 151308 543526
rect 151924 539963 151952 557506
rect 153384 549976 153436 549982
rect 153384 549918 153436 549924
rect 152648 544468 152700 544474
rect 152648 544410 152700 544416
rect 152660 539963 152688 544410
rect 153396 539963 153424 549918
rect 154592 544814 154620 559778
rect 156052 559768 156104 559774
rect 156052 559710 156104 559716
rect 154672 558408 154724 558414
rect 154672 558350 154724 558356
rect 154684 557534 154712 558350
rect 156064 557534 156092 559710
rect 154684 557506 154896 557534
rect 156064 557506 156276 557534
rect 154580 544808 154632 544814
rect 154580 544750 154632 544756
rect 154120 542428 154172 542434
rect 154120 542370 154172 542376
rect 154132 539963 154160 542370
rect 154868 539963 154896 557506
rect 155500 544808 155552 544814
rect 155500 544750 155552 544756
rect 155512 539963 155540 544750
rect 156248 539963 156276 557506
rect 156432 556986 156460 560102
rect 157984 559904 158036 559910
rect 157984 559846 158036 559852
rect 156420 556980 156472 556986
rect 156420 556922 156472 556928
rect 157892 555620 157944 555626
rect 157892 555562 157944 555568
rect 157708 543516 157760 543522
rect 157708 543458 157760 543464
rect 156972 543448 157024 543454
rect 156972 543390 157024 543396
rect 156984 539963 157012 543390
rect 157720 539963 157748 543458
rect 157904 543130 157932 555562
rect 157996 543250 158024 559846
rect 159364 558476 159416 558482
rect 159364 558418 159416 558424
rect 158720 558272 158772 558278
rect 158720 558214 158772 558220
rect 158732 543930 158760 558214
rect 159088 551336 159140 551342
rect 159088 551278 159140 551284
rect 158720 543924 158772 543930
rect 158720 543866 158772 543872
rect 157984 543244 158036 543250
rect 157984 543186 158036 543192
rect 157904 543102 158392 543130
rect 158364 539963 158392 543102
rect 159100 539963 159128 551278
rect 159376 543658 159404 558418
rect 159836 556986 159864 560238
rect 162320 560102 162610 560130
rect 161664 559700 161716 559706
rect 161664 559642 161716 559648
rect 161572 558816 161624 558822
rect 161572 558758 161624 558764
rect 160744 558544 160796 558550
rect 160744 558486 160796 558492
rect 159824 556980 159876 556986
rect 159824 556922 159876 556928
rect 160100 556912 160152 556918
rect 160100 556854 160152 556860
rect 160112 543946 160140 556854
rect 160652 552764 160704 552770
rect 160652 552706 160704 552712
rect 159824 543924 159876 543930
rect 160112 543918 160600 543946
rect 159824 543866 159876 543872
rect 159364 543652 159416 543658
rect 159364 543594 159416 543600
rect 159836 539963 159864 543866
rect 160572 539963 160600 543918
rect 160664 543130 160692 552706
rect 160756 543250 160784 558486
rect 161388 544536 161440 544542
rect 161388 544478 161440 544484
rect 160744 543244 160796 543250
rect 160744 543186 160796 543192
rect 160664 543102 161336 543130
rect 161308 539963 161336 543102
rect 161400 542434 161428 544478
rect 161584 543930 161612 558758
rect 161676 557534 161704 559642
rect 162320 558686 162348 560102
rect 164332 560040 164384 560046
rect 164332 559982 164384 559988
rect 162308 558680 162360 558686
rect 162308 558622 162360 558628
rect 161676 557506 161980 557534
rect 161572 543924 161624 543930
rect 161572 543866 161624 543872
rect 161388 542428 161440 542434
rect 161388 542370 161440 542376
rect 161952 539963 161980 557506
rect 164344 543930 164372 559982
rect 165632 559722 165660 560238
rect 168406 560102 168512 560130
rect 165632 559694 165752 559722
rect 165620 559632 165672 559638
rect 165620 559574 165672 559580
rect 164884 558612 164936 558618
rect 164884 558554 164936 558560
rect 162676 543924 162728 543930
rect 162676 543866 162728 543872
rect 164332 543924 164384 543930
rect 164332 543866 164384 543872
rect 162688 539963 162716 543866
rect 163412 543652 163464 543658
rect 163412 543594 163464 543600
rect 163424 539963 163452 543594
rect 164896 543590 164924 558554
rect 165528 543924 165580 543930
rect 165528 543866 165580 543872
rect 164884 543584 164936 543590
rect 164884 543526 164936 543532
rect 164148 543448 164200 543454
rect 164148 543390 164200 543396
rect 164160 539963 164188 543390
rect 164884 543380 164936 543386
rect 164884 543322 164936 543328
rect 164896 539963 164924 543322
rect 165540 539963 165568 543866
rect 165632 543538 165660 559574
rect 165724 543658 165752 559694
rect 168484 558822 168512 560102
rect 171336 560102 171626 560130
rect 174004 560102 174202 560130
rect 177040 560102 177422 560130
rect 179616 560102 179998 560130
rect 182928 560102 183218 560130
rect 185504 560102 185794 560130
rect 188632 560102 189014 560130
rect 190564 560102 191590 560130
rect 168472 558816 168524 558822
rect 168472 558758 168524 558764
rect 171336 558414 171364 560102
rect 173900 558816 173952 558822
rect 173900 558758 173952 558764
rect 171324 558408 171376 558414
rect 171324 558350 171376 558356
rect 173440 556980 173492 556986
rect 173440 556922 173492 556928
rect 168380 555688 168432 555694
rect 168380 555630 168432 555636
rect 167092 549908 167144 549914
rect 167092 549850 167144 549856
rect 165712 543652 165764 543658
rect 165712 543594 165764 543600
rect 165632 543510 166304 543538
rect 166276 539963 166304 543510
rect 167104 540138 167132 549850
rect 167736 543244 167788 543250
rect 167736 543186 167788 543192
rect 167028 540110 167132 540138
rect 167028 539920 167056 540110
rect 167748 539963 167776 543186
rect 168392 539963 168420 555630
rect 169116 555552 169168 555558
rect 169116 555494 169168 555500
rect 169128 539963 169156 555494
rect 171324 544604 171376 544610
rect 171324 544546 171376 544552
rect 169852 543652 169904 543658
rect 169852 543594 169904 543600
rect 169864 539963 169892 543594
rect 170588 543244 170640 543250
rect 170588 543186 170640 543192
rect 170600 539963 170628 543186
rect 171336 539963 171364 544546
rect 172704 543584 172756 543590
rect 172704 543526 172756 543532
rect 171968 543176 172020 543182
rect 171968 543118 172020 543124
rect 171980 539963 172008 543118
rect 172716 539963 172744 543526
rect 173452 539963 173480 556922
rect 173912 543266 173940 558758
rect 174004 543454 174032 560102
rect 177040 558210 177068 560102
rect 179616 558822 179644 560102
rect 182364 559972 182416 559978
rect 182364 559914 182416 559920
rect 179696 559700 179748 559706
rect 179696 559642 179748 559648
rect 179604 558816 179656 558822
rect 179604 558758 179656 558764
rect 177028 558204 177080 558210
rect 177028 558146 177080 558152
rect 177304 558204 177356 558210
rect 177304 558146 177356 558152
rect 174912 552696 174964 552702
rect 174912 552638 174964 552644
rect 173992 543448 174044 543454
rect 173992 543390 174044 543396
rect 173912 543238 174216 543266
rect 174188 539963 174216 543238
rect 174924 539963 174952 552638
rect 176660 551608 176712 551614
rect 176660 551550 176712 551556
rect 176672 543946 176700 551550
rect 176752 550180 176804 550186
rect 176752 550122 176804 550128
rect 176764 544082 176792 550122
rect 177316 544406 177344 558146
rect 179708 557534 179736 559642
rect 180800 559632 180852 559638
rect 180800 559574 180852 559580
rect 179708 557506 179920 557534
rect 178040 557116 178092 557122
rect 178040 557058 178092 557064
rect 177304 544400 177356 544406
rect 177304 544342 177356 544348
rect 176764 544054 177804 544082
rect 176672 543918 177068 543946
rect 175556 543312 175608 543318
rect 175556 543254 175608 543260
rect 175568 539963 175596 543254
rect 176292 543176 176344 543182
rect 176292 543118 176344 543124
rect 176304 539963 176332 543118
rect 177040 539963 177068 543918
rect 177776 539963 177804 544054
rect 178052 543946 178080 557058
rect 179512 556912 179564 556918
rect 179512 556854 179564 556860
rect 179144 552696 179196 552702
rect 179144 552638 179196 552644
rect 178052 543918 178540 543946
rect 178512 539963 178540 543918
rect 179156 539963 179184 552638
rect 179524 543930 179552 556854
rect 179512 543924 179564 543930
rect 179512 543866 179564 543872
rect 179892 539963 179920 557506
rect 180812 543930 180840 559574
rect 182376 557534 182404 559914
rect 182928 558278 182956 560102
rect 182916 558272 182968 558278
rect 182916 558214 182968 558220
rect 185504 557938 185532 560102
rect 188344 558476 188396 558482
rect 188344 558418 188396 558424
rect 187884 558408 187936 558414
rect 187884 558350 187936 558356
rect 184204 557932 184256 557938
rect 184204 557874 184256 557880
rect 185492 557932 185544 557938
rect 185492 557874 185544 557880
rect 182376 557506 183508 557534
rect 181352 555552 181404 555558
rect 181352 555494 181404 555500
rect 180616 543924 180668 543930
rect 180616 543866 180668 543872
rect 180800 543924 180852 543930
rect 180800 543866 180852 543872
rect 180628 539963 180656 543866
rect 181364 539963 181392 555494
rect 182272 554056 182324 554062
rect 182272 553998 182324 554004
rect 181996 543924 182048 543930
rect 182284 543912 182312 553998
rect 182284 543884 182772 543912
rect 181996 543866 182048 543872
rect 182008 539963 182036 543866
rect 182744 539963 182772 543884
rect 183480 539963 183508 557506
rect 184216 547194 184244 557874
rect 186320 551336 186372 551342
rect 186320 551278 186372 551284
rect 185584 547256 185636 547262
rect 185584 547198 185636 547204
rect 184204 547188 184256 547194
rect 184204 547130 184256 547136
rect 184940 546032 184992 546038
rect 184940 545974 184992 545980
rect 184204 544400 184256 544406
rect 184204 544342 184256 544348
rect 184216 539963 184244 544342
rect 184952 539963 184980 545974
rect 185596 539963 185624 547198
rect 186332 539963 186360 551278
rect 187056 549908 187108 549914
rect 187056 549850 187108 549856
rect 187068 539963 187096 549850
rect 187792 547188 187844 547194
rect 187792 547130 187844 547136
rect 187804 539963 187832 547130
rect 187896 543912 187924 558350
rect 188356 547398 188384 558418
rect 188632 558210 188660 560102
rect 190460 558272 190512 558278
rect 190460 558214 190512 558220
rect 188620 558204 188672 558210
rect 188620 558146 188672 558152
rect 189080 549976 189132 549982
rect 189080 549918 189132 549924
rect 188344 547392 188396 547398
rect 188344 547334 188396 547340
rect 189092 543912 189120 549918
rect 189908 548684 189960 548690
rect 189908 548626 189960 548632
rect 187896 543884 188568 543912
rect 189092 543884 189212 543912
rect 188540 539963 188568 543884
rect 189184 539963 189212 543884
rect 189920 539963 189948 548626
rect 190472 547874 190500 558214
rect 190564 550050 190592 560102
rect 191840 558204 191892 558210
rect 191840 558146 191892 558152
rect 190552 550044 190604 550050
rect 190552 549986 190604 549992
rect 190472 547846 191420 547874
rect 190644 547392 190696 547398
rect 190644 547334 190696 547340
rect 190656 539963 190684 547334
rect 191392 539963 191420 547846
rect 191852 543930 191880 558146
rect 194612 557534 194640 560238
rect 197386 560102 197492 560130
rect 197464 558346 197492 560102
rect 200224 560102 200606 560130
rect 200224 558482 200252 560102
rect 200212 558476 200264 558482
rect 200212 558418 200264 558424
rect 197452 558340 197504 558346
rect 197452 558282 197504 558288
rect 194612 557506 194732 557534
rect 194600 556980 194652 556986
rect 194600 556922 194652 556928
rect 193220 555756 193272 555762
rect 193220 555698 193272 555704
rect 192116 551676 192168 551682
rect 192116 551618 192168 551624
rect 191840 543924 191892 543930
rect 191840 543866 191892 543872
rect 192128 539963 192156 551618
rect 193232 543930 193260 555698
rect 193496 550044 193548 550050
rect 193496 549986 193548 549992
rect 192760 543924 192812 543930
rect 192760 543866 192812 543872
rect 193220 543924 193272 543930
rect 193220 543866 193272 543872
rect 192772 539963 192800 543866
rect 193508 539963 193536 549986
rect 194612 543946 194640 556922
rect 194704 545766 194732 557506
rect 200684 555694 200712 622390
rect 200762 598360 200818 598369
rect 200762 598295 200818 598304
rect 200672 555688 200724 555694
rect 200672 555630 200724 555636
rect 195980 554124 196032 554130
rect 195980 554066 196032 554072
rect 194692 545760 194744 545766
rect 194692 545702 194744 545708
rect 194232 543924 194284 543930
rect 194612 543918 195008 543946
rect 195992 543930 196020 554066
rect 196348 552764 196400 552770
rect 196348 552706 196400 552712
rect 194232 543866 194284 543872
rect 194244 539963 194272 543866
rect 194980 539963 195008 543918
rect 195980 543924 196032 543930
rect 195980 543866 196032 543872
rect 195612 543312 195664 543318
rect 195612 543254 195664 543260
rect 195624 539963 195652 543254
rect 196360 539963 196388 552706
rect 200672 551404 200724 551410
rect 200672 551346 200724 551352
rect 199200 548752 199252 548758
rect 199200 548694 199252 548700
rect 198556 545828 198608 545834
rect 198556 545770 198608 545776
rect 197820 545760 197872 545766
rect 197820 545702 197872 545708
rect 197084 543924 197136 543930
rect 197084 543866 197136 543872
rect 197096 539963 197124 543866
rect 197832 539963 197860 545702
rect 198568 539963 198596 545770
rect 199212 539963 199240 548694
rect 199936 543380 199988 543386
rect 199936 543322 199988 543328
rect 199948 539963 199976 543322
rect 200684 539963 200712 551346
rect 200776 545970 200804 598295
rect 200868 560046 200896 625126
rect 201590 619984 201646 619993
rect 201590 619919 201646 619928
rect 200948 598052 201000 598058
rect 200948 597994 201000 598000
rect 200856 560040 200908 560046
rect 200856 559982 200908 559988
rect 200764 545964 200816 545970
rect 200764 545906 200816 545912
rect 200960 543046 200988 597994
rect 201498 571024 201554 571033
rect 201498 570959 201554 570968
rect 201130 568304 201186 568313
rect 201130 568239 201186 568248
rect 201040 560516 201092 560522
rect 201040 560458 201092 560464
rect 201052 543250 201080 560458
rect 201144 552838 201172 568239
rect 201222 562184 201278 562193
rect 201222 562119 201278 562128
rect 201132 552832 201184 552838
rect 201132 552774 201184 552780
rect 201236 547330 201264 562119
rect 201512 548554 201540 570959
rect 201604 551478 201632 619919
rect 201696 559842 201724 625194
rect 204260 623824 204312 623830
rect 204260 623766 204312 623772
rect 202236 622396 202288 622402
rect 202236 622338 202288 622344
rect 201774 613864 201830 613873
rect 201774 613799 201830 613808
rect 201684 559836 201736 559842
rect 201684 559778 201736 559784
rect 201788 551546 201816 613799
rect 201866 605024 201922 605033
rect 201866 604959 201922 604968
rect 201880 554198 201908 604959
rect 201958 592784 202014 592793
rect 201958 592719 202014 592728
rect 201868 554192 201920 554198
rect 201868 554134 201920 554140
rect 201776 551540 201828 551546
rect 201776 551482 201828 551488
rect 201592 551472 201644 551478
rect 201592 551414 201644 551420
rect 201500 548548 201552 548554
rect 201500 548490 201552 548496
rect 201224 547324 201276 547330
rect 201224 547266 201276 547272
rect 201972 544474 202000 592719
rect 202142 586664 202198 586673
rect 202142 586599 202198 586608
rect 202050 583264 202106 583273
rect 202050 583199 202106 583208
rect 202064 545902 202092 583199
rect 202156 557054 202184 586599
rect 202144 557048 202196 557054
rect 202144 556990 202196 556996
rect 202052 545896 202104 545902
rect 202052 545838 202104 545844
rect 201960 544468 202012 544474
rect 201960 544410 202012 544416
rect 201408 543720 201460 543726
rect 201408 543662 201460 543668
rect 201040 543244 201092 543250
rect 201040 543186 201092 543192
rect 200948 543040 201000 543046
rect 200948 542982 201000 542988
rect 201420 539963 201448 543662
rect 202248 543658 202276 622338
rect 202878 617264 202934 617273
rect 202878 617199 202934 617208
rect 202326 580544 202382 580553
rect 202326 580479 202382 580488
rect 202340 550118 202368 580479
rect 202892 560522 202920 617199
rect 203062 611144 203118 611153
rect 203062 611079 203118 611088
rect 202970 607744 203026 607753
rect 202970 607679 203026 607688
rect 202880 560516 202932 560522
rect 202880 560458 202932 560464
rect 202984 554266 203012 607679
rect 203076 598058 203104 611079
rect 203154 601624 203210 601633
rect 203154 601559 203210 601568
rect 203064 598052 203116 598058
rect 203064 597994 203116 598000
rect 203062 595504 203118 595513
rect 203062 595439 203118 595448
rect 202972 554260 203024 554266
rect 202972 554202 203024 554208
rect 202328 550112 202380 550118
rect 202328 550054 202380 550060
rect 203076 544542 203104 595439
rect 203168 552906 203196 601559
rect 203246 589384 203302 589393
rect 203246 589319 203248 589328
rect 203300 589319 203302 589328
rect 203248 589290 203300 589296
rect 203338 577144 203394 577153
rect 203338 577079 203394 577088
rect 203246 574424 203302 574433
rect 203246 574359 203302 574368
rect 203260 555626 203288 574359
rect 203352 559910 203380 577079
rect 203430 564904 203486 564913
rect 203430 564839 203486 564848
rect 203340 559904 203392 559910
rect 203340 559846 203392 559852
rect 203248 555620 203300 555626
rect 203248 555562 203300 555568
rect 203156 552900 203208 552906
rect 203156 552842 203208 552848
rect 203444 544610 203472 564839
rect 203432 544604 203484 544610
rect 203432 544546 203484 544552
rect 203064 544536 203116 544542
rect 203064 544478 203116 544484
rect 202236 543652 202288 543658
rect 202236 543594 202288 543600
rect 203524 543652 203576 543658
rect 203524 543594 203576 543600
rect 202144 543244 202196 543250
rect 202144 543186 202196 543192
rect 202156 539963 202184 543186
rect 202788 543108 202840 543114
rect 202788 543050 202840 543056
rect 202800 539963 202828 543050
rect 203536 539963 203564 543594
rect 204272 539963 204300 623766
rect 204352 622736 204404 622742
rect 204352 622678 204404 622684
rect 204364 543946 204392 622678
rect 204456 559774 204484 625330
rect 206284 623892 206336 623898
rect 206284 623834 206336 623840
rect 204904 607232 204956 607238
rect 204904 607174 204956 607180
rect 204536 589348 204588 589354
rect 204536 589290 204588 589296
rect 204548 560250 204576 589290
rect 204536 560244 204588 560250
rect 204536 560186 204588 560192
rect 204444 559768 204496 559774
rect 204444 559710 204496 559716
rect 204916 547398 204944 607174
rect 205640 548616 205692 548622
rect 205640 548558 205692 548564
rect 204904 547392 204956 547398
rect 204904 547334 204956 547340
rect 204364 543918 205036 543946
rect 205008 539963 205036 543918
rect 205652 539963 205680 548558
rect 206296 543726 206324 623834
rect 206376 622600 206428 622606
rect 206376 622542 206428 622548
rect 206388 547874 206416 622542
rect 206480 548690 206508 625670
rect 212540 625660 212592 625666
rect 212540 625602 212592 625608
rect 209780 625388 209832 625394
rect 209780 625330 209832 625336
rect 208400 622668 208452 622674
rect 208400 622610 208452 622616
rect 207020 593428 207072 593434
rect 207020 593370 207072 593376
rect 206560 574116 206612 574122
rect 206560 574058 206612 574064
rect 206572 557122 206600 574058
rect 207032 557534 207060 593370
rect 207032 557506 207888 557534
rect 206560 557116 206612 557122
rect 206560 557058 206612 557064
rect 206468 548684 206520 548690
rect 206468 548626 206520 548632
rect 206388 547846 206508 547874
rect 206376 545964 206428 545970
rect 206376 545906 206428 545912
rect 206284 543720 206336 543726
rect 206284 543662 206336 543668
rect 206388 539963 206416 545906
rect 206480 543318 206508 547846
rect 207112 543720 207164 543726
rect 207112 543662 207164 543668
rect 206468 543312 206520 543318
rect 206468 543254 206520 543260
rect 207124 539963 207152 543662
rect 207860 539963 207888 557506
rect 208412 543930 208440 622610
rect 208492 616888 208544 616894
rect 208492 616830 208544 616836
rect 208504 557534 208532 616830
rect 209044 562352 209096 562358
rect 209044 562294 209096 562300
rect 208504 557506 208624 557534
rect 208400 543924 208452 543930
rect 208400 543866 208452 543872
rect 208596 539963 208624 557506
rect 209056 543726 209084 562294
rect 209792 543946 209820 625330
rect 210424 623960 210476 623966
rect 210424 623902 210476 623908
rect 210148 548548 210200 548554
rect 210148 548490 210200 548496
rect 209228 543924 209280 543930
rect 209792 543918 210004 543946
rect 209228 543866 209280 543872
rect 209044 543720 209096 543726
rect 209044 543662 209096 543668
rect 209240 539963 209268 543866
rect 209976 539963 210004 543918
rect 210160 543266 210188 548490
rect 210436 543386 210464 623902
rect 211804 622532 211856 622538
rect 211804 622474 211856 622480
rect 210516 589348 210568 589354
rect 210516 589290 210568 589296
rect 210528 551614 210556 589290
rect 211160 586900 211212 586906
rect 211160 586842 211212 586848
rect 210608 571396 210660 571402
rect 210608 571338 210660 571344
rect 210516 551608 210568 551614
rect 210516 551550 210568 551556
rect 210620 545766 210648 571338
rect 211068 547392 211120 547398
rect 211068 547334 211120 547340
rect 210608 545760 210660 545766
rect 210608 545702 210660 545708
rect 210424 543380 210476 543386
rect 210424 543322 210476 543328
rect 210160 543238 210740 543266
rect 210712 539963 210740 543238
rect 211080 543114 211108 547334
rect 211172 543946 211200 586842
rect 211620 551472 211672 551478
rect 211620 551414 211672 551420
rect 211172 543918 211476 543946
rect 211068 543108 211120 543114
rect 211068 543050 211120 543056
rect 211448 539963 211476 543918
rect 211632 543538 211660 551414
rect 211816 543658 211844 622474
rect 212552 543930 212580 625602
rect 213184 619676 213236 619682
rect 213184 619618 213236 619624
rect 212632 558476 212684 558482
rect 212632 558418 212684 558424
rect 212644 557534 212672 558418
rect 212644 557506 212856 557534
rect 212540 543924 212592 543930
rect 212540 543866 212592 543872
rect 211804 543652 211856 543658
rect 211804 543594 211856 543600
rect 211632 543510 212212 543538
rect 212184 539963 212212 543510
rect 212828 539963 212856 557506
rect 213196 550050 213224 619618
rect 213184 550044 213236 550050
rect 213184 549986 213236 549992
rect 213932 543930 213960 625738
rect 214012 625320 214064 625326
rect 214012 625262 214064 625268
rect 214024 557534 214052 625262
rect 215300 624096 215352 624102
rect 215300 624038 215352 624044
rect 214564 622804 214616 622810
rect 214564 622746 214616 622752
rect 214024 557506 214328 557534
rect 213552 543924 213604 543930
rect 213552 543866 213604 543872
rect 213920 543924 213972 543930
rect 213920 543866 213972 543872
rect 213564 539963 213592 543866
rect 214300 539963 214328 557506
rect 214576 543182 214604 622746
rect 215312 563054 215340 624038
rect 217324 622396 217376 622402
rect 217324 622338 217376 622344
rect 216678 620664 216734 620673
rect 216678 620599 216734 620608
rect 216692 619682 216720 620599
rect 216680 619676 216732 619682
rect 216680 619618 216732 619624
rect 216678 617808 216734 617817
rect 216678 617743 216734 617752
rect 216692 616894 216720 617743
rect 216680 616888 216732 616894
rect 216680 616830 216732 616836
rect 215942 611688 215998 611697
rect 215942 611623 215998 611632
rect 215312 563026 215800 563054
rect 215024 543924 215076 543930
rect 215024 543866 215076 543872
rect 214564 543176 214616 543182
rect 214564 543118 214616 543124
rect 215036 539963 215064 543866
rect 215772 539963 215800 563026
rect 215956 548758 215984 611623
rect 216678 608288 216734 608297
rect 216678 608223 216734 608232
rect 216692 607238 216720 608223
rect 216680 607232 216732 607238
rect 216680 607174 216732 607180
rect 217230 602168 217286 602177
rect 217230 602103 217286 602112
rect 216678 593464 216734 593473
rect 216678 593399 216680 593408
rect 216732 593399 216734 593408
rect 216680 593370 216732 593376
rect 216678 589928 216734 589937
rect 216678 589863 216734 589872
rect 216692 589354 216720 589863
rect 216680 589348 216732 589354
rect 216680 589290 216732 589296
rect 216678 587208 216734 587217
rect 216678 587143 216734 587152
rect 216692 586906 216720 587143
rect 216680 586900 216732 586906
rect 216680 586842 216732 586848
rect 216034 577688 216090 577697
rect 216034 577623 216090 577632
rect 215944 548752 215996 548758
rect 215944 548694 215996 548700
rect 216048 546038 216076 577623
rect 216678 574968 216734 574977
rect 216678 574903 216734 574912
rect 216692 574122 216720 574903
rect 216680 574116 216732 574122
rect 216680 574058 216732 574064
rect 216678 571568 216734 571577
rect 216678 571503 216734 571512
rect 216692 571402 216720 571503
rect 216680 571396 216732 571402
rect 216680 571338 216732 571344
rect 217138 562728 217194 562737
rect 217138 562663 217194 562672
rect 216128 559836 216180 559842
rect 216128 559778 216180 559784
rect 216036 546032 216088 546038
rect 216036 545974 216088 545980
rect 216140 543250 216168 559778
rect 216128 543244 216180 543250
rect 216128 543186 216180 543192
rect 216404 543108 216456 543114
rect 216404 543050 216456 543056
rect 216416 539963 216444 543050
rect 217152 539963 217180 562663
rect 217244 543726 217272 602103
rect 217336 551682 217364 622338
rect 217690 614408 217746 614417
rect 217690 614343 217746 614352
rect 217414 583808 217470 583817
rect 217414 583743 217470 583752
rect 217428 562358 217456 583743
rect 217704 581738 217732 614343
rect 217796 599593 217824 629886
rect 217876 625592 217928 625598
rect 217876 625534 217928 625540
rect 217782 599584 217838 599593
rect 217782 599519 217838 599528
rect 217692 581732 217744 581738
rect 217692 581674 217744 581680
rect 217690 581088 217746 581097
rect 217690 581023 217746 581032
rect 217598 565448 217654 565457
rect 217598 565383 217654 565392
rect 217416 562352 217468 562358
rect 217416 562294 217468 562300
rect 217324 551676 217376 551682
rect 217324 551618 217376 551624
rect 217232 543720 217284 543726
rect 217232 543662 217284 543668
rect 217612 543658 217640 565383
rect 217704 560318 217732 581023
rect 217692 560312 217744 560318
rect 217692 560254 217744 560260
rect 217888 559366 217916 625534
rect 217968 622872 218020 622878
rect 217968 622814 218020 622820
rect 217876 559360 217928 559366
rect 217876 559302 217928 559308
rect 217876 545896 217928 545902
rect 217876 545838 217928 545844
rect 217600 543652 217652 543658
rect 217600 543594 217652 543600
rect 217888 539963 217916 545838
rect 217980 543250 218008 622814
rect 218716 622470 218744 630634
rect 280712 630012 280764 630018
rect 280712 629954 280764 629960
rect 225420 625796 225472 625802
rect 225420 625738 225472 625744
rect 218888 625524 218940 625530
rect 218888 625466 218940 625472
rect 218796 625456 218848 625462
rect 218796 625398 218848 625404
rect 218704 622464 218756 622470
rect 218704 622406 218756 622412
rect 218716 596193 218744 622406
rect 218702 596184 218758 596193
rect 218702 596119 218758 596128
rect 218704 581732 218756 581738
rect 218704 581674 218756 581680
rect 218612 543720 218664 543726
rect 218612 543662 218664 543668
rect 217968 543244 218020 543250
rect 217968 543186 218020 543192
rect 218624 539963 218652 543662
rect 218716 543046 218744 581674
rect 218808 555762 218836 625398
rect 218900 559978 218928 625466
rect 219348 625252 219400 625258
rect 219348 625194 219400 625200
rect 219254 605568 219310 605577
rect 219254 605503 219310 605512
rect 219162 568848 219218 568857
rect 219162 568783 219218 568792
rect 218888 559972 218940 559978
rect 218888 559914 218940 559920
rect 218796 555756 218848 555762
rect 218796 555698 218848 555704
rect 219176 544542 219204 568783
rect 219268 557530 219296 605503
rect 219360 559094 219388 625194
rect 219624 624028 219676 624034
rect 219624 623970 219676 623976
rect 219636 615494 219664 623970
rect 225432 623098 225460 625738
rect 231308 625728 231360 625734
rect 231308 625670 231360 625676
rect 231320 623098 231348 625670
rect 271880 625660 271932 625666
rect 271880 625602 271932 625608
rect 242900 625592 242952 625598
rect 242900 625534 242952 625540
rect 234620 624096 234672 624102
rect 234620 624038 234672 624044
rect 234632 623098 234660 624038
rect 237564 623960 237616 623966
rect 237564 623902 237616 623908
rect 225432 623070 225814 623098
rect 231320 623070 231610 623098
rect 234632 623070 234830 623098
rect 237576 622962 237604 623902
rect 242912 623098 242940 625534
rect 251916 625524 251968 625530
rect 251916 625466 251968 625472
rect 246028 624028 246080 624034
rect 246028 623970 246080 623976
rect 246040 623098 246068 623970
rect 251928 623098 251956 625466
rect 263600 625456 263652 625462
rect 263600 625398 263652 625404
rect 260196 625388 260248 625394
rect 260196 625330 260248 625336
rect 254492 623892 254544 623898
rect 254492 623834 254544 623840
rect 254504 623098 254532 623834
rect 260208 623098 260236 625330
rect 263612 623098 263640 625398
rect 269212 625320 269264 625326
rect 269212 625262 269264 625268
rect 269224 623098 269252 625262
rect 271892 623098 271920 625602
rect 275100 625252 275152 625258
rect 275100 625194 275152 625200
rect 275112 623098 275140 625194
rect 277676 623824 277728 623830
rect 277676 623766 277728 623772
rect 277688 623098 277716 623766
rect 242912 623070 243202 623098
rect 246040 623070 246422 623098
rect 251928 623070 252218 623098
rect 254504 623070 254794 623098
rect 260208 623070 260590 623098
rect 263612 623070 263810 623098
rect 269224 623070 269606 623098
rect 271892 623070 272182 623098
rect 275112 623070 275402 623098
rect 277688 623070 277978 623098
rect 237406 622934 237604 622962
rect 228732 622872 228784 622878
rect 228784 622820 229034 622826
rect 228732 622814 229034 622820
rect 228744 622798 229034 622814
rect 257632 622810 258014 622826
rect 257620 622804 258014 622810
rect 257672 622798 258014 622804
rect 257620 622746 257672 622752
rect 222844 622736 222896 622742
rect 222896 622684 223238 622690
rect 222844 622678 223238 622684
rect 222856 622662 223238 622678
rect 240336 622674 240626 622690
rect 240324 622668 240626 622674
rect 240376 622662 240626 622668
rect 240324 622610 240376 622616
rect 248696 622600 248748 622606
rect 248748 622548 248998 622554
rect 248696 622542 248998 622548
rect 248708 622526 248998 622542
rect 266280 622538 266386 622554
rect 280724 622538 280752 629954
rect 266268 622532 266386 622538
rect 266320 622526 266386 622532
rect 280712 622532 280764 622538
rect 266268 622474 266320 622480
rect 280712 622474 280764 622480
rect 219728 622402 220018 622418
rect 219716 622396 220018 622402
rect 219768 622390 220018 622396
rect 280554 622390 280844 622418
rect 219716 622338 219768 622344
rect 280712 622328 280764 622334
rect 280712 622270 280764 622276
rect 219636 615466 219756 615494
rect 219728 563054 219756 615466
rect 219728 563026 219848 563054
rect 219348 559088 219400 559094
rect 219348 559030 219400 559036
rect 219256 557524 219308 557530
rect 219256 557466 219308 557472
rect 219532 556776 219584 556782
rect 219532 556718 219584 556724
rect 219164 544536 219216 544542
rect 219164 544478 219216 544484
rect 219544 543726 219572 556718
rect 219820 553394 219848 563026
rect 220176 560312 220228 560318
rect 220176 560254 220228 560260
rect 219912 560102 220018 560130
rect 219912 556782 219940 560102
rect 219900 556776 219952 556782
rect 219900 556718 219952 556724
rect 220188 553394 220216 560254
rect 222594 560102 222976 560130
rect 222200 559360 222252 559366
rect 222200 559302 222252 559308
rect 219728 553366 219848 553394
rect 220096 553366 220216 553394
rect 219728 543946 219756 553366
rect 219728 543918 220032 543946
rect 219532 543720 219584 543726
rect 219532 543662 219584 543668
rect 219256 543652 219308 543658
rect 219256 543594 219308 543600
rect 218704 543040 218756 543046
rect 218704 542982 218756 542988
rect 219268 539963 219296 543594
rect 220004 539963 220032 543918
rect 220096 543182 220124 553366
rect 220728 544468 220780 544474
rect 220728 544410 220780 544416
rect 220084 543176 220136 543182
rect 220084 543118 220136 543124
rect 220740 539963 220768 544410
rect 222212 543930 222240 559302
rect 222292 558544 222344 558550
rect 222292 558486 222344 558492
rect 222200 543924 222252 543930
rect 222200 543866 222252 543872
rect 221464 543720 221516 543726
rect 221464 543662 221516 543668
rect 221476 539963 221504 543662
rect 222304 540138 222332 558486
rect 222948 557598 222976 560102
rect 225064 560102 225170 560130
rect 228008 560102 228390 560130
rect 230492 560102 230966 560130
rect 233896 560102 234186 560130
rect 236012 560102 236762 560130
rect 238772 560102 239982 560130
rect 241532 560102 242558 560130
rect 245672 560102 245778 560130
rect 247144 560102 248354 560130
rect 251192 560102 251574 560130
rect 253952 560102 254150 560130
rect 257080 560102 257370 560130
rect 259656 560102 259946 560130
rect 262784 560102 263166 560130
rect 265360 560102 265742 560130
rect 268672 560102 268962 560130
rect 271248 560102 271538 560130
rect 274652 560102 274758 560130
rect 276952 560102 277334 560130
rect 280264 560102 280554 560130
rect 223580 559088 223632 559094
rect 223580 559030 223632 559036
rect 222936 557592 222988 557598
rect 222936 557534 222988 557540
rect 222844 543924 222896 543930
rect 222844 543866 222896 543872
rect 222228 540110 222332 540138
rect 222228 539920 222256 540110
rect 222856 539963 222884 543866
rect 223592 539963 223620 559030
rect 224408 557592 224460 557598
rect 224408 557534 224460 557540
rect 223672 557524 223724 557530
rect 223672 557466 223724 557472
rect 223684 543946 223712 557466
rect 223684 543918 224356 543946
rect 224328 539963 224356 543918
rect 224420 543726 224448 557534
rect 225064 550186 225092 560102
rect 228008 558822 228036 560102
rect 225144 558816 225196 558822
rect 225144 558758 225196 558764
rect 227996 558816 228048 558822
rect 227996 558758 228048 558764
rect 225052 550180 225104 550186
rect 225052 550122 225104 550128
rect 224408 543720 224460 543726
rect 224408 543662 224460 543668
rect 225156 540138 225184 558758
rect 227720 558340 227772 558346
rect 227720 558282 227772 558288
rect 226432 552968 226484 552974
rect 226432 552910 226484 552916
rect 225788 543720 225840 543726
rect 225788 543662 225840 543668
rect 225080 540110 225184 540138
rect 225080 539920 225108 540110
rect 225800 539963 225828 543662
rect 226444 539963 226472 552910
rect 227168 544536 227220 544542
rect 227168 544478 227220 544484
rect 227180 539963 227208 544478
rect 227732 543946 227760 558282
rect 230492 557534 230520 560102
rect 231952 558612 232004 558618
rect 231952 558554 232004 558560
rect 231964 557534 231992 558554
rect 233896 558414 233924 560102
rect 233884 558408 233936 558414
rect 233884 558350 233936 558356
rect 230492 557506 230796 557534
rect 231964 557506 232268 557534
rect 229284 557048 229336 557054
rect 229284 556990 229336 556996
rect 228640 550180 228692 550186
rect 228640 550122 228692 550128
rect 227732 543918 227944 543946
rect 227916 539963 227944 543918
rect 228652 539963 228680 550122
rect 229296 539963 229324 556990
rect 230020 543244 230072 543250
rect 230020 543186 230072 543192
rect 230032 539963 230060 543186
rect 230768 539963 230796 557506
rect 231492 543244 231544 543250
rect 231492 543186 231544 543192
rect 231504 539963 231532 543186
rect 232240 539963 232268 557506
rect 236012 547398 236040 560102
rect 236000 547392 236052 547398
rect 236000 547334 236052 547340
rect 235080 547324 235132 547330
rect 235080 547266 235132 547272
rect 234344 545760 234396 545766
rect 234344 545702 234396 545708
rect 232872 543176 232924 543182
rect 232872 543118 232924 543124
rect 232884 539963 232912 543118
rect 233608 543040 233660 543046
rect 233608 542982 233660 542988
rect 233620 539963 233648 542982
rect 234356 539963 234384 545702
rect 235092 539963 235120 547266
rect 237932 543788 237984 543794
rect 237932 543730 237984 543736
rect 237196 543516 237248 543522
rect 237196 543458 237248 543464
rect 235816 541884 235868 541890
rect 235816 541826 235868 541832
rect 235828 539963 235856 541826
rect 236460 541204 236512 541210
rect 236460 541146 236512 541152
rect 236472 539963 236500 541146
rect 237208 539963 237236 543458
rect 237944 539963 237972 543730
rect 238772 543250 238800 560102
rect 240784 555688 240836 555694
rect 240784 555630 240836 555636
rect 238760 543244 238812 543250
rect 238760 543186 238812 543192
rect 238668 543176 238720 543182
rect 238668 543118 238720 543124
rect 238680 539963 238708 543118
rect 240796 543114 240824 555630
rect 241532 545970 241560 560102
rect 245672 558346 245700 560102
rect 247040 559768 247092 559774
rect 247040 559710 247092 559716
rect 245660 558340 245712 558346
rect 245660 558282 245712 558288
rect 245108 555620 245160 555626
rect 245108 555562 245160 555568
rect 242900 550044 242952 550050
rect 242900 549986 242952 549992
rect 241520 545964 241572 545970
rect 241520 545906 241572 545912
rect 242256 543312 242308 543318
rect 242256 543254 242308 543260
rect 240784 543108 240836 543114
rect 240784 543050 240836 543056
rect 239402 543008 239458 543017
rect 239402 542943 239458 542952
rect 240784 542972 240836 542978
rect 239416 539963 239444 542943
rect 240784 542914 240836 542920
rect 240048 541340 240100 541346
rect 240048 541282 240100 541288
rect 240060 539963 240088 541282
rect 240796 539963 240824 542914
rect 241518 542600 241574 542609
rect 241518 542535 241574 542544
rect 241532 539963 241560 542535
rect 242268 539963 242296 543254
rect 242912 539963 242940 549986
rect 243636 541544 243688 541550
rect 243636 541486 243688 541492
rect 243648 539963 243676 541486
rect 244372 541476 244424 541482
rect 244372 541418 244424 541424
rect 244384 539963 244412 541418
rect 245120 539963 245148 555562
rect 246488 554260 246540 554266
rect 246488 554202 246540 554208
rect 245844 543108 245896 543114
rect 245844 543050 245896 543056
rect 245856 539963 245884 543050
rect 246500 539963 246528 554202
rect 247052 543946 247080 559710
rect 247144 544474 247172 560102
rect 251192 558482 251220 560102
rect 253952 558550 253980 560102
rect 253940 558544 253992 558550
rect 253940 558486 253992 558492
rect 251180 558476 251232 558482
rect 251180 558418 251232 558424
rect 249800 558340 249852 558346
rect 249800 558282 249852 558288
rect 247132 544468 247184 544474
rect 247132 544410 247184 544416
rect 249812 543946 249840 558282
rect 257080 558278 257108 560102
rect 258080 559904 258132 559910
rect 258080 559846 258132 559852
rect 257068 558272 257120 558278
rect 257068 558214 257120 558220
rect 258092 557534 258120 559846
rect 259656 558618 259684 560102
rect 260840 559972 260892 559978
rect 260840 559914 260892 559920
rect 260104 558816 260156 558822
rect 260104 558758 260156 558764
rect 259644 558612 259696 558618
rect 259644 558554 259696 558560
rect 258092 557506 258764 557534
rect 256700 552900 256752 552906
rect 256700 552842 256752 552848
rect 250812 552832 250864 552838
rect 250812 552774 250864 552780
rect 247052 543918 248000 543946
rect 249812 543918 250116 543946
rect 247224 541068 247276 541074
rect 247224 541010 247276 541016
rect 247236 539963 247264 541010
rect 247972 539963 248000 543918
rect 248694 542736 248750 542745
rect 248694 542671 248750 542680
rect 248708 539963 248736 542671
rect 249432 541136 249484 541142
rect 249432 541078 249484 541084
rect 249444 539963 249472 541078
rect 250088 539963 250116 543918
rect 250824 539963 250852 552774
rect 253664 551540 253716 551546
rect 253664 551482 253716 551488
rect 251548 550112 251600 550118
rect 251548 550054 251600 550060
rect 251560 539963 251588 550054
rect 252284 543856 252336 543862
rect 252284 543798 252336 543804
rect 252296 539963 252324 543798
rect 252928 543380 252980 543386
rect 252928 543322 252980 543328
rect 252940 539963 252968 543322
rect 253676 539963 253704 551482
rect 256712 543930 256740 552842
rect 256700 543924 256752 543930
rect 256700 543866 256752 543872
rect 257988 543924 258040 543930
rect 257988 543866 258040 543872
rect 255134 543280 255190 543289
rect 255134 543215 255190 543224
rect 254400 541272 254452 541278
rect 254400 541214 254452 541220
rect 254412 539963 254440 541214
rect 255148 539963 255176 543215
rect 256514 543144 256570 543153
rect 256514 543079 256570 543088
rect 255872 541408 255924 541414
rect 255872 541350 255924 541356
rect 255884 539963 255912 541350
rect 256528 539963 256556 543079
rect 257252 542700 257304 542706
rect 257252 542642 257304 542648
rect 257264 539963 257292 542642
rect 258000 539963 258028 543866
rect 258736 539963 258764 557506
rect 260012 551608 260064 551614
rect 260012 551550 260064 551556
rect 259552 547392 259604 547398
rect 259552 547334 259604 547340
rect 259564 540138 259592 547334
rect 260024 545714 260052 551550
rect 260116 545902 260144 558758
rect 260852 557534 260880 559914
rect 262784 558822 262812 560102
rect 262772 558816 262824 558822
rect 262772 558758 262824 558764
rect 265360 557938 265388 560102
rect 264244 557932 264296 557938
rect 264244 557874 264296 557880
rect 265348 557932 265400 557938
rect 265348 557874 265400 557880
rect 262864 557660 262916 557666
rect 262864 557602 262916 557608
rect 260852 557506 261616 557534
rect 260104 545896 260156 545902
rect 260104 545838 260156 545844
rect 260024 545686 260144 545714
rect 259488 540110 259592 540138
rect 259488 539920 259516 540110
rect 260116 539963 260144 545686
rect 260840 541612 260892 541618
rect 260840 541554 260892 541560
rect 260852 539963 260880 541554
rect 261588 539963 261616 557506
rect 262876 549982 262904 557602
rect 263692 554192 263744 554198
rect 263692 554134 263744 554140
rect 262864 549976 262916 549982
rect 262864 549918 262916 549924
rect 263048 540320 263100 540326
rect 263048 540262 263100 540268
rect 262312 540184 262364 540190
rect 262312 540126 262364 540132
rect 262324 539963 262352 540126
rect 263060 539963 263088 540262
rect 263704 539963 263732 554134
rect 264256 548622 264284 557874
rect 268672 557666 268700 560102
rect 268660 557660 268712 557666
rect 268660 557602 268712 557608
rect 267740 557592 267792 557598
rect 267740 557534 267792 557540
rect 267752 557506 268056 557534
rect 266544 555756 266596 555762
rect 266544 555698 266596 555704
rect 264244 548616 264296 548622
rect 264244 548558 264296 548564
rect 265900 541680 265952 541686
rect 265900 541622 265952 541628
rect 264426 541104 264482 541113
rect 264426 541039 264482 541048
rect 264440 539963 264468 541039
rect 265164 540388 265216 540394
rect 265164 540330 265216 540336
rect 265176 539963 265204 540330
rect 265912 539963 265940 541622
rect 266556 539963 266584 555698
rect 267280 545964 267332 545970
rect 267280 545906 267332 545912
rect 267292 539963 267320 545906
rect 268028 539963 268056 557506
rect 269488 557116 269540 557122
rect 269488 557058 269540 557064
rect 268752 541816 268804 541822
rect 268752 541758 268804 541764
rect 268764 539963 268792 541758
rect 269500 539963 269528 557058
rect 271248 552702 271276 560102
rect 273260 558272 273312 558278
rect 273260 558214 273312 558220
rect 271236 552696 271288 552702
rect 271236 552638 271288 552644
rect 271604 549976 271656 549982
rect 271604 549918 271656 549924
rect 270132 544536 270184 544542
rect 270132 544478 270184 544484
rect 270144 539963 270172 544478
rect 270868 542904 270920 542910
rect 270868 542846 270920 542852
rect 270880 539963 270908 542846
rect 271616 539963 271644 549918
rect 273272 547126 273300 558214
rect 274652 547262 274680 560102
rect 276952 558210 276980 560102
rect 280264 558822 280292 560102
rect 278044 558816 278096 558822
rect 278044 558758 278096 558764
rect 280252 558816 280304 558822
rect 280252 558758 280304 558764
rect 276940 558204 276992 558210
rect 276940 558146 276992 558152
rect 274640 547256 274692 547262
rect 274640 547198 274692 547204
rect 273260 547120 273312 547126
rect 273260 547062 273312 547068
rect 274456 547120 274508 547126
rect 274456 547062 274508 547068
rect 273720 542836 273772 542842
rect 273720 542778 273772 542784
rect 272340 541000 272392 541006
rect 272340 540942 272392 540948
rect 272352 539963 272380 540942
rect 273076 540252 273128 540258
rect 273076 540194 273128 540200
rect 273088 539963 273116 540194
rect 273732 539963 273760 542778
rect 274468 539963 274496 547062
rect 275192 545896 275244 545902
rect 275192 545838 275244 545844
rect 275204 539963 275232 545838
rect 278056 545834 278084 558758
rect 280724 547874 280752 622270
rect 280816 552974 280844 622390
rect 280894 616992 280950 617001
rect 280894 616927 280950 616936
rect 280804 552968 280856 552974
rect 280804 552910 280856 552916
rect 280908 550186 280936 616927
rect 280986 594960 281042 594969
rect 280986 594895 281042 594904
rect 281000 551478 281028 594895
rect 280988 551472 281040 551478
rect 280988 551414 281040 551420
rect 280896 550180 280948 550186
rect 280896 550122 280948 550128
rect 280724 547846 280936 547874
rect 278044 545828 278096 545834
rect 278044 545770 278096 545776
rect 279516 544468 279568 544474
rect 279516 544410 279568 544416
rect 277308 543448 277360 543454
rect 277308 543390 277360 543396
rect 275928 542972 275980 542978
rect 275928 542914 275980 542920
rect 275940 539963 275968 542914
rect 276572 542768 276624 542774
rect 276572 542710 276624 542716
rect 276584 539963 276612 542710
rect 277320 539963 277348 543390
rect 278044 543244 278096 543250
rect 278044 543186 278096 543192
rect 278056 539963 278084 543186
rect 278780 540456 278832 540462
rect 278780 540398 278832 540404
rect 278792 539963 278820 540398
rect 279528 539963 279556 544410
rect 280160 542496 280212 542502
rect 280160 542438 280212 542444
rect 280172 539963 280200 542438
rect 280908 539963 280936 547846
rect 281092 543114 281120 632159
rect 284944 631372 284996 631378
rect 284944 631314 284996 631320
rect 281906 619984 281962 619993
rect 281906 619919 281962 619928
rect 281630 611144 281686 611153
rect 281630 611079 281686 611088
rect 281170 592784 281226 592793
rect 281170 592719 281226 592728
rect 281184 548554 281212 592719
rect 281538 568304 281594 568313
rect 281538 568239 281594 568248
rect 281262 564904 281318 564913
rect 281262 564839 281318 564848
rect 281276 557054 281304 564839
rect 281552 559706 281580 568239
rect 281540 559700 281592 559706
rect 281540 559642 281592 559648
rect 281264 557048 281316 557054
rect 281264 556990 281316 556996
rect 281540 551676 281592 551682
rect 281540 551618 281592 551624
rect 281172 548548 281224 548554
rect 281172 548490 281224 548496
rect 281552 543946 281580 551618
rect 281644 544406 281672 611079
rect 281722 586664 281778 586673
rect 281722 586599 281778 586608
rect 281736 555558 281764 586599
rect 281814 580544 281870 580553
rect 281814 580479 281870 580488
rect 281724 555552 281776 555558
rect 281724 555494 281776 555500
rect 281828 551410 281856 580479
rect 281920 556918 281948 619919
rect 282918 613864 282974 613873
rect 282918 613799 282974 613808
rect 281998 562184 282054 562193
rect 281998 562119 282054 562128
rect 281908 556912 281960 556918
rect 281908 556854 281960 556860
rect 282012 554062 282040 562119
rect 282932 559842 282960 613799
rect 283010 607744 283066 607753
rect 283010 607679 283066 607688
rect 282920 559836 282972 559842
rect 282920 559778 282972 559784
rect 282000 554056 282052 554062
rect 282000 553998 282052 554004
rect 282920 551472 282972 551478
rect 282920 551414 282972 551420
rect 281816 551404 281868 551410
rect 281816 551346 281868 551352
rect 281632 544400 281684 544406
rect 281632 544342 281684 544348
rect 282932 543946 282960 551414
rect 283024 547194 283052 607679
rect 283194 605024 283250 605033
rect 283194 604959 283250 604968
rect 283102 601624 283158 601633
rect 283102 601559 283158 601568
rect 283116 549914 283144 601559
rect 283208 559638 283236 604959
rect 283286 598904 283342 598913
rect 283286 598839 283342 598848
rect 283196 559632 283248 559638
rect 283196 559574 283248 559580
rect 283300 552770 283328 598839
rect 283654 589384 283710 589393
rect 283654 589319 283656 589328
rect 283708 589319 283710 589328
rect 283656 589290 283708 589296
rect 283378 583264 283434 583273
rect 283378 583199 283434 583208
rect 283392 554130 283420 583199
rect 283562 577144 283618 577153
rect 283562 577079 283618 577088
rect 283470 574424 283526 574433
rect 283470 574359 283526 574368
rect 283484 555694 283512 574359
rect 283472 555688 283524 555694
rect 283472 555630 283524 555636
rect 283380 554124 283432 554130
rect 283380 554066 283432 554072
rect 283288 552764 283340 552770
rect 283288 552706 283340 552712
rect 283576 551342 283604 577079
rect 283654 571024 283710 571033
rect 283654 570959 283710 570968
rect 283668 556986 283696 570959
rect 283656 556980 283708 556986
rect 283656 556922 283708 556928
rect 283564 551336 283616 551342
rect 283564 551278 283616 551284
rect 283104 549908 283156 549914
rect 283104 549850 283156 549856
rect 283012 547188 283064 547194
rect 283012 547130 283064 547136
rect 281552 543918 282408 543946
rect 282932 543918 283788 543946
rect 281080 543108 281132 543114
rect 281080 543050 281132 543056
rect 281632 541748 281684 541754
rect 281632 541690 281684 541696
rect 281644 539963 281672 541690
rect 282380 539963 282408 543918
rect 283104 542632 283156 542638
rect 283104 542574 283156 542580
rect 283116 539963 283144 542574
rect 283760 539963 283788 543918
rect 284300 543516 284352 543522
rect 284300 543458 284352 543464
rect 284312 541657 284340 543458
rect 284956 543046 284984 631314
rect 285036 631304 285088 631310
rect 285036 631246 285088 631252
rect 285048 543153 285076 631246
rect 287060 630896 287112 630902
rect 287060 630838 287112 630844
rect 286324 615528 286376 615534
rect 286324 615470 286376 615476
rect 286336 559570 286364 615470
rect 286324 559564 286376 559570
rect 286324 559506 286376 559512
rect 287072 557534 287100 630838
rect 287704 610020 287756 610026
rect 287704 609962 287756 609968
rect 287072 557506 287560 557534
rect 287532 544354 287560 557506
rect 287716 554266 287744 609962
rect 287796 596216 287848 596222
rect 287796 596158 287848 596164
rect 287704 554260 287756 554266
rect 287704 554202 287756 554208
rect 287808 544542 287836 596158
rect 288452 557534 288480 633422
rect 289084 625184 289136 625190
rect 289084 625126 289136 625132
rect 288452 557506 288848 557534
rect 287796 544536 287848 544542
rect 287796 544478 287848 544484
rect 287532 544326 288112 544354
rect 287428 544128 287480 544134
rect 287428 544070 287480 544076
rect 285220 543924 285272 543930
rect 285220 543866 285272 543872
rect 285034 543144 285090 543153
rect 285034 543079 285090 543088
rect 284944 543040 284996 543046
rect 284944 542982 284996 542988
rect 284484 542564 284536 542570
rect 284484 542506 284536 542512
rect 284298 541648 284354 541657
rect 284298 541583 284354 541592
rect 284496 539963 284524 542506
rect 285232 539963 285260 543866
rect 285954 542872 286010 542881
rect 285954 542807 286010 542816
rect 285968 539963 285996 542807
rect 286690 542464 286746 542473
rect 286690 542399 286746 542408
rect 286704 539963 286732 542399
rect 287440 540138 287468 544070
rect 287364 540110 287468 540138
rect 287364 539920 287392 540110
rect 288084 539963 288112 544326
rect 288820 539963 288848 557506
rect 289096 549982 289124 625126
rect 289176 571396 289228 571402
rect 289176 571338 289228 571344
rect 289188 551614 289216 571338
rect 289832 557534 289860 633558
rect 296720 633548 296772 633554
rect 296720 633490 296772 633496
rect 291200 631100 291252 631106
rect 291200 631042 291252 631048
rect 289832 557506 290228 557534
rect 289176 551608 289228 551614
rect 289176 551550 289228 551556
rect 289084 549976 289136 549982
rect 289084 549918 289136 549924
rect 289544 545148 289596 545154
rect 289544 545090 289596 545096
rect 289556 539963 289584 545090
rect 290200 539963 290228 557506
rect 290924 544196 290976 544202
rect 290924 544138 290976 544144
rect 290936 539963 290964 544138
rect 291212 543998 291240 631042
rect 293960 630964 294012 630970
rect 293960 630906 294012 630912
rect 293224 586560 293276 586566
rect 293224 586502 293276 586508
rect 293236 551682 293264 586502
rect 293224 551676 293276 551682
rect 293224 551618 293276 551624
rect 293972 543998 294000 630906
rect 294604 600364 294656 600370
rect 294604 600306 294656 600312
rect 294616 558346 294644 600306
rect 294604 558340 294656 558346
rect 294604 558282 294656 558288
rect 296732 557534 296760 633490
rect 296732 557506 297404 557534
rect 291200 543992 291252 543998
rect 291200 543934 291252 543940
rect 292396 543992 292448 543998
rect 292396 543934 292448 543940
rect 293960 543992 294012 543998
rect 293960 543934 294012 543940
rect 295248 543992 295300 543998
rect 295248 543934 295300 543940
rect 291658 541376 291714 541385
rect 291658 541311 291714 541320
rect 291672 539963 291700 541311
rect 292408 539963 292436 543934
rect 294510 541240 294566 541249
rect 294510 541175 294566 541184
rect 293776 540592 293828 540598
rect 293776 540534 293828 540540
rect 293132 540524 293184 540530
rect 293132 540466 293184 540472
rect 293144 539963 293172 540466
rect 293788 539963 293816 540534
rect 294524 539963 294552 541175
rect 295260 539963 295288 543934
rect 296720 542428 296772 542434
rect 296720 542370 296772 542376
rect 295984 540796 296036 540802
rect 295984 540738 296036 540744
rect 295996 539963 296024 540738
rect 296732 539963 296760 542370
rect 297376 539963 297404 557506
rect 298112 541822 298140 633626
rect 300124 632936 300176 632942
rect 300124 632878 300176 632884
rect 298192 631236 298244 631242
rect 298192 631178 298244 631184
rect 298100 541816 298152 541822
rect 298100 541758 298152 541764
rect 298204 540138 298232 631178
rect 300136 545970 300164 632878
rect 304264 605872 304316 605878
rect 304264 605814 304316 605820
rect 302240 589960 302292 589966
rect 302240 589902 302292 589908
rect 302252 589354 302280 589902
rect 302240 589348 302292 589354
rect 302240 589290 302292 589296
rect 300216 576904 300268 576910
rect 300216 576846 300268 576852
rect 300228 557122 300256 576846
rect 302252 560250 302280 589290
rect 302240 560244 302292 560250
rect 302240 560186 302292 560192
rect 300216 557116 300268 557122
rect 300216 557058 300268 557064
rect 300124 545964 300176 545970
rect 300124 545906 300176 545912
rect 301780 543380 301832 543386
rect 301780 543322 301832 543328
rect 301596 543312 301648 543318
rect 301596 543254 301648 543260
rect 299572 543040 299624 543046
rect 299572 542982 299624 542988
rect 298836 541816 298888 541822
rect 298836 541758 298888 541764
rect 298128 540110 298232 540138
rect 298128 539920 298156 540110
rect 298848 539963 298876 541758
rect 299584 539963 299612 542982
rect 300584 542904 300636 542910
rect 300584 542846 300636 542852
rect 300214 542736 300270 542745
rect 300214 542671 300270 542680
rect 300400 542700 300452 542706
rect 300124 542632 300176 542638
rect 300124 542574 300176 542580
rect 300136 517206 300164 542574
rect 300228 518809 300256 542671
rect 300400 542642 300452 542648
rect 300308 541680 300360 541686
rect 300308 541622 300360 541628
rect 300214 518800 300270 518809
rect 300214 518735 300270 518744
rect 300320 518430 300348 541622
rect 300412 520062 300440 542642
rect 300492 541000 300544 541006
rect 300492 540942 300544 540948
rect 300400 520056 300452 520062
rect 300400 519998 300452 520004
rect 300308 518424 300360 518430
rect 300308 518366 300360 518372
rect 300504 518022 300532 540942
rect 300596 520130 300624 542846
rect 301502 542464 301558 542473
rect 301502 542399 301558 542408
rect 300676 541544 300728 541550
rect 300676 541486 300728 541492
rect 300688 529922 300716 541486
rect 300860 540456 300912 540462
rect 300860 540398 300912 540404
rect 300872 539578 300900 540398
rect 300860 539572 300912 539578
rect 300860 539514 300912 539520
rect 300676 529916 300728 529922
rect 300676 529858 300728 529864
rect 300584 520124 300636 520130
rect 300584 520066 300636 520072
rect 300492 518016 300544 518022
rect 300492 517958 300544 517964
rect 300124 517200 300176 517206
rect 300124 517142 300176 517148
rect 301516 516118 301544 542399
rect 301608 517138 301636 543254
rect 301688 542564 301740 542570
rect 301688 542506 301740 542512
rect 301596 517132 301648 517138
rect 301596 517074 301648 517080
rect 301700 517070 301728 542506
rect 301792 518158 301820 543322
rect 301964 542972 302016 542978
rect 301964 542914 302016 542920
rect 301872 542496 301924 542502
rect 301872 542438 301924 542444
rect 301884 519994 301912 542438
rect 301872 519988 301924 519994
rect 301872 519930 301924 519936
rect 301976 519246 302004 542914
rect 302056 541884 302108 541890
rect 302056 541826 302108 541832
rect 301964 519240 302016 519246
rect 301964 519182 302016 519188
rect 302068 518498 302096 541826
rect 302056 518492 302108 518498
rect 302056 518434 302108 518440
rect 301780 518152 301832 518158
rect 301780 518094 301832 518100
rect 301688 517064 301740 517070
rect 301688 517006 301740 517012
rect 301504 516112 301556 516118
rect 301504 516054 301556 516060
rect 57702 509960 57758 509969
rect 42708 509924 42760 509930
rect 57702 509895 57704 509904
rect 42708 509866 42760 509872
rect 57756 509895 57758 509904
rect 57886 509960 57942 509969
rect 57886 509895 57942 509904
rect 57704 509866 57756 509872
rect 42432 470280 42484 470286
rect 42432 470222 42484 470228
rect 42340 470144 42392 470150
rect 42340 470086 42392 470092
rect 42156 469056 42208 469062
rect 42156 468998 42208 469004
rect 42168 373969 42196 468998
rect 42248 464364 42300 464370
rect 42248 464306 42300 464312
rect 42154 373960 42210 373969
rect 42154 373895 42210 373904
rect 42260 267646 42288 464306
rect 42248 267640 42300 267646
rect 42248 267582 42300 267588
rect 42352 267510 42380 470086
rect 42340 267504 42392 267510
rect 42340 267446 42392 267452
rect 42444 263566 42472 470222
rect 42524 468920 42576 468926
rect 42524 468862 42576 468868
rect 42432 263560 42484 263566
rect 42432 263502 42484 263508
rect 42064 202836 42116 202842
rect 42064 202778 42116 202784
rect 42536 164422 42564 468862
rect 42614 466304 42670 466313
rect 42614 466239 42670 466248
rect 42524 164416 42576 164422
rect 42524 164358 42576 164364
rect 41328 164280 41380 164286
rect 41328 164222 41380 164228
rect 42628 58818 42656 466239
rect 42720 382226 42748 509866
rect 302252 502489 302280 560186
rect 304276 551478 304304 605814
rect 304356 582412 304408 582418
rect 304356 582354 304408 582360
rect 304368 561134 304396 582354
rect 304356 561128 304408 561134
rect 304356 561070 304408 561076
rect 304264 551472 304316 551478
rect 304264 551414 304316 551420
rect 303068 543448 303120 543454
rect 303068 543390 303120 543396
rect 302884 542428 302936 542434
rect 302884 542370 302936 542376
rect 302330 532400 302386 532409
rect 302330 532335 302386 532344
rect 302344 532234 302372 532335
rect 302332 532228 302384 532234
rect 302332 532170 302384 532176
rect 302606 517440 302662 517449
rect 302606 517375 302662 517384
rect 302620 516186 302648 517375
rect 302896 517342 302924 542370
rect 302976 541476 303028 541482
rect 302976 541418 303028 541424
rect 302988 518090 303016 541418
rect 303080 519926 303108 543390
rect 304264 542836 304316 542842
rect 304264 542778 304316 542784
rect 303160 541340 303212 541346
rect 303160 541282 303212 541288
rect 303172 525774 303200 541282
rect 303160 525768 303212 525774
rect 303160 525710 303212 525716
rect 303068 519920 303120 519926
rect 303068 519862 303120 519868
rect 304276 519110 304304 542778
rect 304356 541204 304408 541210
rect 304356 541146 304408 541152
rect 304368 535430 304396 541146
rect 304356 535424 304408 535430
rect 304356 535366 304408 535372
rect 304356 532228 304408 532234
rect 304356 532170 304408 532176
rect 304264 519104 304316 519110
rect 304264 519046 304316 519052
rect 302976 518084 303028 518090
rect 302976 518026 303028 518032
rect 302884 517336 302936 517342
rect 302884 517278 302936 517284
rect 302608 516180 302660 516186
rect 302608 516122 302660 516128
rect 304368 515438 304396 532170
rect 305656 519178 305684 700334
rect 317052 639600 317104 639606
rect 317052 639542 317104 639548
rect 316868 634908 316920 634914
rect 316868 634850 316920 634856
rect 316684 633004 316736 633010
rect 316684 632946 316736 632952
rect 312544 632800 312596 632806
rect 312544 632742 312596 632748
rect 307024 632596 307076 632602
rect 307024 632538 307076 632544
rect 307036 555762 307064 632538
rect 309784 629332 309836 629338
rect 309784 629274 309836 629280
rect 307024 555756 307076 555762
rect 307024 555698 307076 555704
rect 309796 547398 309824 629274
rect 311164 619676 311216 619682
rect 311164 619618 311216 619624
rect 309784 547392 309836 547398
rect 309784 547334 309836 547340
rect 311176 544474 311204 619618
rect 312556 545902 312584 632742
rect 313924 632528 313976 632534
rect 313924 632470 313976 632476
rect 313936 550118 313964 632470
rect 314016 632324 314068 632330
rect 314016 632266 314068 632272
rect 313924 550112 313976 550118
rect 313924 550054 313976 550060
rect 314028 550050 314056 632266
rect 315304 632256 315356 632262
rect 315304 632198 315356 632204
rect 315316 554198 315344 632198
rect 315304 554192 315356 554198
rect 315304 554134 315356 554140
rect 316696 551546 316724 632946
rect 316776 632392 316828 632398
rect 316776 632334 316828 632340
rect 316788 552906 316816 632334
rect 316880 559910 316908 634850
rect 316960 634840 317012 634846
rect 316960 634782 317012 634788
rect 316972 559978 317000 634782
rect 317064 568313 317092 639542
rect 318800 634092 318852 634098
rect 318800 634034 318852 634040
rect 318248 632868 318300 632874
rect 318248 632810 318300 632816
rect 318156 632664 318208 632670
rect 318156 632606 318208 632612
rect 318064 631032 318116 631038
rect 318064 630974 318116 630980
rect 317786 629640 317842 629649
rect 317786 629575 317842 629584
rect 317800 629338 317828 629575
rect 317788 629332 317840 629338
rect 317788 629274 317840 629280
rect 317602 625288 317658 625297
rect 317602 625223 317658 625232
rect 317616 625190 317644 625223
rect 317604 625184 317656 625190
rect 317604 625126 317656 625132
rect 317970 620120 318026 620129
rect 317970 620055 318026 620064
rect 317984 619682 318012 620055
rect 317972 619676 318024 619682
rect 317972 619618 318024 619624
rect 317970 615632 318026 615641
rect 317970 615567 318026 615576
rect 317984 615534 318012 615567
rect 317972 615528 318024 615534
rect 317972 615470 318024 615476
rect 317878 610600 317934 610609
rect 317878 610535 317934 610544
rect 317892 610026 317920 610535
rect 317880 610020 317932 610026
rect 317880 609962 317932 609968
rect 317970 606112 318026 606121
rect 317970 606047 318026 606056
rect 317984 605878 318012 606047
rect 317972 605872 318024 605878
rect 317972 605814 318024 605820
rect 317602 601080 317658 601089
rect 317602 601015 317658 601024
rect 317616 600370 317644 601015
rect 317604 600364 317656 600370
rect 317604 600306 317656 600312
rect 317602 596456 317658 596465
rect 317602 596391 317658 596400
rect 317616 596222 317644 596391
rect 317604 596216 317656 596222
rect 317604 596158 317656 596164
rect 317420 586560 317472 586566
rect 317418 586528 317420 586537
rect 317472 586528 317474 586537
rect 317418 586463 317474 586472
rect 317970 582584 318026 582593
rect 317970 582519 318026 582528
rect 317984 582418 318012 582519
rect 317972 582412 318024 582418
rect 317972 582354 318024 582360
rect 317878 577280 317934 577289
rect 317878 577215 317934 577224
rect 317892 576910 317920 577215
rect 317880 576904 317932 576910
rect 317880 576846 317932 576852
rect 317970 571840 318026 571849
rect 317970 571775 318026 571784
rect 317984 571402 318012 571775
rect 317972 571396 318024 571402
rect 317972 571338 318024 571344
rect 317050 568304 317106 568313
rect 317050 568239 317106 568248
rect 316960 559972 317012 559978
rect 316960 559914 317012 559920
rect 316868 559904 316920 559910
rect 316868 559846 316920 559852
rect 317418 557696 317474 557705
rect 317418 557631 317474 557640
rect 317432 557598 317460 557631
rect 317420 557592 317472 557598
rect 317420 557534 317472 557540
rect 317970 553480 318026 553489
rect 317970 553415 317972 553424
rect 318024 553415 318026 553424
rect 317972 553386 318024 553392
rect 316776 552900 316828 552906
rect 316776 552842 316828 552848
rect 316684 551540 316736 551546
rect 316684 551482 316736 551488
rect 314016 550044 314068 550050
rect 314016 549986 314068 549992
rect 317972 549228 318024 549234
rect 317972 549170 318024 549176
rect 317984 549137 318012 549170
rect 317970 549128 318026 549137
rect 317970 549063 318026 549072
rect 312544 545896 312596 545902
rect 312544 545838 312596 545844
rect 313924 545148 313976 545154
rect 313924 545090 313976 545096
rect 311164 544468 311216 544474
rect 311164 544410 311216 544416
rect 307024 540320 307076 540326
rect 307024 540262 307076 540268
rect 305644 519172 305696 519178
rect 305644 519114 305696 519120
rect 307036 518634 307064 540262
rect 312544 540116 312596 540122
rect 312544 540058 312596 540064
rect 307024 518628 307076 518634
rect 307024 518570 307076 518576
rect 312556 518537 312584 540058
rect 312542 518528 312598 518537
rect 312542 518463 312598 518472
rect 313936 515778 313964 545090
rect 314016 544060 314068 544066
rect 314016 544002 314068 544008
rect 314028 515982 314056 544002
rect 314384 543992 314436 543998
rect 314384 543934 314436 543940
rect 314108 543924 314160 543930
rect 314108 543866 314160 543872
rect 314016 515976 314068 515982
rect 314016 515918 314068 515924
rect 314120 515914 314148 543866
rect 314198 541376 314254 541385
rect 314198 541311 314254 541320
rect 314212 517274 314240 541311
rect 314292 540592 314344 540598
rect 314292 540534 314344 540540
rect 314200 517268 314252 517274
rect 314200 517210 314252 517216
rect 314108 515908 314160 515914
rect 314108 515850 314160 515856
rect 314304 515846 314332 540534
rect 314396 520266 314424 543934
rect 317972 543856 318024 543862
rect 317970 543824 317972 543833
rect 318024 543824 318026 543833
rect 316684 543788 316736 543794
rect 317970 543759 318026 543768
rect 316684 543730 316736 543736
rect 314476 540524 314528 540530
rect 314476 540466 314528 540472
rect 314384 520260 314436 520266
rect 314384 520202 314436 520208
rect 314488 517478 314516 540466
rect 314476 517472 314528 517478
rect 314476 517414 314528 517420
rect 314292 515840 314344 515846
rect 314292 515782 314344 515788
rect 313924 515772 313976 515778
rect 313924 515714 313976 515720
rect 304356 515432 304408 515438
rect 304356 515374 304408 515380
rect 316696 514758 316724 543730
rect 318076 543046 318104 630974
rect 318168 555626 318196 632606
rect 318260 558278 318288 632810
rect 318812 592793 318840 634034
rect 337384 632800 337436 632806
rect 337384 632742 337436 632748
rect 319444 632732 319496 632738
rect 319444 632674 319496 632680
rect 319076 630828 319128 630834
rect 319076 630770 319128 630776
rect 319088 629950 319116 630770
rect 319076 629944 319128 629950
rect 319076 629886 319128 629892
rect 318798 592784 318854 592793
rect 318798 592719 318854 592728
rect 318338 562320 318394 562329
rect 318338 562255 318394 562264
rect 318248 558272 318300 558278
rect 318248 558214 318300 558220
rect 318352 556850 318380 562255
rect 318340 556844 318392 556850
rect 318340 556786 318392 556792
rect 318156 555620 318208 555626
rect 318156 555562 318208 555568
rect 319456 545766 319484 632674
rect 319720 632460 319772 632466
rect 319720 632402 319772 632408
rect 319534 632360 319590 632369
rect 319534 632295 319590 632304
rect 319548 547330 319576 632295
rect 319628 632120 319680 632126
rect 319628 632062 319680 632068
rect 319640 552838 319668 632062
rect 319732 559774 319760 632402
rect 332876 632256 332928 632262
rect 332876 632198 332928 632204
rect 320364 632188 320416 632194
rect 320364 632130 320416 632136
rect 319812 631168 319864 631174
rect 319812 631110 319864 631116
rect 319824 589966 319852 631110
rect 320376 630494 320404 632130
rect 323860 632120 323912 632126
rect 323860 632062 323912 632068
rect 323872 630972 323900 632062
rect 332888 630972 332916 632198
rect 337396 630972 337424 632742
rect 364352 632738 364380 702406
rect 400680 641028 400732 641034
rect 400680 640970 400732 640976
rect 396632 633004 396684 633010
rect 396632 632946 396684 632952
rect 378600 632936 378652 632942
rect 378600 632878 378652 632884
rect 355416 632732 355468 632738
rect 355416 632674 355468 632680
rect 364340 632732 364392 632738
rect 364340 632674 364392 632680
rect 350908 632596 350960 632602
rect 350908 632538 350960 632544
rect 341892 632188 341944 632194
rect 341892 632130 341944 632136
rect 341904 630972 341932 632130
rect 346398 632088 346454 632097
rect 346398 632023 346454 632032
rect 346412 630972 346440 632023
rect 350920 630972 350948 632538
rect 355428 630972 355456 632674
rect 359924 632664 359976 632670
rect 359924 632606 359976 632612
rect 359936 630972 359964 632606
rect 364432 632528 364484 632534
rect 364432 632470 364484 632476
rect 364444 630972 364472 632470
rect 373448 632460 373500 632466
rect 373448 632402 373500 632408
rect 368940 631372 368992 631378
rect 368940 631314 368992 631320
rect 368952 630972 368980 631314
rect 373460 630972 373488 632402
rect 378612 630972 378640 632878
rect 383108 632392 383160 632398
rect 383108 632334 383160 632340
rect 392122 632360 392178 632369
rect 383120 630972 383148 632334
rect 387616 632324 387668 632330
rect 392122 632295 392178 632304
rect 387616 632266 387668 632272
rect 387628 630972 387656 632266
rect 392136 630972 392164 632295
rect 396644 630972 396672 632946
rect 400692 630986 400720 640970
rect 428188 632868 428240 632874
rect 428188 632810 428240 632816
rect 423680 632732 423732 632738
rect 423680 632674 423732 632680
rect 414664 632120 414716 632126
rect 414664 632062 414716 632068
rect 414676 630986 414704 632062
rect 419172 631304 419224 631310
rect 419172 631246 419224 631252
rect 400692 630958 401166 630986
rect 414584 630972 414704 630986
rect 419184 630972 419212 631246
rect 423692 630972 423720 632674
rect 428200 630972 428228 632810
rect 414584 630958 414690 630972
rect 328090 630864 328146 630873
rect 328146 630822 328394 630850
rect 328090 630799 328146 630808
rect 409880 630760 409932 630766
rect 405370 630728 405426 630737
rect 405426 630686 405674 630714
rect 409932 630708 410182 630714
rect 409880 630702 410182 630708
rect 409892 630686 410182 630702
rect 414584 630698 414612 630958
rect 414572 630692 414624 630698
rect 405370 630663 405426 630672
rect 414572 630634 414624 630640
rect 320364 630488 320416 630494
rect 320364 630430 320416 630436
rect 319812 589960 319864 589966
rect 319812 589902 319864 589908
rect 319720 559768 319772 559774
rect 319720 559710 319772 559716
rect 428370 558240 428426 558249
rect 428370 558175 428426 558184
rect 319720 555484 319772 555490
rect 319720 555426 319772 555432
rect 319628 552832 319680 552838
rect 319628 552774 319680 552780
rect 319536 547324 319588 547330
rect 319536 547266 319588 547272
rect 319444 545760 319496 545766
rect 319444 545702 319496 545708
rect 318246 543280 318302 543289
rect 318246 543215 318302 543224
rect 319628 543244 319680 543250
rect 318064 543040 318116 543046
rect 318064 542982 318116 542988
rect 317050 542872 317106 542881
rect 317050 542807 317106 542816
rect 316868 541748 316920 541754
rect 316868 541690 316920 541696
rect 316774 541648 316830 541657
rect 316774 541583 316830 541592
rect 316684 514752 316736 514758
rect 316684 514694 316736 514700
rect 316788 514690 316816 541583
rect 316880 515710 316908 541690
rect 316958 541240 317014 541249
rect 316958 541175 317014 541184
rect 316972 516050 317000 541175
rect 317064 517410 317092 542807
rect 318156 542768 318208 542774
rect 318156 542710 318208 542716
rect 317144 541612 317196 541618
rect 317144 541554 317196 541560
rect 317156 518226 317184 541554
rect 317972 541408 318024 541414
rect 317972 541350 318024 541356
rect 317236 540660 317288 540666
rect 317236 540602 317288 540608
rect 317248 520198 317276 540602
rect 317984 538214 318012 541350
rect 318064 539572 318116 539578
rect 318064 539514 318116 539520
rect 318076 539345 318104 539514
rect 318062 539336 318118 539345
rect 318062 539271 318118 539280
rect 317984 538186 318104 538214
rect 317604 535424 317656 535430
rect 317604 535366 317656 535372
rect 317616 534993 317644 535366
rect 317602 534984 317658 534993
rect 317602 534919 317658 534928
rect 317604 529916 317656 529922
rect 317604 529858 317656 529864
rect 317616 529825 317644 529858
rect 317602 529816 317658 529825
rect 317602 529751 317658 529760
rect 317696 525768 317748 525774
rect 317696 525710 317748 525716
rect 317708 525473 317736 525710
rect 317694 525464 317750 525473
rect 317694 525399 317750 525408
rect 317236 520192 317288 520198
rect 317236 520134 317288 520140
rect 318076 518566 318104 538186
rect 318168 519042 318196 542710
rect 318260 520169 318288 543215
rect 319628 543186 319680 543192
rect 319444 543176 319496 543182
rect 319444 543118 319496 543124
rect 318340 541136 318392 541142
rect 318340 541078 318392 541084
rect 318246 520160 318302 520169
rect 318246 520095 318302 520104
rect 318156 519036 318208 519042
rect 318156 518978 318208 518984
rect 318352 518702 318380 541078
rect 318800 540388 318852 540394
rect 318800 540330 318852 540336
rect 318432 540184 318484 540190
rect 318432 540126 318484 540132
rect 318444 518770 318472 540126
rect 318812 520742 318840 540330
rect 319352 540252 319404 540258
rect 319352 540194 319404 540200
rect 319364 524754 319392 540194
rect 319352 524748 319404 524754
rect 319352 524690 319404 524696
rect 319456 524634 319484 543118
rect 319536 541884 319588 541890
rect 319536 541826 319588 541832
rect 319272 524606 319484 524634
rect 319168 523728 319220 523734
rect 319168 523670 319220 523676
rect 318800 520736 318852 520742
rect 318800 520678 318852 520684
rect 318432 518764 318484 518770
rect 318432 518706 318484 518712
rect 318340 518696 318392 518702
rect 318340 518638 318392 518644
rect 318064 518560 318116 518566
rect 318064 518502 318116 518508
rect 319180 518294 319208 523670
rect 319272 519858 319300 524606
rect 319352 524544 319404 524550
rect 319352 524486 319404 524492
rect 319260 519852 319312 519858
rect 319260 519794 319312 519800
rect 319364 518362 319392 524486
rect 319444 524476 319496 524482
rect 319444 524418 319496 524424
rect 319456 519790 319484 524418
rect 319444 519784 319496 519790
rect 319444 519726 319496 519732
rect 319548 518838 319576 541826
rect 319640 541210 319668 543186
rect 319628 541204 319680 541210
rect 319628 541146 319680 541152
rect 319628 541068 319680 541074
rect 319628 541010 319680 541016
rect 319640 523734 319668 541010
rect 319628 523728 319680 523734
rect 319628 523670 319680 523676
rect 319536 518832 319588 518838
rect 319536 518774 319588 518780
rect 319732 518401 319760 555426
rect 319812 541272 319864 541278
rect 319864 541220 319944 541226
rect 319812 541214 319944 541220
rect 319824 541198 319944 541214
rect 319812 541136 319864 541142
rect 319812 541078 319864 541084
rect 319824 524482 319852 541078
rect 319812 524476 319864 524482
rect 319812 524418 319864 524424
rect 319916 520826 319944 541198
rect 319824 520798 319944 520826
rect 319824 518906 319852 520798
rect 319904 520736 319956 520742
rect 319956 520684 320022 520690
rect 319904 520678 320022 520684
rect 319916 520662 320022 520678
rect 427818 520296 427874 520305
rect 356086 520254 356284 520282
rect 324530 520118 324912 520146
rect 324884 518974 324912 520118
rect 328748 520118 329038 520146
rect 333256 520118 333546 520146
rect 337672 520118 338054 520146
rect 342272 520118 342562 520146
rect 346688 520118 347070 520146
rect 351288 520118 351578 520146
rect 324872 518968 324924 518974
rect 324872 518910 324924 518916
rect 319812 518900 319864 518906
rect 319812 518842 319864 518848
rect 328748 518770 328776 520118
rect 333256 518838 333284 520118
rect 333244 518832 333296 518838
rect 333244 518774 333296 518780
rect 328736 518764 328788 518770
rect 328736 518706 328788 518712
rect 337672 518401 337700 520118
rect 319718 518392 319774 518401
rect 319352 518356 319404 518362
rect 319718 518327 319774 518336
rect 337658 518392 337714 518401
rect 337658 518327 337714 518336
rect 319352 518298 319404 518304
rect 319168 518288 319220 518294
rect 319168 518230 319220 518236
rect 342272 518226 342300 520118
rect 346688 518906 346716 520118
rect 351288 519246 351316 520118
rect 351276 519240 351328 519246
rect 351276 519182 351328 519188
rect 346676 518900 346728 518906
rect 346676 518842 346728 518848
rect 356256 518537 356284 520254
rect 427818 520231 427874 520240
rect 360304 520118 360594 520146
rect 364720 520118 365102 520146
rect 369320 520118 369610 520146
rect 374472 520118 374762 520146
rect 378152 520118 379270 520146
rect 383672 520118 383778 520146
rect 387904 520118 388286 520146
rect 391952 520118 392794 520146
rect 396920 520118 397302 520146
rect 401612 520118 401810 520146
rect 406028 520118 406318 520146
rect 410536 520118 410826 520146
rect 414952 520118 415334 520146
rect 419552 520118 419842 520146
rect 423968 520118 424350 520146
rect 356242 518528 356298 518537
rect 356242 518463 356298 518472
rect 360304 518294 360332 520118
rect 364720 518362 364748 520118
rect 369320 519178 369348 520118
rect 369308 519172 369360 519178
rect 369308 519114 369360 519120
rect 374472 518673 374500 520118
rect 374458 518664 374514 518673
rect 374458 518599 374514 518608
rect 364708 518356 364760 518362
rect 364708 518298 364760 518304
rect 360292 518288 360344 518294
rect 360292 518230 360344 518236
rect 317144 518220 317196 518226
rect 317144 518162 317196 518168
rect 342260 518220 342312 518226
rect 342260 518162 342312 518168
rect 317052 517404 317104 517410
rect 317052 517346 317104 517352
rect 316960 516044 317012 516050
rect 316960 515986 317012 515992
rect 316868 515704 316920 515710
rect 316868 515646 316920 515652
rect 316776 514684 316828 514690
rect 316776 514626 316828 514632
rect 302238 502480 302294 502489
rect 302238 502415 302294 502424
rect 302882 487520 302938 487529
rect 302882 487455 302938 487464
rect 302896 487218 302924 487455
rect 302884 487212 302936 487218
rect 302884 487154 302936 487160
rect 366362 480856 366418 480865
rect 366362 480791 366418 480800
rect 59740 480134 60214 480162
rect 299782 480134 299888 480162
rect 59740 480094 59768 480134
rect 59648 480066 59768 480094
rect 158720 480072 158772 480078
rect 50988 478984 51040 478990
rect 50988 478926 51040 478932
rect 50896 478780 50948 478786
rect 50896 478722 50948 478728
rect 50068 478644 50120 478650
rect 50068 478586 50120 478592
rect 43812 478168 43864 478174
rect 43812 478110 43864 478116
rect 43720 470212 43772 470218
rect 43720 470154 43772 470160
rect 43444 469872 43496 469878
rect 43444 469814 43496 469820
rect 43260 460692 43312 460698
rect 43260 460634 43312 460640
rect 42708 382220 42760 382226
rect 42708 382162 42760 382168
rect 43272 373833 43300 460634
rect 43352 460624 43404 460630
rect 43352 460566 43404 460572
rect 43258 373824 43314 373833
rect 43258 373759 43314 373768
rect 43364 371210 43392 460566
rect 43456 373726 43484 469814
rect 43628 468716 43680 468722
rect 43628 468658 43680 468664
rect 43536 465724 43588 465730
rect 43536 465666 43588 465672
rect 43444 373720 43496 373726
rect 43444 373662 43496 373668
rect 43352 371204 43404 371210
rect 43352 371146 43404 371152
rect 43548 269550 43576 465666
rect 43536 269544 43588 269550
rect 43536 269486 43588 269492
rect 43640 267714 43668 468658
rect 43628 267708 43680 267714
rect 43628 267650 43680 267656
rect 43732 264858 43760 470154
rect 43824 267578 43852 478110
rect 48044 475992 48096 475998
rect 46846 475960 46902 475969
rect 48044 475934 48096 475940
rect 46846 475895 46902 475904
rect 46388 475652 46440 475658
rect 46388 475594 46440 475600
rect 45468 473136 45520 473142
rect 45468 473078 45520 473084
rect 43994 472968 44050 472977
rect 43994 472903 44050 472912
rect 43904 470348 43956 470354
rect 43904 470290 43956 470296
rect 43812 267572 43864 267578
rect 43812 267514 43864 267520
rect 43720 264852 43772 264858
rect 43720 264794 43772 264800
rect 43916 249762 43944 470290
rect 43904 249756 43956 249762
rect 43904 249698 43956 249704
rect 44008 173874 44036 472903
rect 45376 468648 45428 468654
rect 45376 468590 45428 468596
rect 45284 468580 45336 468586
rect 45284 468522 45336 468528
rect 45192 467220 45244 467226
rect 45192 467162 45244 467168
rect 45008 465860 45060 465866
rect 45008 465802 45060 465808
rect 44732 465588 44784 465594
rect 44732 465530 44784 465536
rect 44088 460216 44140 460222
rect 44088 460158 44140 460164
rect 43996 173868 44048 173874
rect 43996 173810 44048 173816
rect 42616 58812 42668 58818
rect 42616 58754 42668 58760
rect 44100 57798 44128 460158
rect 44640 409896 44692 409902
rect 44640 409838 44692 409844
rect 44652 373998 44680 409838
rect 44640 373992 44692 373998
rect 44640 373934 44692 373940
rect 44744 371958 44772 465530
rect 44824 465520 44876 465526
rect 44824 465462 44876 465468
rect 44732 371952 44784 371958
rect 44732 371894 44784 371900
rect 44836 371278 44864 465462
rect 44916 460420 44968 460426
rect 44916 460362 44968 460368
rect 44824 371272 44876 371278
rect 44824 371214 44876 371220
rect 44928 269482 44956 460362
rect 44916 269476 44968 269482
rect 44916 269418 44968 269424
rect 45020 269414 45048 465802
rect 45100 465792 45152 465798
rect 45100 465734 45152 465740
rect 45008 269408 45060 269414
rect 45008 269350 45060 269356
rect 45112 269346 45140 465734
rect 45204 269754 45232 467162
rect 45192 269748 45244 269754
rect 45192 269690 45244 269696
rect 45100 269340 45152 269346
rect 45100 269282 45152 269288
rect 45296 269210 45324 468522
rect 45388 269278 45416 468590
rect 45376 269272 45428 269278
rect 45376 269214 45428 269220
rect 45284 269204 45336 269210
rect 45284 269146 45336 269152
rect 45480 269074 45508 473078
rect 46296 472728 46348 472734
rect 46296 472670 46348 472676
rect 46112 472660 46164 472666
rect 46112 472602 46164 472608
rect 46020 458312 46072 458318
rect 46020 458254 46072 458260
rect 46032 412622 46060 458254
rect 46020 412616 46072 412622
rect 46020 412558 46072 412564
rect 46124 385014 46152 472602
rect 46204 469940 46256 469946
rect 46204 469882 46256 469888
rect 46112 385008 46164 385014
rect 46112 384950 46164 384956
rect 46216 373590 46244 469882
rect 46204 373584 46256 373590
rect 46204 373526 46256 373532
rect 46308 373318 46336 472670
rect 46296 373312 46348 373318
rect 46296 373254 46348 373260
rect 46296 371272 46348 371278
rect 46296 371214 46348 371220
rect 46204 269680 46256 269686
rect 46204 269622 46256 269628
rect 45468 269068 45520 269074
rect 45468 269010 45520 269016
rect 46216 145586 46244 269622
rect 46308 267481 46336 371214
rect 46400 268122 46428 475594
rect 46478 475552 46534 475561
rect 46478 475487 46534 475496
rect 46756 475516 46808 475522
rect 46492 268938 46520 475487
rect 46756 475458 46808 475464
rect 46572 473272 46624 473278
rect 46572 473214 46624 473220
rect 46480 268932 46532 268938
rect 46480 268874 46532 268880
rect 46388 268116 46440 268122
rect 46388 268058 46440 268064
rect 46294 267472 46350 267481
rect 46294 267407 46350 267416
rect 46308 266393 46336 267407
rect 46294 266384 46350 266393
rect 46294 266319 46350 266328
rect 46204 145580 46256 145586
rect 46204 145522 46256 145528
rect 46400 145382 46428 268058
rect 46478 266384 46534 266393
rect 46478 266319 46534 266328
rect 46492 148646 46520 266319
rect 46584 264518 46612 473214
rect 46664 472592 46716 472598
rect 46664 472534 46716 472540
rect 46676 264586 46704 472534
rect 46768 264654 46796 475458
rect 46756 264648 46808 264654
rect 46756 264590 46808 264596
rect 46664 264580 46716 264586
rect 46664 264522 46716 264528
rect 46572 264512 46624 264518
rect 46572 264454 46624 264460
rect 46480 148640 46532 148646
rect 46480 148582 46532 148588
rect 46388 145376 46440 145382
rect 46388 145318 46440 145324
rect 46860 69018 46888 475895
rect 47860 475720 47912 475726
rect 47860 475662 47912 475668
rect 47768 472796 47820 472802
rect 47768 472738 47820 472744
rect 47584 462868 47636 462874
rect 47584 462810 47636 462816
rect 47492 408536 47544 408542
rect 47492 408478 47544 408484
rect 47400 407176 47452 407182
rect 47400 407118 47452 407124
rect 47412 373930 47440 407118
rect 47504 375057 47532 408478
rect 47490 375048 47546 375057
rect 47490 374983 47546 374992
rect 47400 373924 47452 373930
rect 47400 373866 47452 373872
rect 47596 371890 47624 462810
rect 47676 462800 47728 462806
rect 47676 462742 47728 462748
rect 47688 372026 47716 462742
rect 47780 373862 47808 472738
rect 47768 373856 47820 373862
rect 47768 373798 47820 373804
rect 47676 372020 47728 372026
rect 47676 371962 47728 371968
rect 47584 371884 47636 371890
rect 47584 371826 47636 371832
rect 47596 364334 47624 371826
rect 47688 370138 47716 371962
rect 47688 370110 47808 370138
rect 47596 364306 47716 364334
rect 47688 266558 47716 364306
rect 47780 266830 47808 370110
rect 47872 298110 47900 475662
rect 47952 468988 48004 468994
rect 47952 468930 48004 468936
rect 47860 298104 47912 298110
rect 47860 298046 47912 298052
rect 47964 266937 47992 468930
rect 48056 268598 48084 475934
rect 49056 475924 49108 475930
rect 49056 475866 49108 475872
rect 48136 475788 48188 475794
rect 48136 475730 48188 475736
rect 48044 268592 48096 268598
rect 48044 268534 48096 268540
rect 48148 268258 48176 475730
rect 48964 475584 49016 475590
rect 48964 475526 49016 475532
rect 48228 473340 48280 473346
rect 48228 473282 48280 473288
rect 48136 268252 48188 268258
rect 48136 268194 48188 268200
rect 47950 266928 48006 266937
rect 47950 266863 48006 266872
rect 48044 266892 48096 266898
rect 48044 266834 48096 266840
rect 47768 266824 47820 266830
rect 47768 266766 47820 266772
rect 47676 266552 47728 266558
rect 47676 266494 47728 266500
rect 47780 146266 47808 266766
rect 48056 266558 48084 266834
rect 48044 266552 48096 266558
rect 48044 266494 48096 266500
rect 47952 264988 48004 264994
rect 47952 264930 48004 264936
rect 47858 249112 47914 249121
rect 47858 249047 47914 249056
rect 47872 160750 47900 249047
rect 47964 163810 47992 264930
rect 47952 163804 48004 163810
rect 47952 163746 48004 163752
rect 47860 160744 47912 160750
rect 47860 160686 47912 160692
rect 48056 148714 48084 266494
rect 48044 148708 48096 148714
rect 48044 148650 48096 148656
rect 47768 146260 47820 146266
rect 47768 146202 47820 146208
rect 48148 145450 48176 268194
rect 48240 264722 48268 473282
rect 48872 472864 48924 472870
rect 48872 472806 48924 472812
rect 48780 470008 48832 470014
rect 48780 469950 48832 469956
rect 48792 373454 48820 469950
rect 48780 373448 48832 373454
rect 48780 373390 48832 373396
rect 48884 373182 48912 472806
rect 48872 373176 48924 373182
rect 48872 373118 48924 373124
rect 48872 371952 48924 371958
rect 48872 371894 48924 371900
rect 48884 371550 48912 371894
rect 48872 371544 48924 371550
rect 48872 371486 48924 371492
rect 48884 267345 48912 371486
rect 48976 268054 49004 475526
rect 49068 268462 49096 475866
rect 49148 475448 49200 475454
rect 49148 475390 49200 475396
rect 49056 268456 49108 268462
rect 49056 268398 49108 268404
rect 48964 268048 49016 268054
rect 48964 267990 49016 267996
rect 48870 267336 48926 267345
rect 48870 267271 48926 267280
rect 48884 266393 48912 267271
rect 48870 266384 48926 266393
rect 48870 266319 48926 266328
rect 48228 264716 48280 264722
rect 48228 264658 48280 264664
rect 48976 145790 49004 267990
rect 49160 267306 49188 475390
rect 49240 473204 49292 473210
rect 49240 473146 49292 473152
rect 49148 267300 49200 267306
rect 49148 267242 49200 267248
rect 49146 266384 49202 266393
rect 49146 266319 49202 266328
rect 49160 148578 49188 266319
rect 49252 264790 49280 473146
rect 49424 466336 49476 466342
rect 49424 466278 49476 466284
rect 49332 463616 49384 463622
rect 49332 463558 49384 463564
rect 49240 264784 49292 264790
rect 49240 264726 49292 264732
rect 49148 148572 49200 148578
rect 49148 148514 49200 148520
rect 48964 145784 49016 145790
rect 48964 145726 49016 145732
rect 48136 145444 48188 145450
rect 48136 145386 48188 145392
rect 49252 144634 49280 264726
rect 49344 162042 49372 463558
rect 49436 164014 49464 466278
rect 49516 460556 49568 460562
rect 49516 460498 49568 460504
rect 49424 164008 49476 164014
rect 49424 163950 49476 163956
rect 49332 162036 49384 162042
rect 49332 161978 49384 161984
rect 49240 144628 49292 144634
rect 49240 144570 49292 144576
rect 46848 69012 46900 69018
rect 46848 68954 46900 68960
rect 49528 59430 49556 460498
rect 49608 460352 49660 460358
rect 49608 460294 49660 460300
rect 49516 59424 49568 59430
rect 49516 59366 49568 59372
rect 44088 57792 44140 57798
rect 44088 57734 44140 57740
rect 39948 57520 40000 57526
rect 39948 57462 40000 57468
rect 49620 55894 49648 460294
rect 50080 58750 50108 478586
rect 50908 477601 50936 478722
rect 50894 477592 50950 477601
rect 50894 477527 50950 477536
rect 50342 475688 50398 475697
rect 50342 475623 50398 475632
rect 50160 472932 50212 472938
rect 50160 472874 50212 472880
rect 50172 373386 50200 472874
rect 50252 465996 50304 466002
rect 50252 465938 50304 465944
rect 50160 373380 50212 373386
rect 50160 373322 50212 373328
rect 50264 267034 50292 465938
rect 50356 269074 50384 475623
rect 50436 472524 50488 472530
rect 50436 472466 50488 472472
rect 50344 269068 50396 269074
rect 50344 269010 50396 269016
rect 50252 267028 50304 267034
rect 50252 266970 50304 266976
rect 50344 266416 50396 266422
rect 50344 266358 50396 266364
rect 50356 144702 50384 266358
rect 50448 265742 50476 472466
rect 51000 470594 51028 478926
rect 52092 478916 52144 478922
rect 52092 478858 52144 478864
rect 52000 478304 52052 478310
rect 52000 478246 52052 478252
rect 51908 476060 51960 476066
rect 51908 476002 51960 476008
rect 50908 470566 51028 470594
rect 50620 466404 50672 466410
rect 50620 466346 50672 466352
rect 50528 460284 50580 460290
rect 50528 460226 50580 460232
rect 50436 265736 50488 265742
rect 50436 265678 50488 265684
rect 50540 162858 50568 460226
rect 50632 164694 50660 466346
rect 50802 466032 50858 466041
rect 50802 465967 50858 465976
rect 50712 460896 50764 460902
rect 50712 460838 50764 460844
rect 50724 459649 50752 460838
rect 50710 459640 50766 459649
rect 50710 459575 50766 459584
rect 50712 456136 50764 456142
rect 50712 456078 50764 456084
rect 50620 164688 50672 164694
rect 50620 164630 50672 164636
rect 50528 162852 50580 162858
rect 50528 162794 50580 162800
rect 50724 162625 50752 456078
rect 50816 163742 50844 465967
rect 50908 163946 50936 470566
rect 51540 470076 51592 470082
rect 51540 470018 51592 470024
rect 50986 463040 51042 463049
rect 50986 462975 51042 462984
rect 51000 456142 51028 462975
rect 50988 456136 51040 456142
rect 50988 456078 51040 456084
rect 51552 373658 51580 470018
rect 51816 466200 51868 466206
rect 51816 466142 51868 466148
rect 51724 459060 51776 459066
rect 51724 459002 51776 459008
rect 51632 404388 51684 404394
rect 51632 404330 51684 404336
rect 51644 375086 51672 404330
rect 51736 404326 51764 459002
rect 51724 404320 51776 404326
rect 51724 404262 51776 404268
rect 51724 379568 51776 379574
rect 51724 379510 51776 379516
rect 51632 375080 51684 375086
rect 51632 375022 51684 375028
rect 51540 373652 51592 373658
rect 51540 373594 51592 373600
rect 51632 372632 51684 372638
rect 51632 372574 51684 372580
rect 51448 269816 51500 269822
rect 51448 269758 51500 269764
rect 50986 268424 51042 268433
rect 50986 268359 51042 268368
rect 51000 267510 51028 268359
rect 51460 268274 51488 269758
rect 51540 269612 51592 269618
rect 51540 269554 51592 269560
rect 51552 268394 51580 269554
rect 51540 268388 51592 268394
rect 51540 268330 51592 268336
rect 51460 268246 51580 268274
rect 51448 267776 51500 267782
rect 51448 267718 51500 267724
rect 50988 267504 51040 267510
rect 50988 267446 51040 267452
rect 51000 266422 51028 267446
rect 50988 266416 51040 266422
rect 50988 266358 51040 266364
rect 50896 163940 50948 163946
rect 50896 163882 50948 163888
rect 50804 163736 50856 163742
rect 50804 163678 50856 163684
rect 50710 162616 50766 162625
rect 50710 162551 50766 162560
rect 51460 160886 51488 267718
rect 51448 160880 51500 160886
rect 51448 160822 51500 160828
rect 51552 144809 51580 268246
rect 51644 264926 51672 372574
rect 51736 269618 51764 379510
rect 51724 269612 51776 269618
rect 51724 269554 51776 269560
rect 51724 269068 51776 269074
rect 51724 269010 51776 269016
rect 51736 267782 51764 269010
rect 51724 267776 51776 267782
rect 51724 267718 51776 267724
rect 51828 267170 51856 466142
rect 51920 268530 51948 476002
rect 51908 268524 51960 268530
rect 51908 268466 51960 268472
rect 52012 267238 52040 478246
rect 52000 267232 52052 267238
rect 52000 267174 52052 267180
rect 51816 267164 51868 267170
rect 51816 267106 51868 267112
rect 52104 267102 52132 478858
rect 54576 478848 54628 478854
rect 54576 478790 54628 478796
rect 52828 478508 52880 478514
rect 52828 478450 52880 478456
rect 52276 465656 52328 465662
rect 52276 465598 52328 465604
rect 52184 461644 52236 461650
rect 52184 461586 52236 461592
rect 52092 267096 52144 267102
rect 52092 267038 52144 267044
rect 51908 266212 51960 266218
rect 51908 266154 51960 266160
rect 51632 264920 51684 264926
rect 51632 264862 51684 264868
rect 51816 146260 51868 146266
rect 51816 146202 51868 146208
rect 51828 145518 51856 146202
rect 51816 145512 51868 145518
rect 51816 145454 51868 145460
rect 51538 144800 51594 144809
rect 51538 144735 51594 144744
rect 50344 144696 50396 144702
rect 50344 144638 50396 144644
rect 50068 58744 50120 58750
rect 50068 58686 50120 58692
rect 51828 57254 51856 145454
rect 51920 144770 51948 266154
rect 52000 265872 52052 265878
rect 52000 265814 52052 265820
rect 52012 144838 52040 265814
rect 52196 163878 52224 461586
rect 52288 164082 52316 465598
rect 52368 403028 52420 403034
rect 52368 402970 52420 402976
rect 52380 375442 52408 402970
rect 52380 375414 52500 375442
rect 52366 375320 52422 375329
rect 52366 375255 52422 375264
rect 52276 164076 52328 164082
rect 52276 164018 52328 164024
rect 52184 163872 52236 163878
rect 52184 163814 52236 163820
rect 52276 163804 52328 163810
rect 52276 163746 52328 163752
rect 52288 162994 52316 163746
rect 52276 162988 52328 162994
rect 52276 162930 52328 162936
rect 52092 148708 52144 148714
rect 52092 148650 52144 148656
rect 52000 144832 52052 144838
rect 52000 144774 52052 144780
rect 51908 144764 51960 144770
rect 51908 144706 51960 144712
rect 51816 57248 51868 57254
rect 51816 57190 51868 57196
rect 52104 55962 52132 148650
rect 52184 148368 52236 148374
rect 52184 148310 52236 148316
rect 52092 55956 52144 55962
rect 52092 55898 52144 55904
rect 49608 55888 49660 55894
rect 49608 55830 49660 55836
rect 52196 55010 52224 148310
rect 52288 55146 52316 162930
rect 52380 57866 52408 375255
rect 52472 374921 52500 375414
rect 52458 374912 52514 374921
rect 52458 374847 52514 374856
rect 52368 57860 52420 57866
rect 52368 57802 52420 57808
rect 52840 57730 52868 478450
rect 53472 478372 53524 478378
rect 53472 478314 53524 478320
rect 53484 477601 53512 478314
rect 53470 477592 53526 477601
rect 53470 477527 53526 477536
rect 53564 473068 53616 473074
rect 53564 473010 53616 473016
rect 53470 466168 53526 466177
rect 53196 466132 53248 466138
rect 53470 466103 53526 466112
rect 53196 466074 53248 466080
rect 53104 466064 53156 466070
rect 53104 466006 53156 466012
rect 53012 463004 53064 463010
rect 53012 462946 53064 462952
rect 52920 458856 52972 458862
rect 52920 458798 52972 458804
rect 52932 269618 52960 458798
rect 52920 269612 52972 269618
rect 52920 269554 52972 269560
rect 53024 267306 53052 462946
rect 53116 267442 53144 466006
rect 53104 267436 53156 267442
rect 53104 267378 53156 267384
rect 53208 267374 53236 466074
rect 53288 463412 53340 463418
rect 53288 463354 53340 463360
rect 53196 267368 53248 267374
rect 53196 267310 53248 267316
rect 52920 267300 52972 267306
rect 52920 267242 52972 267248
rect 53012 267300 53064 267306
rect 53012 267242 53064 267248
rect 52932 267073 52960 267242
rect 52918 267064 52974 267073
rect 52918 266999 52974 267008
rect 52932 161022 52960 266999
rect 53104 265736 53156 265742
rect 53104 265678 53156 265684
rect 53116 264586 53144 265678
rect 53104 264580 53156 264586
rect 53104 264522 53156 264528
rect 52920 161016 52972 161022
rect 52920 160958 52972 160964
rect 53116 146198 53144 264522
rect 53196 163056 53248 163062
rect 53196 162998 53248 163004
rect 53104 146192 53156 146198
rect 53104 146134 53156 146140
rect 52828 57724 52880 57730
rect 52828 57666 52880 57672
rect 52276 55140 52328 55146
rect 52276 55082 52328 55088
rect 52184 55004 52236 55010
rect 52184 54946 52236 54952
rect 53116 54942 53144 146134
rect 53208 56506 53236 162998
rect 53300 162314 53328 463354
rect 53380 463072 53432 463078
rect 53380 463014 53432 463020
rect 53392 162382 53420 463014
rect 53380 162376 53432 162382
rect 53380 162318 53432 162324
rect 53288 162308 53340 162314
rect 53288 162250 53340 162256
rect 53484 162110 53512 466103
rect 53576 409834 53604 473010
rect 54392 470484 54444 470490
rect 54392 470426 54444 470432
rect 53748 460828 53800 460834
rect 53748 460770 53800 460776
rect 53656 460760 53708 460766
rect 53656 460702 53708 460708
rect 53564 409828 53616 409834
rect 53564 409770 53616 409776
rect 53564 405748 53616 405754
rect 53564 405690 53616 405696
rect 53576 375426 53604 405690
rect 53564 375420 53616 375426
rect 53564 375362 53616 375368
rect 53562 375320 53618 375329
rect 53562 375255 53618 375264
rect 53472 162104 53524 162110
rect 53472 162046 53524 162052
rect 53380 148640 53432 148646
rect 53380 148582 53432 148588
rect 53288 148572 53340 148578
rect 53288 148514 53340 148520
rect 53196 56500 53248 56506
rect 53196 56442 53248 56448
rect 53300 56030 53328 148514
rect 53288 56024 53340 56030
rect 53288 55966 53340 55972
rect 53104 54936 53156 54942
rect 53104 54878 53156 54884
rect 53392 54670 53420 148582
rect 53576 58682 53604 375255
rect 53564 58676 53616 58682
rect 53564 58618 53616 58624
rect 53668 57390 53696 460702
rect 53760 459649 53788 460770
rect 53746 459640 53802 459649
rect 53746 459575 53802 459584
rect 54404 414254 54432 470426
rect 54484 458924 54536 458930
rect 54484 458866 54536 458872
rect 54392 414248 54444 414254
rect 54392 414190 54444 414196
rect 54392 411936 54444 411942
rect 54392 411878 54444 411884
rect 53840 404320 53892 404326
rect 53840 404262 53892 404268
rect 53852 379574 53880 404262
rect 53840 379568 53892 379574
rect 53840 379510 53892 379516
rect 53748 375352 53800 375358
rect 53748 375294 53800 375300
rect 53760 375018 53788 375294
rect 53748 375012 53800 375018
rect 53748 374954 53800 374960
rect 54404 372638 54432 411878
rect 54496 374066 54524 458866
rect 54484 374060 54536 374066
rect 54484 374002 54536 374008
rect 54392 372632 54444 372638
rect 54392 372574 54444 372580
rect 54588 371142 54616 478790
rect 56416 478712 56468 478718
rect 56416 478654 56468 478660
rect 56324 478440 56376 478446
rect 56324 478382 56376 478388
rect 54760 475312 54812 475318
rect 54760 475254 54812 475260
rect 54668 459128 54720 459134
rect 54668 459070 54720 459076
rect 54576 371136 54628 371142
rect 54576 371078 54628 371084
rect 54576 369572 54628 369578
rect 54576 369514 54628 369520
rect 54484 368688 54536 368694
rect 54484 368630 54536 368636
rect 54392 352572 54444 352578
rect 54392 352514 54444 352520
rect 54404 270494 54432 352514
rect 54312 270466 54432 270494
rect 54312 269498 54340 270466
rect 54496 269822 54524 368630
rect 54484 269816 54536 269822
rect 54484 269758 54536 269764
rect 54312 269470 54432 269498
rect 54404 269113 54432 269470
rect 54588 269226 54616 369514
rect 54496 269198 54616 269226
rect 54390 269104 54446 269113
rect 54390 269039 54446 269048
rect 53746 268560 53802 268569
rect 53746 268495 53802 268504
rect 53760 268394 53788 268495
rect 53748 268388 53800 268394
rect 53748 268330 53800 268336
rect 53760 146305 53788 268330
rect 54208 268184 54260 268190
rect 54208 268126 54260 268132
rect 54220 267850 54248 268126
rect 54300 267980 54352 267986
rect 54300 267922 54352 267928
rect 54208 267844 54260 267850
rect 54208 267786 54260 267792
rect 54220 161294 54248 267786
rect 54208 161288 54260 161294
rect 54208 161230 54260 161236
rect 54312 160954 54340 267922
rect 54404 165578 54432 269039
rect 54496 268190 54524 269198
rect 54680 269090 54708 459070
rect 54588 269062 54708 269090
rect 54484 268184 54536 268190
rect 54484 268126 54536 268132
rect 54588 266286 54616 269062
rect 54668 268932 54720 268938
rect 54668 268874 54720 268880
rect 54680 267986 54708 268874
rect 54668 267980 54720 267986
rect 54668 267922 54720 267928
rect 54772 266966 54800 475254
rect 55862 472560 55918 472569
rect 55862 472495 55918 472504
rect 55680 470552 55732 470558
rect 55680 470494 55732 470500
rect 54944 463480 54996 463486
rect 54944 463422 54996 463428
rect 54852 462936 54904 462942
rect 54852 462878 54904 462884
rect 54760 266960 54812 266966
rect 54760 266902 54812 266908
rect 54576 266280 54628 266286
rect 54576 266222 54628 266228
rect 54484 266076 54536 266082
rect 54484 266018 54536 266024
rect 54496 264654 54524 266018
rect 54576 265940 54628 265946
rect 54576 265882 54628 265888
rect 54484 264648 54536 264654
rect 54484 264590 54536 264596
rect 54392 165572 54444 165578
rect 54392 165514 54444 165520
rect 54300 160948 54352 160954
rect 54300 160890 54352 160896
rect 53746 146296 53802 146305
rect 53746 146231 53802 146240
rect 54392 145784 54444 145790
rect 54392 145726 54444 145732
rect 54404 59566 54432 145726
rect 54496 144906 54524 264590
rect 54588 264518 54616 265882
rect 54576 264512 54628 264518
rect 54576 264454 54628 264460
rect 54588 161474 54616 264454
rect 54864 161906 54892 462878
rect 54956 162518 54984 463422
rect 55128 463344 55180 463350
rect 55128 463286 55180 463292
rect 55036 463276 55088 463282
rect 55036 463218 55088 463224
rect 55048 162586 55076 463218
rect 55140 162722 55168 463286
rect 55692 415313 55720 470494
rect 55772 458992 55824 458998
rect 55772 458934 55824 458940
rect 55678 415304 55734 415313
rect 55678 415239 55734 415248
rect 55588 414248 55640 414254
rect 55588 414190 55640 414196
rect 55494 375320 55550 375329
rect 55494 375255 55550 375264
rect 55220 269816 55272 269822
rect 55220 269758 55272 269764
rect 55232 268394 55260 269758
rect 55220 268388 55272 268394
rect 55220 268330 55272 268336
rect 55128 162716 55180 162722
rect 55128 162658 55180 162664
rect 55036 162580 55088 162586
rect 55036 162522 55088 162528
rect 54944 162512 54996 162518
rect 54944 162454 54996 162460
rect 54852 161900 54904 161906
rect 54852 161842 54904 161848
rect 54588 161446 54892 161474
rect 54760 148504 54812 148510
rect 54760 148446 54812 148452
rect 54576 145444 54628 145450
rect 54576 145386 54628 145392
rect 54484 144900 54536 144906
rect 54484 144842 54536 144848
rect 54588 59634 54616 145386
rect 54668 145376 54720 145382
rect 54668 145318 54720 145324
rect 54576 59628 54628 59634
rect 54576 59570 54628 59576
rect 54392 59560 54444 59566
rect 54392 59502 54444 59508
rect 53656 57384 53708 57390
rect 53656 57326 53708 57332
rect 54680 57186 54708 145318
rect 54772 58886 54800 148446
rect 54864 145994 54892 161446
rect 55036 161288 55088 161294
rect 55036 161230 55088 161236
rect 54944 148436 54996 148442
rect 54944 148378 54996 148384
rect 54852 145988 54904 145994
rect 54852 145930 54904 145936
rect 54760 58880 54812 58886
rect 54760 58822 54812 58828
rect 54668 57180 54720 57186
rect 54668 57122 54720 57128
rect 54864 56098 54892 145930
rect 54956 57662 54984 148378
rect 55048 59498 55076 161230
rect 55128 160880 55180 160886
rect 55128 160822 55180 160828
rect 55036 59492 55088 59498
rect 55036 59434 55088 59440
rect 54944 57656 54996 57662
rect 54944 57598 54996 57604
rect 55140 57458 55168 160822
rect 55128 57452 55180 57458
rect 55128 57394 55180 57400
rect 55508 57322 55536 375255
rect 55600 373017 55628 414190
rect 55784 373114 55812 458934
rect 55772 373108 55824 373114
rect 55772 373050 55824 373056
rect 55586 373008 55642 373017
rect 55586 372943 55642 372952
rect 55678 372736 55734 372745
rect 55678 372671 55734 372680
rect 55692 278730 55720 372671
rect 55876 368694 55904 472495
rect 56048 463684 56100 463690
rect 56048 463626 56100 463632
rect 55956 459264 56008 459270
rect 55956 459206 56008 459212
rect 55864 368688 55916 368694
rect 55864 368630 55916 368636
rect 55864 353388 55916 353394
rect 55864 353330 55916 353336
rect 55680 278724 55732 278730
rect 55680 278666 55732 278672
rect 55876 267510 55904 353330
rect 55864 267504 55916 267510
rect 55864 267446 55916 267452
rect 55772 266348 55824 266354
rect 55772 266290 55824 266296
rect 55680 164620 55732 164626
rect 55680 164562 55732 164568
rect 55496 57316 55548 57322
rect 55496 57258 55548 57264
rect 54852 56092 54904 56098
rect 54852 56034 54904 56040
rect 55692 55078 55720 164562
rect 55784 162926 55812 266290
rect 55864 266280 55916 266286
rect 55864 266222 55916 266228
rect 55876 265810 55904 266222
rect 55864 265804 55916 265810
rect 55864 265746 55916 265752
rect 55772 162920 55824 162926
rect 55772 162862 55824 162868
rect 55784 55214 55812 162862
rect 55876 161474 55904 265746
rect 55968 164490 55996 459206
rect 55956 164484 56008 164490
rect 55956 164426 56008 164432
rect 56060 162246 56088 463626
rect 56232 463548 56284 463554
rect 56232 463490 56284 463496
rect 56140 463208 56192 463214
rect 56140 463150 56192 463156
rect 56152 162790 56180 463150
rect 56140 162784 56192 162790
rect 56140 162726 56192 162732
rect 56244 162450 56272 463490
rect 56336 162654 56364 478382
rect 56324 162648 56376 162654
rect 56324 162590 56376 162596
rect 56232 162444 56284 162450
rect 56232 162386 56284 162392
rect 56048 162240 56100 162246
rect 56048 162182 56100 162188
rect 56428 161974 56456 478654
rect 59176 478576 59228 478582
rect 59176 478518 59228 478524
rect 58808 475244 58860 475250
rect 58808 475186 58860 475192
rect 57336 475108 57388 475114
rect 57336 475050 57388 475056
rect 57060 473000 57112 473006
rect 57060 472942 57112 472948
rect 56508 466268 56560 466274
rect 56508 466210 56560 466216
rect 56520 374950 56548 466210
rect 56968 412616 57020 412622
rect 56968 412558 57020 412564
rect 56980 412321 57008 412558
rect 56966 412312 57022 412321
rect 56966 412247 57022 412256
rect 57072 410854 57100 472942
rect 57244 471368 57296 471374
rect 57244 471310 57296 471316
rect 57152 470416 57204 470422
rect 57152 470358 57204 470364
rect 57060 410848 57112 410854
rect 57060 410790 57112 410796
rect 57058 410408 57114 410417
rect 57058 410343 57114 410352
rect 57072 409902 57100 410343
rect 57060 409896 57112 409902
rect 57060 409838 57112 409844
rect 56876 409828 56928 409834
rect 56876 409770 56928 409776
rect 56888 404274 56916 409770
rect 57058 408640 57114 408649
rect 57058 408575 57114 408584
rect 57072 408542 57100 408575
rect 57060 408536 57112 408542
rect 57060 408478 57112 408484
rect 56966 407416 57022 407425
rect 56966 407351 57022 407360
rect 56980 407182 57008 407351
rect 56968 407176 57020 407182
rect 56968 407118 57020 407124
rect 57058 405784 57114 405793
rect 57058 405719 57060 405728
rect 57112 405719 57114 405728
rect 57060 405690 57112 405696
rect 57058 404424 57114 404433
rect 57058 404359 57060 404368
rect 57112 404359 57114 404368
rect 57060 404330 57112 404336
rect 56888 404246 57100 404274
rect 56966 403064 57022 403073
rect 56966 402999 56968 403008
rect 57020 402999 57022 403008
rect 56968 402970 57020 402976
rect 56968 385008 57020 385014
rect 56966 384976 56968 384985
rect 57020 384976 57022 384985
rect 56966 384911 57022 384920
rect 56968 383648 57020 383654
rect 56968 383590 57020 383596
rect 56874 383344 56930 383353
rect 56874 383279 56930 383288
rect 56888 382226 56916 383279
rect 56876 382220 56928 382226
rect 56876 382162 56928 382168
rect 56508 374944 56560 374950
rect 56508 374886 56560 374892
rect 56980 374134 57008 383590
rect 56968 374128 57020 374134
rect 56968 374070 57020 374076
rect 57072 373250 57100 404246
rect 57164 383654 57192 470358
rect 57256 383654 57284 471310
rect 57348 383654 57376 475050
rect 57888 474020 57940 474026
rect 57888 473962 57940 473968
rect 57796 467288 57848 467294
rect 57796 467230 57848 467236
rect 57428 464432 57480 464438
rect 57428 464374 57480 464380
rect 57152 383648 57204 383654
rect 57152 383590 57204 383596
rect 57244 383648 57296 383654
rect 57244 383590 57296 383596
rect 57336 383648 57388 383654
rect 57336 383590 57388 383596
rect 57152 383512 57204 383518
rect 57152 383454 57204 383460
rect 57244 383512 57296 383518
rect 57440 383466 57468 464374
rect 57612 463140 57664 463146
rect 57612 463082 57664 463088
rect 57520 459196 57572 459202
rect 57520 459138 57572 459144
rect 57244 383454 57296 383460
rect 57164 383081 57192 383454
rect 57150 383072 57206 383081
rect 57150 383007 57206 383016
rect 57256 382378 57284 383454
rect 57164 382350 57284 382378
rect 57348 383438 57468 383466
rect 57164 378622 57192 382350
rect 57244 382220 57296 382226
rect 57244 382162 57296 382168
rect 57152 378616 57204 378622
rect 57152 378558 57204 378564
rect 57060 373244 57112 373250
rect 57060 373186 57112 373192
rect 56506 372872 56562 372881
rect 56506 372807 56562 372816
rect 56520 369578 56548 372807
rect 56968 372632 57020 372638
rect 56968 372574 57020 372580
rect 56508 369572 56560 369578
rect 56508 369514 56560 369520
rect 56876 351960 56928 351966
rect 56876 351902 56928 351908
rect 56690 303648 56746 303657
rect 56690 303583 56746 303592
rect 56704 198801 56732 303583
rect 56782 302288 56838 302297
rect 56782 302223 56838 302232
rect 56690 198792 56746 198801
rect 56690 198727 56746 198736
rect 56796 197441 56824 302223
rect 56888 266354 56916 351902
rect 56980 268977 57008 372574
rect 57150 305008 57206 305017
rect 57150 304943 57206 304952
rect 57058 300520 57114 300529
rect 57058 300455 57114 300464
rect 56966 268968 57022 268977
rect 56966 268903 57022 268912
rect 56876 266348 56928 266354
rect 56876 266290 56928 266296
rect 56980 258074 57008 268903
rect 56888 258046 57008 258074
rect 56782 197432 56838 197441
rect 56782 197367 56838 197376
rect 56508 165572 56560 165578
rect 56508 165514 56560 165520
rect 56520 164626 56548 165514
rect 56508 164620 56560 164626
rect 56508 164562 56560 164568
rect 56416 161968 56468 161974
rect 56416 161910 56468 161916
rect 55876 161446 56180 161474
rect 56046 145616 56102 145625
rect 56046 145551 56102 145560
rect 55956 144900 56008 144906
rect 55956 144842 56008 144848
rect 55864 144696 55916 144702
rect 55864 144638 55916 144644
rect 55876 58954 55904 144638
rect 55968 59362 55996 144842
rect 55956 59356 56008 59362
rect 55956 59298 56008 59304
rect 56060 59022 56088 145551
rect 56152 145314 56180 161446
rect 56888 161430 56916 258046
rect 56968 249008 57020 249014
rect 56968 248950 57020 248956
rect 56876 161424 56928 161430
rect 56876 161366 56928 161372
rect 56888 160177 56916 161366
rect 56874 160168 56930 160177
rect 56874 160103 56930 160112
rect 56322 146296 56378 146305
rect 56232 146260 56284 146266
rect 56322 146231 56378 146240
rect 56232 146202 56284 146208
rect 56140 145308 56192 145314
rect 56140 145250 56192 145256
rect 56048 59016 56100 59022
rect 56048 58958 56100 58964
rect 55864 58948 55916 58954
rect 55864 58890 55916 58896
rect 56152 56166 56180 145250
rect 56140 56160 56192 56166
rect 56140 56102 56192 56108
rect 55772 55208 55824 55214
rect 55772 55150 55824 55156
rect 55680 55072 55732 55078
rect 55680 55014 55732 55020
rect 56244 54806 56272 146202
rect 56336 145625 56364 146231
rect 56980 146130 57008 248950
rect 57072 195265 57100 300455
rect 57164 200977 57192 304943
rect 57256 278769 57284 382162
rect 57348 378706 57376 383438
rect 57532 383348 57560 459138
rect 57440 383320 57560 383348
rect 57440 378842 57468 383320
rect 57440 378814 57560 378842
rect 57348 378678 57468 378706
rect 57336 378616 57388 378622
rect 57336 378558 57388 378564
rect 57348 373794 57376 378558
rect 57336 373788 57388 373794
rect 57336 373730 57388 373736
rect 57440 306921 57468 378678
rect 57426 306912 57482 306921
rect 57426 306847 57482 306856
rect 57440 306374 57468 306847
rect 57348 306346 57468 306374
rect 57242 278760 57298 278769
rect 57242 278695 57298 278704
rect 57244 263560 57296 263566
rect 57244 263502 57296 263508
rect 57256 262313 57284 263502
rect 57242 262304 57298 262313
rect 57242 262239 57298 262248
rect 57348 201929 57376 306346
rect 57532 301345 57560 378814
rect 57624 302297 57652 463082
rect 57704 461712 57756 461718
rect 57704 461654 57756 461660
rect 57610 302288 57666 302297
rect 57610 302223 57666 302232
rect 57518 301336 57574 301345
rect 57440 301294 57518 301322
rect 57334 201920 57390 201929
rect 57334 201855 57390 201864
rect 57150 200968 57206 200977
rect 57150 200903 57206 200912
rect 57058 195256 57114 195265
rect 57058 195191 57114 195200
rect 57060 147552 57112 147558
rect 57058 147520 57060 147529
rect 57112 147520 57114 147529
rect 57058 147455 57114 147464
rect 56968 146124 57020 146130
rect 56968 146066 57020 146072
rect 56414 145888 56470 145897
rect 56414 145823 56470 145832
rect 56508 145852 56560 145858
rect 56322 145616 56378 145625
rect 56322 145551 56378 145560
rect 56428 144702 56456 145823
rect 56508 145794 56560 145800
rect 56520 144906 56548 145794
rect 57060 145648 57112 145654
rect 57060 145590 57112 145596
rect 56508 144900 56560 144906
rect 56508 144842 56560 144848
rect 57072 144770 57100 145590
rect 57060 144764 57112 144770
rect 57060 144706 57112 144712
rect 56416 144696 56468 144702
rect 56416 144638 56468 144644
rect 56876 69012 56928 69018
rect 56876 68954 56928 68960
rect 56888 68105 56916 68954
rect 56874 68096 56930 68105
rect 56874 68031 56930 68040
rect 57072 56234 57100 144706
rect 57164 96529 57192 200903
rect 57348 200114 57376 201855
rect 57256 200086 57376 200114
rect 57256 97481 57284 200086
rect 57334 197432 57390 197441
rect 57334 197367 57390 197376
rect 57242 97472 57298 97481
rect 57242 97407 57298 97416
rect 57150 96520 57206 96529
rect 57150 96455 57206 96464
rect 57348 93401 57376 197367
rect 57440 196081 57468 301294
rect 57518 301271 57574 301280
rect 57716 300529 57744 461654
rect 57808 303657 57836 467230
rect 57900 305969 57928 473962
rect 58624 472456 58676 472462
rect 58624 472398 58676 472404
rect 58532 469804 58584 469810
rect 58532 469746 58584 469752
rect 58440 469736 58492 469742
rect 58440 469678 58492 469684
rect 58452 411942 58480 469678
rect 58440 411936 58492 411942
rect 58440 411878 58492 411884
rect 58440 410848 58492 410854
rect 58440 410790 58492 410796
rect 58452 373522 58480 410790
rect 58440 373516 58492 373522
rect 58440 373458 58492 373464
rect 58544 372638 58572 469746
rect 58636 372745 58664 472398
rect 58716 465928 58768 465934
rect 58716 465870 58768 465876
rect 58622 372736 58678 372745
rect 58622 372671 58678 372680
rect 58532 372632 58584 372638
rect 58532 372574 58584 372580
rect 58624 353320 58676 353326
rect 58624 353262 58676 353268
rect 58532 350600 58584 350606
rect 58532 350542 58584 350548
rect 57886 305960 57942 305969
rect 57886 305895 57942 305904
rect 57900 305017 57928 305895
rect 57886 305008 57942 305017
rect 57886 304943 57942 304952
rect 57794 303648 57850 303657
rect 57794 303583 57850 303592
rect 57702 300520 57758 300529
rect 57702 300455 57758 300464
rect 57518 298208 57574 298217
rect 57518 298143 57574 298152
rect 57532 298110 57560 298143
rect 57520 298104 57572 298110
rect 57520 298046 57572 298052
rect 57426 196072 57482 196081
rect 57426 196007 57482 196016
rect 57426 195256 57482 195265
rect 57426 195191 57482 195200
rect 57334 93392 57390 93401
rect 57334 93327 57390 93336
rect 57440 90545 57468 195191
rect 57532 193225 57560 298046
rect 57886 278760 57942 278769
rect 57886 278695 57942 278704
rect 57796 264240 57848 264246
rect 57796 264182 57848 264188
rect 57808 263566 57836 264182
rect 57796 263560 57848 263566
rect 57796 263502 57848 263508
rect 57610 198792 57666 198801
rect 57610 198727 57666 198736
rect 57518 193216 57574 193225
rect 57518 193151 57574 193160
rect 57426 90536 57482 90545
rect 57426 90471 57482 90480
rect 57532 88233 57560 193151
rect 57624 93809 57652 198727
rect 57702 196072 57758 196081
rect 57702 196007 57758 196016
rect 57610 93800 57666 93809
rect 57610 93735 57666 93744
rect 57716 91089 57744 196007
rect 57796 173868 57848 173874
rect 57796 173810 57848 173816
rect 57808 173097 57836 173810
rect 57900 173369 57928 278695
rect 58544 268666 58572 350542
rect 58532 268660 58584 268666
rect 58532 268602 58584 268608
rect 58636 266354 58664 353262
rect 58728 279993 58756 465870
rect 58714 279984 58770 279993
rect 58714 279919 58770 279928
rect 58716 278724 58768 278730
rect 58716 278666 58768 278672
rect 58728 267918 58756 278666
rect 58820 278089 58848 475186
rect 58990 472832 59046 472841
rect 58990 472767 59046 472776
rect 58900 459332 58952 459338
rect 58900 459274 58952 459280
rect 58806 278080 58862 278089
rect 58806 278015 58862 278024
rect 58716 267912 58768 267918
rect 58716 267854 58768 267860
rect 57980 266348 58032 266354
rect 57980 266290 58032 266296
rect 58624 266348 58676 266354
rect 58624 266290 58676 266296
rect 57992 266218 58020 266290
rect 57980 266212 58032 266218
rect 57980 266154 58032 266160
rect 57980 266008 58032 266014
rect 57980 265950 58032 265956
rect 57992 264722 58020 265950
rect 57980 264716 58032 264722
rect 57980 264658 58032 264664
rect 57886 173360 57942 173369
rect 57886 173295 57942 173304
rect 57794 173088 57850 173097
rect 57794 173023 57850 173032
rect 57796 161016 57848 161022
rect 57796 160958 57848 160964
rect 57702 91080 57758 91089
rect 57702 91015 57758 91024
rect 57518 88224 57574 88233
rect 57518 88159 57574 88168
rect 57808 59226 57836 160958
rect 57900 68921 57928 173295
rect 57992 146266 58020 264658
rect 58716 250572 58768 250578
rect 58716 250514 58768 250520
rect 58624 250504 58676 250510
rect 58624 250446 58676 250452
rect 58636 249801 58664 250446
rect 58622 249792 58678 249801
rect 58728 249762 58756 250514
rect 58622 249727 58678 249736
rect 58716 249756 58768 249762
rect 58636 161362 58664 249727
rect 58716 249698 58768 249704
rect 58624 161356 58676 161362
rect 58624 161298 58676 161304
rect 58636 160138 58664 161298
rect 58728 160614 58756 249698
rect 58912 163606 58940 459274
rect 59004 175273 59032 472767
rect 59082 463312 59138 463321
rect 59082 463247 59138 463256
rect 58990 175264 59046 175273
rect 58990 175199 59046 175208
rect 59096 163674 59124 463247
rect 59188 164558 59216 478518
rect 59648 470594 59676 480066
rect 60568 476882 60596 480037
rect 60844 480023 61042 480051
rect 61120 480023 61502 480051
rect 60556 476876 60608 476882
rect 60556 476818 60608 476824
rect 59820 475856 59872 475862
rect 59820 475798 59872 475804
rect 59728 475176 59780 475182
rect 59728 475118 59780 475124
rect 59372 470566 59676 470594
rect 59372 467158 59400 470566
rect 59360 467152 59412 467158
rect 59360 467094 59412 467100
rect 59268 460148 59320 460154
rect 59268 460090 59320 460096
rect 59176 164552 59228 164558
rect 59176 164494 59228 164500
rect 59084 163668 59136 163674
rect 59084 163610 59136 163616
rect 58900 163600 58952 163606
rect 58900 163542 58952 163548
rect 59084 160948 59136 160954
rect 59084 160890 59136 160896
rect 58716 160608 58768 160614
rect 58716 160550 58768 160556
rect 58624 160132 58676 160138
rect 58624 160074 58676 160080
rect 57980 146260 58032 146266
rect 57980 146202 58032 146208
rect 58900 146260 58952 146266
rect 58900 146202 58952 146208
rect 57992 146062 58020 146202
rect 57980 146056 58032 146062
rect 57980 145998 58032 146004
rect 58622 146024 58678 146033
rect 58622 145959 58678 145968
rect 58636 144634 58664 145959
rect 58716 145920 58768 145926
rect 58716 145862 58768 145868
rect 58728 144838 58756 145862
rect 58716 144832 58768 144838
rect 58716 144774 58768 144780
rect 58624 144628 58676 144634
rect 58624 144570 58676 144576
rect 57886 68912 57942 68921
rect 57886 68847 57942 68856
rect 57796 59220 57848 59226
rect 57796 59162 57848 59168
rect 57900 57934 57928 68847
rect 57888 57928 57940 57934
rect 57888 57870 57940 57876
rect 57900 57594 57928 57870
rect 58072 57656 58124 57662
rect 58072 57598 58124 57604
rect 57244 57588 57296 57594
rect 57244 57530 57296 57536
rect 57888 57588 57940 57594
rect 57888 57530 57940 57536
rect 57060 56228 57112 56234
rect 57060 56170 57112 56176
rect 56232 54800 56284 54806
rect 56232 54742 56284 54748
rect 53380 54664 53432 54670
rect 53380 54606 53432 54612
rect 2780 20392 2832 20398
rect 2780 20334 2832 20340
rect 4804 20392 4856 20398
rect 4804 20334 4856 20340
rect 2792 19417 2820 20334
rect 2778 19408 2834 19417
rect 2778 19343 2834 19352
rect 57256 3466 57284 57530
rect 58084 57322 58112 57598
rect 58072 57316 58124 57322
rect 58072 57258 58124 57264
rect 58636 54874 58664 144570
rect 58728 56574 58756 144774
rect 58912 59090 58940 146202
rect 58992 146124 59044 146130
rect 58992 146066 59044 146072
rect 59004 145722 59032 146066
rect 58992 145716 59044 145722
rect 58992 145658 59044 145664
rect 58900 59084 58952 59090
rect 58900 59026 58952 59032
rect 58716 56568 58768 56574
rect 58716 56510 58768 56516
rect 58624 54868 58676 54874
rect 58624 54810 58676 54816
rect 59004 54738 59032 145658
rect 59096 59158 59124 160890
rect 59176 160132 59228 160138
rect 59176 160074 59228 160080
rect 59084 59152 59136 59158
rect 59084 59094 59136 59100
rect 59188 56370 59216 160074
rect 59280 57322 59308 460090
rect 59358 407824 59414 407833
rect 59358 407759 59414 407768
rect 59372 351966 59400 407759
rect 59450 373008 59506 373017
rect 59450 372943 59506 372952
rect 59464 352578 59492 372943
rect 59452 352572 59504 352578
rect 59452 352514 59504 352520
rect 59360 351960 59412 351966
rect 59360 351902 59412 351908
rect 59740 350606 59768 475118
rect 59728 350600 59780 350606
rect 59728 350542 59780 350548
rect 59832 269686 59860 475798
rect 60740 475380 60792 475386
rect 60740 475322 60792 475328
rect 60002 463176 60058 463185
rect 60002 463111 60058 463120
rect 59912 460080 59964 460086
rect 59912 460022 59964 460028
rect 59820 269680 59872 269686
rect 59820 269622 59872 269628
rect 59820 267912 59872 267918
rect 59820 267854 59872 267860
rect 59728 265668 59780 265674
rect 59728 265610 59780 265616
rect 59740 264858 59768 265610
rect 59728 264852 59780 264858
rect 59728 264794 59780 264800
rect 59360 160744 59412 160750
rect 59360 160686 59412 160692
rect 59372 140865 59400 160686
rect 59740 147626 59768 264794
rect 59728 147620 59780 147626
rect 59728 147562 59780 147568
rect 59740 146146 59768 147562
rect 59832 146266 59860 267854
rect 59924 163810 59952 460022
rect 59912 163804 59964 163810
rect 59912 163746 59964 163752
rect 60016 163538 60044 463111
rect 60752 460698 60780 475322
rect 60844 468518 60872 480023
rect 61120 475386 61148 480023
rect 61108 475380 61160 475386
rect 61108 475322 61160 475328
rect 61948 471306 61976 480037
rect 62224 480023 62330 480051
rect 62120 475380 62172 475386
rect 62120 475322 62172 475328
rect 61936 471300 61988 471306
rect 61936 471242 61988 471248
rect 60832 468512 60884 468518
rect 60832 468454 60884 468460
rect 60740 460692 60792 460698
rect 60740 460634 60792 460640
rect 62132 460630 62160 475322
rect 62224 469062 62252 480023
rect 62776 478242 62804 480037
rect 62960 480023 63250 480051
rect 62764 478236 62816 478242
rect 62764 478178 62816 478184
rect 62960 475386 62988 480023
rect 63696 478854 63724 480037
rect 63684 478848 63736 478854
rect 63684 478790 63736 478796
rect 64156 478106 64184 480037
rect 64248 480023 64538 480051
rect 64892 480023 64998 480051
rect 65076 480023 65458 480051
rect 65536 480023 65918 480051
rect 64144 478100 64196 478106
rect 64144 478042 64196 478048
rect 62948 475380 63000 475386
rect 62948 475322 63000 475328
rect 63040 475380 63092 475386
rect 63040 475322 63092 475328
rect 63052 475114 63080 475322
rect 63040 475108 63092 475114
rect 63040 475050 63092 475056
rect 64248 470594 64276 480023
rect 63696 470566 64276 470594
rect 62212 469056 62264 469062
rect 62212 468998 62264 469004
rect 63696 462806 63724 470566
rect 64892 462874 64920 480023
rect 65076 475402 65104 480023
rect 64984 475374 65104 475402
rect 64984 465526 65012 475374
rect 65536 470594 65564 480023
rect 66258 478272 66314 478281
rect 66258 478207 66314 478216
rect 66272 477873 66300 478207
rect 66258 477864 66314 477873
rect 66258 477799 66314 477808
rect 66364 475969 66392 480037
rect 66456 480023 66746 480051
rect 66824 480023 67206 480051
rect 66350 475960 66406 475969
rect 66350 475895 66406 475904
rect 66260 475108 66312 475114
rect 66260 475050 66312 475056
rect 65076 470566 65564 470594
rect 65076 465594 65104 470566
rect 65064 465588 65116 465594
rect 65064 465530 65116 465536
rect 64972 465520 65024 465526
rect 64972 465462 65024 465468
rect 64880 462868 64932 462874
rect 64880 462810 64932 462816
rect 63684 462800 63736 462806
rect 63684 462742 63736 462748
rect 62120 460624 62172 460630
rect 62120 460566 62172 460572
rect 66272 460494 66300 475050
rect 66456 470594 66484 480023
rect 66824 475114 66852 480023
rect 67652 475402 67680 480037
rect 67560 475374 67680 475402
rect 67928 480023 68126 480051
rect 68204 480023 68494 480051
rect 68664 480023 68954 480051
rect 69032 480023 69414 480051
rect 69492 480023 69874 480051
rect 69952 480023 70334 480051
rect 70504 480023 70702 480051
rect 70872 480023 71162 480051
rect 71240 480023 71622 480051
rect 67560 475130 67588 475374
rect 66812 475108 66864 475114
rect 67560 475102 67772 475130
rect 66812 475050 66864 475056
rect 67640 475040 67692 475046
rect 67640 474982 67692 474988
rect 66364 470566 66484 470594
rect 66364 460766 66392 470566
rect 66352 460760 66404 460766
rect 66352 460702 66404 460708
rect 66260 460488 66312 460494
rect 66260 460430 66312 460436
rect 67652 459105 67680 474982
rect 67744 460154 67772 475102
rect 67824 475108 67876 475114
rect 67824 475050 67876 475056
rect 67836 460737 67864 475050
rect 67928 475046 67956 480023
rect 67916 475040 67968 475046
rect 67916 474982 67968 474988
rect 68204 470594 68232 480023
rect 68284 478848 68336 478854
rect 68284 478790 68336 478796
rect 67928 470566 68232 470594
rect 67928 461689 67956 470566
rect 67914 461680 67970 461689
rect 67914 461615 67970 461624
rect 67822 460728 67878 460737
rect 67822 460663 67878 460672
rect 67732 460148 67784 460154
rect 67732 460090 67784 460096
rect 68296 460086 68324 478790
rect 68664 475114 68692 480023
rect 68652 475108 68704 475114
rect 68652 475050 68704 475056
rect 68284 460080 68336 460086
rect 68284 460022 68336 460028
rect 67638 459096 67694 459105
rect 67638 459031 67694 459040
rect 69032 458833 69060 480023
rect 69492 475402 69520 480023
rect 69124 475374 69520 475402
rect 69124 458969 69152 475374
rect 69952 470594 69980 480023
rect 70400 476128 70452 476134
rect 70400 476070 70452 476076
rect 69216 470566 69980 470594
rect 69216 460873 69244 470566
rect 69202 460864 69258 460873
rect 69202 460799 69258 460808
rect 70412 460562 70440 476070
rect 70504 463457 70532 480023
rect 70872 476134 70900 480023
rect 70860 476128 70912 476134
rect 70860 476070 70912 476076
rect 71240 475402 71268 480023
rect 72068 478825 72096 480037
rect 72054 478816 72110 478825
rect 72054 478751 72110 478760
rect 72424 478100 72476 478106
rect 72424 478042 72476 478048
rect 71320 477896 71372 477902
rect 71320 477838 71372 477844
rect 70596 475374 71268 475402
rect 70596 466313 70624 475374
rect 71332 470594 71360 477838
rect 71780 475108 71832 475114
rect 71780 475050 71832 475056
rect 71056 470566 71360 470594
rect 70582 466304 70638 466313
rect 70582 466239 70638 466248
rect 70490 463448 70546 463457
rect 70490 463383 70546 463392
rect 71056 461650 71084 470566
rect 71044 461644 71096 461650
rect 71044 461586 71096 461592
rect 70400 460556 70452 460562
rect 70400 460498 70452 460504
rect 71792 460222 71820 475050
rect 72436 460222 72464 478042
rect 72528 478009 72556 480037
rect 72620 480023 72910 480051
rect 73264 480023 73370 480051
rect 73448 480023 73830 480051
rect 72514 478000 72570 478009
rect 72514 477935 72570 477944
rect 72620 475114 72648 480023
rect 73158 478816 73214 478825
rect 73158 478751 73160 478760
rect 73212 478751 73214 478760
rect 73160 478722 73212 478728
rect 73158 478680 73214 478689
rect 73158 478615 73214 478624
rect 73172 478378 73200 478615
rect 73160 478372 73212 478378
rect 73160 478314 73212 478320
rect 72608 475108 72660 475114
rect 72608 475050 72660 475056
rect 73264 461553 73292 480023
rect 73448 478961 73476 480023
rect 73434 478952 73490 478961
rect 73434 478887 73490 478896
rect 74276 478514 74304 480037
rect 74264 478508 74316 478514
rect 74264 478450 74316 478456
rect 74356 478508 74408 478514
rect 74356 478450 74408 478456
rect 73896 478372 73948 478378
rect 73896 478314 73948 478320
rect 73804 477556 73856 477562
rect 73804 477498 73856 477504
rect 73250 461544 73306 461553
rect 73250 461479 73306 461488
rect 73816 460426 73844 477498
rect 73908 468994 73936 478314
rect 74080 478100 74132 478106
rect 74080 478042 74132 478048
rect 73988 477964 74040 477970
rect 73988 477906 74040 477912
rect 73896 468988 73948 468994
rect 73896 468930 73948 468936
rect 74000 468926 74028 477906
rect 73988 468920 74040 468926
rect 73988 468862 74040 468868
rect 74092 468858 74120 478042
rect 74172 478032 74224 478038
rect 74172 477974 74224 477980
rect 74080 468852 74132 468858
rect 74080 468794 74132 468800
rect 74184 468790 74212 477974
rect 74368 477562 74396 478450
rect 74644 478417 74672 480037
rect 74736 480023 75118 480051
rect 75288 480023 75578 480051
rect 74630 478408 74686 478417
rect 74630 478343 74686 478352
rect 74356 477556 74408 477562
rect 74356 477498 74408 477504
rect 74540 475108 74592 475114
rect 74540 475050 74592 475056
rect 74172 468784 74224 468790
rect 74172 468726 74224 468732
rect 73804 460420 73856 460426
rect 73804 460362 73856 460368
rect 71780 460216 71832 460222
rect 71780 460158 71832 460164
rect 72424 460216 72476 460222
rect 72424 460158 72476 460164
rect 74552 460057 74580 475050
rect 74736 470594 74764 480023
rect 75288 475114 75316 480023
rect 76024 478281 76052 480037
rect 76010 478272 76066 478281
rect 76010 478207 76066 478216
rect 76484 477873 76512 480037
rect 76576 480023 76866 480051
rect 76470 477864 76526 477873
rect 76470 477799 76526 477808
rect 75276 475108 75328 475114
rect 75276 475050 75328 475056
rect 76576 470594 76604 480023
rect 77312 478650 77340 480037
rect 77772 478689 77800 480037
rect 77864 480023 78246 480051
rect 77758 478680 77814 478689
rect 77300 478644 77352 478650
rect 77758 478615 77814 478624
rect 77300 478586 77352 478592
rect 77864 470594 77892 480023
rect 74644 470566 74764 470594
rect 75932 470566 76604 470594
rect 77404 470566 77892 470594
rect 74644 460465 74672 470566
rect 74630 460456 74686 460465
rect 74630 460391 74686 460400
rect 75932 460329 75960 470566
rect 77404 460601 77432 470566
rect 77390 460592 77446 460601
rect 77390 460527 77446 460536
rect 75918 460320 75974 460329
rect 75918 460255 75974 460264
rect 78692 460193 78720 480037
rect 78876 480023 79074 480051
rect 78772 475108 78824 475114
rect 78772 475050 78824 475056
rect 78784 460834 78812 475050
rect 78772 460828 78824 460834
rect 78772 460770 78824 460776
rect 78876 460358 78904 480023
rect 79520 478825 79548 480037
rect 79704 480023 79994 480051
rect 80072 480023 80454 480051
rect 79506 478816 79562 478825
rect 79506 478751 79562 478760
rect 79704 475114 79732 480023
rect 79692 475108 79744 475114
rect 79692 475050 79744 475056
rect 80072 460902 80100 480023
rect 80808 478145 80836 480037
rect 80794 478136 80850 478145
rect 80794 478071 80850 478080
rect 81268 472977 81296 480037
rect 81728 478718 81756 480037
rect 81912 480023 82202 480051
rect 82280 480023 82662 480051
rect 82832 480023 83030 480051
rect 83108 480023 83490 480051
rect 83568 480023 83950 480051
rect 81716 478712 81768 478718
rect 81716 478654 81768 478660
rect 81254 472968 81310 472977
rect 81254 472903 81310 472912
rect 81532 471232 81584 471238
rect 81532 471174 81584 471180
rect 81544 465905 81572 471174
rect 81912 466454 81940 480023
rect 82280 471238 82308 480023
rect 82832 471238 82860 480023
rect 83108 476114 83136 480023
rect 82924 476086 83136 476114
rect 82268 471232 82320 471238
rect 82268 471174 82320 471180
rect 82820 471232 82872 471238
rect 82820 471174 82872 471180
rect 82820 471096 82872 471102
rect 82820 471038 82872 471044
rect 81636 466426 81940 466454
rect 81530 465896 81586 465905
rect 81530 465831 81586 465840
rect 81636 463622 81664 466426
rect 82832 465662 82860 471038
rect 82924 466342 82952 476086
rect 83004 471232 83056 471238
rect 83004 471174 83056 471180
rect 83016 466410 83044 471174
rect 83568 471102 83596 480023
rect 84396 478990 84424 480037
rect 84384 478984 84436 478990
rect 84384 478926 84436 478932
rect 84856 477902 84884 480037
rect 84948 480023 85238 480051
rect 84844 477896 84896 477902
rect 84844 477838 84896 477844
rect 83556 471096 83608 471102
rect 83556 471038 83608 471044
rect 84948 466454 84976 480023
rect 85580 476128 85632 476134
rect 85580 476070 85632 476076
rect 84304 466426 84976 466454
rect 83004 466404 83056 466410
rect 83004 466346 83056 466352
rect 82912 466336 82964 466342
rect 82912 466278 82964 466284
rect 84304 466041 84332 466426
rect 84290 466032 84346 466041
rect 84290 465967 84346 465976
rect 82820 465656 82872 465662
rect 82820 465598 82872 465604
rect 81624 463616 81676 463622
rect 81624 463558 81676 463564
rect 85592 462942 85620 476070
rect 85684 471322 85712 480037
rect 85776 480023 86158 480051
rect 86328 480023 86618 480051
rect 86972 480023 87078 480051
rect 87156 480023 87446 480051
rect 87524 480023 87906 480051
rect 88366 480023 88656 480051
rect 85776 476134 85804 480023
rect 85764 476128 85816 476134
rect 85764 476070 85816 476076
rect 85684 471294 85804 471322
rect 85672 471232 85724 471238
rect 85672 471174 85724 471180
rect 85684 463418 85712 471174
rect 85776 466177 85804 471294
rect 86328 471238 86356 480023
rect 86316 471232 86368 471238
rect 86316 471174 86368 471180
rect 85762 466168 85818 466177
rect 85762 466103 85818 466112
rect 86972 463690 87000 480023
rect 87156 476114 87184 480023
rect 87064 476086 87184 476114
rect 86960 463684 87012 463690
rect 86960 463626 87012 463632
rect 85672 463412 85724 463418
rect 85672 463354 85724 463360
rect 87064 463078 87092 476086
rect 87524 466454 87552 480023
rect 88524 468172 88576 468178
rect 88524 468114 88576 468120
rect 88432 468036 88484 468042
rect 88432 467978 88484 467984
rect 87156 466426 87552 466454
rect 87156 463486 87184 466426
rect 87144 463480 87196 463486
rect 87144 463422 87196 463428
rect 88444 463282 88472 467978
rect 88536 463350 88564 468114
rect 88628 463554 88656 480023
rect 88720 480023 88826 480051
rect 88720 468042 88748 480023
rect 89180 478446 89208 480037
rect 89272 480023 89654 480051
rect 89824 480023 90114 480051
rect 90192 480023 90574 480051
rect 89168 478440 89220 478446
rect 89168 478382 89220 478388
rect 89272 468178 89300 480023
rect 89260 468172 89312 468178
rect 89260 468114 89312 468120
rect 88708 468036 88760 468042
rect 88708 467978 88760 467984
rect 88616 463548 88668 463554
rect 88616 463490 88668 463496
rect 88524 463344 88576 463350
rect 88524 463286 88576 463292
rect 88432 463276 88484 463282
rect 88432 463218 88484 463224
rect 89824 463214 89852 480023
rect 90192 470594 90220 480023
rect 91020 478582 91048 480037
rect 91008 478576 91060 478582
rect 91008 478518 91060 478524
rect 91388 477970 91416 480037
rect 91848 478854 91876 480037
rect 91940 480023 92322 480051
rect 92492 480023 92782 480051
rect 92860 480023 93242 480051
rect 93320 480023 93610 480051
rect 93964 480023 94070 480051
rect 94240 480023 94530 480051
rect 91836 478848 91888 478854
rect 91836 478790 91888 478796
rect 91376 477964 91428 477970
rect 91376 477906 91428 477912
rect 91940 470594 91968 480023
rect 89916 470566 90220 470594
rect 91204 470566 91968 470594
rect 89812 463208 89864 463214
rect 89812 463150 89864 463156
rect 87052 463072 87104 463078
rect 87052 463014 87104 463020
rect 85580 462936 85632 462942
rect 85580 462878 85632 462884
rect 80060 460896 80112 460902
rect 80060 460838 80112 460844
rect 78864 460352 78916 460358
rect 78864 460294 78916 460300
rect 78678 460184 78734 460193
rect 78678 460119 78734 460128
rect 74538 460048 74594 460057
rect 74538 459983 74594 459992
rect 89916 459270 89944 470566
rect 91204 463321 91232 470566
rect 91190 463312 91246 463321
rect 91190 463247 91246 463256
rect 92492 459338 92520 480023
rect 92572 475108 92624 475114
rect 92572 475050 92624 475056
rect 92584 460290 92612 475050
rect 92860 470594 92888 480023
rect 93320 475114 93348 480023
rect 93308 475108 93360 475114
rect 93308 475050 93360 475056
rect 92676 470566 92888 470594
rect 92676 463185 92704 470566
rect 92662 463176 92718 463185
rect 92662 463111 92718 463120
rect 93964 463049 93992 480023
rect 94240 470594 94268 480023
rect 94976 478038 95004 480037
rect 95344 478106 95372 480037
rect 95332 478100 95384 478106
rect 95332 478042 95384 478048
rect 94964 478032 95016 478038
rect 94964 477974 95016 477980
rect 95804 472841 95832 480037
rect 96264 475250 96292 480037
rect 96724 475318 96752 480037
rect 97184 475998 97212 480037
rect 97172 475992 97224 475998
rect 97172 475934 97224 475940
rect 96712 475312 96764 475318
rect 96712 475254 96764 475260
rect 96252 475244 96304 475250
rect 96252 475186 96304 475192
rect 97552 475182 97580 480037
rect 98012 475930 98040 480037
rect 98472 476066 98500 480037
rect 98564 480023 98946 480051
rect 98460 476060 98512 476066
rect 98460 476002 98512 476008
rect 98000 475924 98052 475930
rect 98000 475866 98052 475872
rect 97540 475176 97592 475182
rect 97540 475118 97592 475124
rect 95790 472832 95846 472841
rect 95790 472767 95846 472776
rect 98564 470594 98592 480023
rect 99392 478922 99420 480037
rect 99484 480023 99774 480051
rect 99380 478916 99432 478922
rect 99380 478858 99432 478864
rect 94056 470566 94268 470594
rect 98196 470566 98592 470594
rect 93950 463040 94006 463049
rect 93950 462975 94006 462984
rect 94056 462913 94084 470566
rect 98196 466002 98224 470566
rect 99484 466206 99512 480023
rect 100220 478310 100248 480037
rect 100312 480023 100694 480051
rect 100772 480023 101154 480051
rect 101232 480023 101522 480051
rect 101600 480023 101982 480051
rect 100208 478304 100260 478310
rect 100208 478246 100260 478252
rect 100312 470594 100340 480023
rect 99576 470566 100340 470594
rect 99472 466200 99524 466206
rect 99472 466142 99524 466148
rect 98184 465996 98236 466002
rect 98184 465938 98236 465944
rect 94042 462904 94098 462913
rect 94042 462839 94098 462848
rect 92572 460284 92624 460290
rect 92572 460226 92624 460232
rect 92480 459332 92532 459338
rect 92480 459274 92532 459280
rect 89904 459264 89956 459270
rect 89904 459206 89956 459212
rect 69110 458960 69166 458969
rect 69110 458895 69166 458904
rect 99576 458862 99604 470566
rect 100772 463010 100800 480023
rect 100852 475312 100904 475318
rect 100852 475254 100904 475260
rect 100864 466070 100892 475254
rect 101232 470594 101260 480023
rect 101600 475318 101628 480023
rect 102428 478174 102456 480037
rect 102520 480023 102902 480051
rect 102980 480023 103362 480051
rect 102416 478168 102468 478174
rect 102416 478110 102468 478116
rect 102520 475402 102548 480023
rect 102244 475374 102548 475402
rect 101588 475312 101640 475318
rect 101588 475254 101640 475260
rect 100956 470566 101260 470594
rect 100956 466138 100984 470566
rect 100944 466132 100996 466138
rect 100944 466074 100996 466080
rect 100852 466064 100904 466070
rect 100852 466006 100904 466012
rect 102244 465769 102272 475374
rect 102980 470594 103008 480023
rect 103612 475312 103664 475318
rect 103612 475254 103664 475260
rect 103520 475244 103572 475250
rect 103520 475186 103572 475192
rect 102336 470566 103008 470594
rect 102230 465760 102286 465769
rect 102230 465695 102286 465704
rect 102336 464370 102364 470566
rect 103532 465730 103560 475186
rect 103624 466274 103652 475254
rect 103716 468722 103744 480037
rect 103808 480023 104190 480051
rect 104360 480023 104650 480051
rect 103808 475318 103836 480023
rect 103796 475312 103848 475318
rect 103796 475254 103848 475260
rect 104360 475250 104388 480023
rect 105096 478514 105124 480037
rect 105188 480023 105570 480051
rect 105648 480023 105938 480051
rect 106398 480023 106504 480051
rect 105084 478508 105136 478514
rect 105084 478450 105136 478456
rect 104992 475312 105044 475318
rect 104992 475254 105044 475260
rect 104348 475244 104400 475250
rect 104348 475186 104400 475192
rect 103704 468716 103756 468722
rect 103704 468658 103756 468664
rect 103612 466268 103664 466274
rect 103612 466210 103664 466216
rect 105004 465798 105032 475254
rect 105188 470594 105216 480023
rect 105648 475318 105676 480023
rect 105636 475312 105688 475318
rect 105636 475254 105688 475260
rect 106372 475312 106424 475318
rect 106372 475254 106424 475260
rect 106280 475244 106332 475250
rect 106280 475186 106332 475192
rect 105096 470566 105216 470594
rect 105096 465866 105124 470566
rect 106292 467226 106320 475186
rect 106384 468586 106412 475254
rect 106476 468654 106504 480023
rect 106568 480023 106858 480051
rect 106936 480023 107318 480051
rect 106568 475318 106596 480023
rect 106556 475312 106608 475318
rect 106556 475254 106608 475260
rect 106936 475250 106964 480023
rect 107764 478961 107792 480037
rect 107856 480023 108146 480051
rect 108224 480023 108606 480051
rect 109066 480023 109172 480051
rect 107750 478952 107806 478961
rect 107750 478887 107806 478896
rect 107856 475300 107884 480023
rect 107672 475272 107884 475300
rect 106924 475244 106976 475250
rect 106924 475186 106976 475192
rect 106464 468648 106516 468654
rect 106464 468590 106516 468596
rect 106372 468580 106424 468586
rect 106372 468522 106424 468528
rect 106280 467220 106332 467226
rect 106280 467162 106332 467168
rect 105084 465860 105136 465866
rect 105084 465802 105136 465808
rect 104992 465792 105044 465798
rect 104992 465734 105044 465740
rect 103520 465724 103572 465730
rect 103520 465666 103572 465672
rect 102324 464364 102376 464370
rect 102324 464306 102376 464312
rect 100760 463004 100812 463010
rect 100760 462946 100812 462952
rect 107672 461650 107700 475272
rect 108224 470594 108252 480023
rect 107764 470566 108252 470594
rect 107764 463078 107792 470566
rect 107752 463072 107804 463078
rect 107752 463014 107804 463020
rect 109144 463010 109172 480023
rect 109512 478922 109540 480037
rect 109604 480023 109894 480051
rect 109500 478916 109552 478922
rect 109500 478858 109552 478864
rect 109604 470594 109632 480023
rect 110340 478378 110368 480037
rect 110616 480023 110814 480051
rect 110328 478372 110380 478378
rect 110328 478314 110380 478320
rect 109328 470566 109632 470594
rect 109132 463004 109184 463010
rect 109132 462946 109184 462952
rect 107660 461644 107712 461650
rect 107660 461586 107712 461592
rect 109328 458862 109356 470566
rect 110616 465934 110644 480023
rect 111260 475658 111288 480037
rect 111720 475794 111748 480037
rect 111708 475788 111760 475794
rect 111708 475730 111760 475736
rect 112088 475726 112116 480037
rect 112180 480023 112562 480051
rect 112640 480023 113022 480051
rect 112076 475720 112128 475726
rect 112076 475662 112128 475668
rect 111248 475652 111300 475658
rect 111248 475594 111300 475600
rect 112180 475300 112208 480023
rect 111904 475272 112208 475300
rect 110604 465928 110656 465934
rect 110604 465870 110656 465876
rect 111904 461718 111932 475272
rect 112640 470594 112668 480023
rect 113272 475312 113324 475318
rect 113272 475254 113324 475260
rect 111996 470566 112668 470594
rect 111892 461712 111944 461718
rect 111892 461654 111944 461660
rect 111996 459202 112024 470566
rect 113284 467294 113312 475254
rect 113468 470642 113496 480037
rect 113560 480023 113942 480051
rect 113560 475318 113588 480023
rect 113548 475312 113600 475318
rect 113548 475254 113600 475260
rect 114296 474026 114324 480037
rect 114284 474020 114336 474026
rect 114284 473962 114336 473968
rect 113376 470614 113496 470642
rect 113272 467288 113324 467294
rect 113272 467230 113324 467236
rect 113376 463146 113404 470614
rect 114756 464438 114784 480037
rect 115216 475590 115244 480037
rect 115204 475584 115256 475590
rect 115204 475526 115256 475532
rect 115676 475522 115704 480037
rect 115664 475516 115716 475522
rect 115664 475458 115716 475464
rect 116044 472530 116072 480037
rect 116308 478236 116360 478242
rect 116308 478178 116360 478184
rect 116320 474065 116348 478178
rect 116306 474056 116362 474065
rect 116306 473991 116362 474000
rect 116504 473278 116532 480037
rect 116492 473272 116544 473278
rect 116492 473214 116544 473220
rect 116964 472598 116992 480037
rect 117438 480023 117544 480051
rect 116952 472592 117004 472598
rect 116952 472534 117004 472540
rect 116032 472524 116084 472530
rect 116032 472466 116084 472472
rect 114744 464432 114796 464438
rect 114744 464374 114796 464380
rect 113364 463140 113416 463146
rect 113364 463082 113416 463088
rect 111984 459196 112036 459202
rect 111984 459138 112036 459144
rect 117516 459134 117544 480023
rect 117884 473346 117912 480037
rect 117872 473340 117924 473346
rect 117872 473282 117924 473288
rect 118252 473142 118280 480037
rect 118240 473136 118292 473142
rect 118240 473078 118292 473084
rect 118712 472462 118740 480037
rect 119172 473210 119200 480037
rect 119632 475862 119660 480037
rect 119620 475856 119672 475862
rect 119620 475798 119672 475804
rect 120092 475454 120120 480037
rect 120460 475561 120488 480037
rect 120920 475697 120948 480037
rect 121380 475833 121408 480037
rect 121366 475824 121422 475833
rect 121366 475759 121422 475768
rect 120906 475688 120962 475697
rect 120906 475623 120962 475632
rect 120446 475552 120502 475561
rect 120446 475487 120502 475496
rect 120080 475448 120132 475454
rect 120080 475390 120132 475396
rect 119160 473204 119212 473210
rect 119160 473146 119212 473152
rect 121840 472569 121868 480037
rect 121932 480023 122222 480051
rect 121826 472560 121882 472569
rect 121826 472495 121882 472504
rect 118700 472456 118752 472462
rect 118700 472398 118752 472404
rect 121932 470594 121960 480023
rect 122668 472705 122696 480037
rect 123036 480023 123142 480051
rect 123312 480023 123602 480051
rect 123680 480023 124062 480051
rect 124324 480023 124430 480051
rect 124508 480023 124890 480051
rect 124968 480023 125350 480051
rect 125704 480023 125810 480051
rect 125888 480023 126270 480051
rect 126348 480023 126638 480051
rect 126992 480023 127098 480051
rect 127176 480023 127558 480051
rect 127728 480023 128018 480051
rect 128372 480023 128478 480051
rect 128556 480023 128846 480051
rect 122840 475448 122892 475454
rect 122840 475390 122892 475396
rect 122654 472696 122710 472705
rect 122654 472631 122710 472640
rect 121472 470566 121960 470594
rect 117504 459128 117556 459134
rect 117504 459070 117556 459076
rect 121472 459066 121500 470566
rect 122852 470354 122880 475390
rect 122932 475312 122984 475318
rect 122932 475254 122984 475260
rect 122840 470348 122892 470354
rect 122840 470290 122892 470296
rect 122944 470286 122972 475254
rect 122932 470280 122984 470286
rect 122932 470222 122984 470228
rect 123036 470150 123064 480023
rect 123312 475318 123340 480023
rect 123680 475454 123708 480023
rect 123668 475448 123720 475454
rect 123668 475390 123720 475396
rect 123300 475312 123352 475318
rect 123300 475254 123352 475260
rect 124220 475312 124272 475318
rect 124220 475254 124272 475260
rect 123024 470144 123076 470150
rect 123024 470086 123076 470092
rect 124232 465769 124260 475254
rect 124324 469985 124352 480023
rect 124508 470594 124536 480023
rect 124968 475318 124996 480023
rect 124956 475312 125008 475318
rect 124956 475254 125008 475260
rect 125600 475312 125652 475318
rect 125600 475254 125652 475260
rect 124416 470566 124536 470594
rect 124416 470218 124444 470566
rect 124404 470212 124456 470218
rect 124404 470154 124456 470160
rect 124310 469976 124366 469985
rect 124310 469911 124366 469920
rect 124218 465760 124274 465769
rect 124218 465695 124274 465704
rect 125612 459066 125640 475254
rect 121460 459060 121512 459066
rect 121460 459002 121512 459008
rect 125600 459060 125652 459066
rect 125600 459002 125652 459008
rect 99564 458856 99616 458862
rect 69018 458824 69074 458833
rect 99564 458798 99616 458804
rect 109316 458856 109368 458862
rect 125704 458833 125732 480023
rect 125888 470594 125916 480023
rect 126348 475318 126376 480023
rect 126336 475312 126388 475318
rect 126336 475254 126388 475260
rect 125796 470566 125916 470594
rect 125796 465730 125824 470566
rect 126992 469742 127020 480023
rect 127176 475300 127204 480023
rect 127084 475272 127204 475300
rect 127084 470490 127112 475272
rect 127728 470594 127756 480023
rect 127176 470566 127756 470594
rect 127072 470484 127124 470490
rect 127072 470426 127124 470432
rect 127176 469810 127204 470566
rect 128372 470558 128400 480023
rect 128360 470552 128412 470558
rect 128360 470494 128412 470500
rect 128556 469849 128584 480023
rect 129292 471374 129320 480037
rect 129752 472870 129780 480037
rect 130028 480023 130226 480051
rect 129740 472864 129792 472870
rect 129740 472806 129792 472812
rect 129280 471368 129332 471374
rect 129280 471310 129332 471316
rect 128542 469840 128598 469849
rect 127164 469804 127216 469810
rect 128542 469775 128598 469784
rect 127164 469746 127216 469752
rect 126980 469736 127032 469742
rect 126980 469678 127032 469684
rect 125784 465724 125836 465730
rect 125784 465666 125836 465672
rect 130028 458998 130056 480023
rect 130580 472734 130608 480037
rect 131040 472802 131068 480037
rect 131500 472938 131528 480037
rect 131960 473074 131988 480037
rect 132144 480023 132434 480051
rect 131948 473068 132000 473074
rect 131948 473010 132000 473016
rect 131488 472932 131540 472938
rect 131488 472874 131540 472880
rect 131028 472796 131080 472802
rect 131028 472738 131080 472744
rect 130568 472728 130620 472734
rect 130568 472670 130620 472676
rect 132144 469878 132172 480023
rect 132788 470422 132816 480037
rect 132880 480023 133262 480051
rect 133432 480023 133722 480051
rect 133984 480023 134182 480051
rect 134352 480023 134642 480051
rect 132776 470416 132828 470422
rect 132776 470358 132828 470364
rect 132880 469946 132908 480023
rect 133144 476876 133196 476882
rect 133144 476818 133196 476824
rect 132868 469940 132920 469946
rect 132868 469882 132920 469888
rect 132132 469872 132184 469878
rect 132132 469814 132184 469820
rect 133156 462330 133184 476818
rect 133432 470014 133460 480023
rect 133984 470082 134012 480023
rect 133972 470076 134024 470082
rect 133972 470018 134024 470024
rect 133420 470008 133472 470014
rect 133420 469950 133472 469956
rect 134352 466454 134380 480023
rect 134996 475386 135024 480037
rect 134984 475380 135036 475386
rect 134984 475322 135036 475328
rect 135456 475250 135484 480037
rect 135916 475522 135944 480037
rect 135904 475516 135956 475522
rect 135904 475458 135956 475464
rect 135444 475244 135496 475250
rect 135444 475186 135496 475192
rect 136376 473006 136404 480037
rect 136744 475454 136772 480037
rect 136928 480023 137218 480051
rect 136732 475448 136784 475454
rect 136732 475390 136784 475396
rect 136364 473000 136416 473006
rect 136364 472942 136416 472948
rect 136928 466454 136956 480023
rect 137664 475726 137692 480037
rect 137652 475720 137704 475726
rect 137652 475662 137704 475668
rect 138124 475590 138152 480037
rect 138584 475658 138612 480037
rect 138952 478174 138980 480037
rect 138940 478168 138992 478174
rect 138940 478110 138992 478116
rect 139412 478038 139440 480037
rect 139504 480023 139886 480051
rect 140056 480023 140346 480051
rect 139400 478032 139452 478038
rect 139400 477974 139452 477980
rect 138572 475652 138624 475658
rect 138572 475594 138624 475600
rect 138112 475584 138164 475590
rect 138112 475526 138164 475532
rect 139400 475380 139452 475386
rect 139400 475322 139452 475328
rect 134076 466426 134380 466454
rect 136652 466426 136956 466454
rect 133144 462324 133196 462330
rect 133144 462266 133196 462272
rect 130016 458992 130068 458998
rect 130016 458934 130068 458940
rect 134076 458930 134104 466426
rect 136652 458998 136680 466426
rect 139412 466002 139440 475322
rect 139504 468586 139532 480023
rect 140056 475386 140084 480023
rect 140792 478990 140820 480037
rect 140976 480023 141174 480051
rect 141344 480023 141634 480051
rect 141712 480023 142094 480051
rect 142264 480023 142554 480051
rect 142632 480023 142922 480051
rect 143000 480023 143382 480051
rect 140780 478984 140832 478990
rect 140780 478926 140832 478932
rect 140044 475380 140096 475386
rect 140044 475322 140096 475328
rect 140872 475380 140924 475386
rect 140872 475322 140924 475328
rect 140780 475312 140832 475318
rect 140780 475254 140832 475260
rect 139492 468580 139544 468586
rect 139492 468522 139544 468528
rect 139400 465996 139452 466002
rect 139400 465938 139452 465944
rect 140792 465866 140820 475254
rect 140780 465860 140832 465866
rect 140780 465802 140832 465808
rect 140884 465798 140912 475322
rect 140976 465934 141004 480023
rect 141344 475318 141372 480023
rect 141712 475386 141740 480023
rect 141700 475380 141752 475386
rect 141700 475322 141752 475328
rect 141332 475312 141384 475318
rect 141332 475254 141384 475260
rect 142160 475176 142212 475182
rect 142160 475118 142212 475124
rect 140964 465928 141016 465934
rect 140964 465870 141016 465876
rect 140872 465792 140924 465798
rect 140872 465734 140924 465740
rect 136640 458992 136692 458998
rect 136640 458934 136692 458940
rect 142172 458930 142200 475118
rect 142264 463146 142292 480023
rect 142632 475182 142660 480023
rect 142620 475176 142672 475182
rect 142620 475118 142672 475124
rect 143000 470594 143028 480023
rect 143632 475312 143684 475318
rect 143632 475254 143684 475260
rect 142356 470566 143028 470594
rect 142356 463214 142384 470566
rect 143644 468489 143672 475254
rect 143828 472666 143856 480037
rect 143920 480023 144302 480051
rect 144472 480023 144762 480051
rect 143816 472660 143868 472666
rect 143816 472602 143868 472608
rect 143920 470594 143948 480023
rect 144472 475318 144500 480023
rect 145116 478145 145144 480037
rect 145576 478281 145604 480037
rect 145562 478272 145618 478281
rect 145562 478207 145618 478216
rect 145102 478136 145158 478145
rect 145102 478071 145158 478080
rect 144460 475312 144512 475318
rect 144460 475254 144512 475260
rect 146036 471345 146064 480037
rect 146404 480023 146510 480051
rect 146680 480023 146970 480051
rect 146300 475312 146352 475318
rect 146300 475254 146352 475260
rect 146022 471336 146078 471345
rect 146022 471271 146078 471280
rect 143736 470566 143948 470594
rect 143630 468480 143686 468489
rect 143630 468415 143686 468424
rect 142344 463208 142396 463214
rect 142344 463150 142396 463156
rect 142252 463140 142304 463146
rect 142252 463082 142304 463088
rect 143736 460329 143764 470566
rect 146312 462913 146340 475254
rect 146404 470642 146432 480023
rect 146680 475318 146708 480023
rect 147324 478553 147352 480037
rect 147310 478544 147366 478553
rect 147310 478479 147366 478488
rect 146668 475312 146720 475318
rect 146668 475254 146720 475260
rect 147784 472666 147812 480037
rect 148244 478417 148272 480037
rect 148336 480023 148718 480051
rect 148230 478408 148286 478417
rect 148230 478343 148286 478352
rect 147772 472660 147824 472666
rect 147772 472602 147824 472608
rect 146404 470614 146524 470642
rect 146496 463049 146524 470614
rect 148336 470594 148364 480023
rect 149164 478378 149192 480037
rect 149532 478718 149560 480037
rect 149992 478854 150020 480037
rect 149980 478848 150032 478854
rect 149980 478790 150032 478796
rect 149520 478712 149572 478718
rect 149520 478654 149572 478660
rect 149152 478372 149204 478378
rect 149152 478314 149204 478320
rect 150452 474201 150480 480037
rect 150544 480023 150926 480051
rect 150438 474192 150494 474201
rect 150438 474127 150494 474136
rect 150544 470594 150572 480023
rect 151280 478446 151308 480037
rect 151268 478440 151320 478446
rect 151268 478382 151320 478388
rect 151740 471209 151768 480037
rect 152200 478582 152228 480037
rect 152188 478576 152240 478582
rect 152188 478518 152240 478524
rect 152660 472569 152688 480037
rect 153120 476785 153148 480037
rect 153488 478650 153516 480037
rect 153580 480023 153962 480051
rect 154040 480023 154422 480051
rect 153476 478644 153528 478650
rect 153476 478586 153528 478592
rect 153106 476776 153162 476785
rect 153106 476711 153162 476720
rect 153580 475402 153608 480023
rect 153212 475374 153608 475402
rect 152646 472560 152702 472569
rect 152646 472495 152702 472504
rect 151726 471200 151782 471209
rect 151726 471135 151782 471144
rect 147692 470566 148364 470594
rect 150452 470566 150572 470594
rect 147692 467129 147720 470566
rect 150452 468625 150480 470566
rect 150438 468616 150494 468625
rect 150438 468551 150494 468560
rect 147678 467120 147734 467129
rect 147678 467055 147734 467064
rect 146482 463040 146538 463049
rect 146482 462975 146538 462984
rect 146298 462904 146354 462913
rect 146298 462839 146354 462848
rect 143722 460320 143778 460329
rect 143722 460255 143778 460264
rect 153212 460193 153240 475374
rect 154040 470594 154068 480023
rect 154868 478514 154896 480037
rect 154960 480023 155342 480051
rect 154856 478508 154908 478514
rect 154856 478450 154908 478456
rect 154960 470594 154988 480023
rect 155696 475561 155724 480037
rect 156156 478786 156184 480037
rect 156248 480023 156630 480051
rect 156144 478780 156196 478786
rect 156144 478722 156196 478728
rect 155682 475552 155738 475561
rect 155682 475487 155738 475496
rect 156248 470594 156276 480023
rect 157076 478310 157104 480037
rect 157352 480023 157458 480051
rect 157536 480023 157918 480051
rect 157064 478304 157116 478310
rect 157064 478246 157116 478252
rect 153304 470566 154068 470594
rect 154592 470566 154988 470594
rect 155972 470566 156276 470594
rect 153304 469849 153332 470566
rect 153290 469840 153346 469849
rect 153290 469775 153346 469784
rect 154592 467265 154620 470566
rect 155972 469985 156000 470566
rect 155958 469976 156014 469985
rect 155958 469911 156014 469920
rect 154578 467256 154634 467265
rect 154578 467191 154634 467200
rect 157352 460465 157380 480023
rect 157536 470594 157564 480023
rect 158364 478242 158392 480037
rect 158996 480072 159048 480078
rect 158838 480023 158868 480051
rect 158720 480014 158772 480020
rect 158352 478236 158404 478242
rect 158352 478178 158404 478184
rect 157444 470566 157564 470594
rect 157444 468761 157472 470566
rect 157430 468752 157486 468761
rect 157430 468687 157486 468696
rect 158732 461718 158760 480014
rect 158840 479890 158868 480023
rect 187792 480072 187844 480078
rect 159048 480023 159298 480051
rect 158996 480014 159048 480020
rect 158840 479862 159036 479890
rect 159008 470642 159036 479862
rect 159652 474026 159680 480037
rect 160112 475794 160140 480037
rect 160204 480023 160586 480051
rect 160664 480023 161046 480051
rect 161506 480023 161536 480051
rect 160100 475788 160152 475794
rect 160100 475730 160152 475736
rect 160204 475402 160232 480023
rect 160112 475374 160232 475402
rect 159640 474020 159692 474026
rect 159640 473962 159692 473968
rect 158840 470614 159036 470642
rect 158840 470594 158868 470614
rect 158824 470566 158868 470594
rect 158824 469878 158852 470566
rect 158812 469872 158864 469878
rect 158812 469814 158864 469820
rect 160112 466041 160140 475374
rect 160664 470594 160692 480023
rect 161508 479874 161536 480023
rect 161584 480023 161874 480051
rect 161952 480023 162334 480051
rect 162504 480023 162794 480051
rect 161496 479868 161548 479874
rect 161496 479810 161548 479816
rect 161584 475538 161612 480023
rect 160204 470566 160692 470594
rect 161492 475510 161612 475538
rect 160204 467226 160232 470566
rect 160192 467220 160244 467226
rect 160192 467162 160244 467168
rect 160098 466032 160154 466041
rect 160098 465967 160154 465976
rect 161492 463282 161520 475510
rect 161952 475402 161980 480023
rect 162032 479868 162084 479874
rect 162032 479810 162084 479816
rect 161584 475374 161980 475402
rect 161584 463350 161612 475374
rect 162044 471374 162072 479810
rect 162032 471368 162084 471374
rect 162032 471310 162084 471316
rect 162504 470594 162532 480023
rect 163240 476950 163268 480037
rect 163608 478689 163636 480037
rect 163594 478680 163650 478689
rect 163594 478615 163650 478624
rect 163228 476944 163280 476950
rect 163228 476886 163280 476892
rect 164068 476882 164096 480037
rect 164252 480023 164542 480051
rect 164620 480023 165002 480051
rect 164056 476876 164108 476882
rect 164056 476818 164108 476824
rect 161676 470566 162532 470594
rect 161676 465905 161704 470566
rect 161662 465896 161718 465905
rect 161662 465831 161718 465840
rect 161572 463344 161624 463350
rect 161572 463286 161624 463292
rect 161480 463276 161532 463282
rect 161480 463218 161532 463224
rect 158720 461712 158772 461718
rect 158720 461654 158772 461660
rect 157338 460456 157394 460465
rect 157338 460391 157394 460400
rect 153198 460184 153254 460193
rect 153198 460119 153254 460128
rect 164252 458969 164280 480023
rect 164620 470594 164648 480023
rect 165448 475862 165476 480037
rect 165724 480023 165830 480051
rect 165436 475856 165488 475862
rect 165436 475798 165488 475804
rect 165620 475312 165672 475318
rect 165620 475254 165672 475260
rect 164344 470566 164648 470594
rect 164344 460601 164372 470566
rect 164330 460592 164386 460601
rect 164330 460527 164386 460536
rect 165632 460358 165660 475254
rect 165724 468654 165752 480023
rect 166276 478106 166304 480037
rect 166368 480023 166750 480051
rect 167012 480023 167210 480051
rect 166264 478100 166316 478106
rect 166264 478042 166316 478048
rect 166368 475318 166396 480023
rect 166356 475312 166408 475318
rect 166356 475254 166408 475260
rect 165712 468648 165764 468654
rect 165712 468590 165764 468596
rect 167012 460737 167040 480023
rect 167656 477018 167684 480037
rect 167748 480023 168038 480051
rect 167644 477012 167696 477018
rect 167644 476954 167696 476960
rect 167748 470594 167776 480023
rect 168380 475312 168432 475318
rect 168380 475254 168432 475260
rect 167196 470566 167776 470594
rect 167196 460873 167224 470566
rect 167182 460864 167238 460873
rect 167182 460799 167238 460808
rect 166998 460728 167054 460737
rect 166998 460663 167054 460672
rect 165620 460352 165672 460358
rect 165620 460294 165672 460300
rect 168392 459105 168420 475254
rect 168484 460426 168512 480037
rect 168576 480023 168958 480051
rect 169128 480023 169418 480051
rect 169772 480023 169878 480051
rect 168472 460420 168524 460426
rect 168472 460362 168524 460368
rect 168576 459377 168604 480023
rect 169024 478032 169076 478038
rect 169024 477974 169076 477980
rect 169036 468722 169064 477974
rect 169128 475318 169156 480023
rect 169116 475312 169168 475318
rect 169116 475254 169168 475260
rect 169024 468716 169076 468722
rect 169024 468658 169076 468664
rect 169772 463418 169800 480023
rect 170232 478825 170260 480037
rect 170324 480023 170706 480051
rect 170218 478816 170274 478825
rect 170218 478751 170274 478760
rect 170324 470594 170352 480023
rect 169864 470566 170352 470594
rect 169864 466177 169892 470566
rect 169850 466168 169906 466177
rect 169850 466103 169906 466112
rect 169760 463412 169812 463418
rect 169760 463354 169812 463360
rect 168562 459368 168618 459377
rect 168562 459303 168618 459312
rect 171152 459241 171180 480037
rect 171612 474337 171640 480037
rect 171704 480023 171994 480051
rect 171598 474328 171654 474337
rect 171598 474263 171654 474272
rect 171704 470594 171732 480023
rect 172440 472734 172468 480037
rect 172624 480023 172914 480051
rect 172992 480023 173374 480051
rect 173544 480023 173834 480051
rect 174004 480023 174202 480051
rect 174280 480023 174662 480051
rect 174740 480023 175122 480051
rect 175384 480023 175582 480051
rect 172520 475312 172572 475318
rect 172520 475254 172572 475260
rect 172428 472728 172480 472734
rect 172428 472670 172480 472676
rect 171244 470566 171732 470594
rect 171244 463185 171272 470566
rect 171230 463176 171286 463185
rect 171230 463111 171286 463120
rect 172532 459513 172560 475254
rect 172624 464409 172652 480023
rect 172992 470594 173020 480023
rect 173544 475318 173572 480023
rect 173532 475312 173584 475318
rect 173532 475254 173584 475260
rect 173900 475312 173952 475318
rect 173900 475254 173952 475260
rect 172716 470566 173020 470594
rect 172716 470121 172744 470566
rect 172702 470112 172758 470121
rect 172702 470047 172758 470056
rect 172610 464400 172666 464409
rect 172610 464335 172666 464344
rect 172518 459504 172574 459513
rect 172518 459439 172574 459448
rect 171138 459232 171194 459241
rect 171138 459167 171194 459176
rect 173912 459134 173940 475254
rect 174004 459270 174032 480023
rect 174280 475318 174308 480023
rect 174268 475312 174320 475318
rect 174268 475254 174320 475260
rect 174740 470594 174768 480023
rect 175280 475312 175332 475318
rect 175280 475254 175332 475260
rect 174096 470566 174768 470594
rect 174096 466070 174124 470566
rect 175292 467294 175320 475254
rect 175384 468790 175412 480023
rect 176028 474094 176056 480037
rect 176120 480023 176410 480051
rect 176672 480023 176870 480051
rect 176948 480023 177330 480051
rect 177408 480023 177790 480051
rect 176120 475318 176148 480023
rect 176108 475312 176160 475318
rect 176108 475254 176160 475260
rect 176016 474088 176068 474094
rect 176016 474030 176068 474036
rect 175372 468784 175424 468790
rect 175372 468726 175424 468732
rect 175280 467288 175332 467294
rect 175280 467230 175332 467236
rect 174084 466064 174136 466070
rect 174084 466006 174136 466012
rect 173992 459264 174044 459270
rect 173992 459206 174044 459212
rect 176672 459202 176700 480023
rect 176948 475402 176976 480023
rect 176764 475374 176976 475402
rect 176764 462058 176792 475374
rect 177408 470594 177436 480023
rect 178144 475998 178172 480037
rect 178236 480023 178618 480051
rect 178696 480023 179078 480051
rect 179432 480023 179538 480051
rect 178132 475992 178184 475998
rect 178132 475934 178184 475940
rect 178236 475402 178264 480023
rect 176856 470566 177436 470594
rect 178052 475374 178264 475402
rect 176856 463690 176884 470566
rect 176844 463684 176896 463690
rect 176844 463626 176896 463632
rect 178052 463486 178080 475374
rect 178696 470594 178724 480023
rect 178144 470566 178724 470594
rect 178144 469946 178172 470566
rect 178132 469940 178184 469946
rect 178132 469882 178184 469888
rect 178040 463480 178092 463486
rect 178040 463422 178092 463428
rect 178316 462324 178368 462330
rect 178316 462266 178368 462272
rect 176752 462052 176804 462058
rect 176752 461994 176804 462000
rect 178328 461417 178356 462266
rect 178314 461408 178370 461417
rect 178314 461343 178370 461352
rect 178328 461038 178356 461343
rect 178316 461032 178368 461038
rect 178316 460974 178368 460980
rect 179432 460834 179460 480023
rect 179984 472705 180012 480037
rect 179970 472696 180026 472705
rect 179970 472631 180026 472640
rect 180352 471442 180380 480037
rect 180340 471436 180392 471442
rect 180340 471378 180392 471384
rect 179512 467152 179564 467158
rect 179512 467094 179564 467100
rect 179524 461786 179552 467094
rect 179512 461780 179564 461786
rect 179512 461722 179564 461728
rect 179524 461689 179552 461722
rect 179510 461680 179566 461689
rect 179510 461615 179566 461624
rect 179420 460828 179472 460834
rect 179420 460770 179472 460776
rect 180812 460562 180840 480037
rect 180904 480023 181286 480051
rect 181456 480023 181746 480051
rect 180904 461854 180932 480023
rect 181456 470594 181484 480023
rect 180996 470566 181484 470594
rect 180996 463554 181024 470566
rect 180984 463548 181036 463554
rect 180984 463490 181036 463496
rect 180892 461848 180944 461854
rect 180892 461790 180944 461796
rect 180800 460556 180852 460562
rect 180800 460498 180852 460504
rect 182192 459338 182220 480037
rect 182376 480023 182574 480051
rect 182744 480023 183034 480051
rect 183112 480023 183494 480051
rect 183572 480023 183954 480051
rect 184032 480023 184322 480051
rect 184400 480023 184782 480051
rect 184952 480023 185242 480051
rect 182272 472932 182324 472938
rect 182272 472874 182324 472880
rect 182284 461922 182312 472874
rect 182376 462874 182404 480023
rect 182744 470594 182772 480023
rect 183112 472938 183140 480023
rect 183100 472932 183152 472938
rect 183100 472874 183152 472880
rect 182468 470566 182772 470594
rect 182468 466206 182496 470566
rect 182456 466200 182508 466206
rect 182456 466142 182508 466148
rect 182364 462868 182416 462874
rect 182364 462810 182416 462816
rect 182272 461916 182324 461922
rect 182272 461858 182324 461864
rect 183572 460698 183600 480023
rect 184032 475402 184060 480023
rect 183664 475374 184060 475402
rect 183664 466342 183692 475374
rect 184400 470594 184428 480023
rect 183756 470566 184428 470594
rect 183652 466336 183704 466342
rect 183652 466278 183704 466284
rect 183756 466274 183784 470566
rect 183744 466268 183796 466274
rect 183744 466210 183796 466216
rect 184952 461990 184980 480023
rect 185584 478168 185636 478174
rect 185584 478110 185636 478116
rect 185596 462194 185624 478110
rect 185688 478009 185716 480037
rect 186148 478038 186176 480037
rect 186424 480023 186530 480051
rect 186136 478032 186188 478038
rect 185674 478000 185730 478009
rect 186136 477974 186188 477980
rect 185674 477935 185730 477944
rect 186424 467158 186452 480023
rect 186976 478038 187004 480037
rect 187160 480023 187450 480051
rect 186504 478032 186556 478038
rect 186504 477974 186556 477980
rect 186964 478032 187016 478038
rect 186964 477974 187016 477980
rect 186516 475930 186544 477974
rect 186504 475924 186556 475930
rect 186504 475866 186556 475872
rect 186412 467152 186464 467158
rect 186412 467094 186464 467100
rect 187160 466454 187188 480023
rect 188068 480072 188120 480078
rect 187910 480023 187940 480051
rect 187792 480014 187844 480020
rect 187700 470348 187752 470354
rect 187700 470290 187752 470296
rect 186332 466426 187188 466454
rect 186332 463321 186360 466426
rect 186318 463312 186374 463321
rect 186318 463247 186374 463256
rect 185584 462188 185636 462194
rect 185584 462130 185636 462136
rect 184940 461984 184992 461990
rect 184940 461926 184992 461932
rect 183560 460692 183612 460698
rect 183560 460634 183612 460640
rect 187712 459542 187740 470290
rect 187804 460630 187832 480014
rect 187912 479890 187940 480023
rect 196298 480066 196664 480094
rect 188120 480023 188370 480051
rect 188448 480023 188738 480051
rect 189092 480023 189198 480051
rect 189276 480023 189658 480051
rect 189736 480023 190118 480051
rect 188068 480014 188120 480020
rect 187912 479862 188108 479890
rect 188080 466454 188108 479862
rect 188448 470354 188476 480023
rect 188436 470348 188488 470354
rect 188436 470290 188488 470296
rect 187896 466426 188108 466454
rect 187896 466313 187924 466426
rect 187882 466304 187938 466313
rect 187882 466239 187938 466248
rect 189092 462942 189120 480023
rect 189172 471232 189224 471238
rect 189172 471174 189224 471180
rect 189184 466410 189212 471174
rect 189172 466404 189224 466410
rect 189172 466346 189224 466352
rect 189276 466138 189304 480023
rect 189736 471238 189764 480023
rect 189724 471232 189776 471238
rect 189724 471174 189776 471180
rect 189264 466132 189316 466138
rect 189264 466074 189316 466080
rect 189080 462936 189132 462942
rect 189080 462878 189132 462884
rect 187792 460624 187844 460630
rect 187792 460566 187844 460572
rect 187700 459536 187752 459542
rect 187700 459478 187752 459484
rect 190472 459406 190500 480037
rect 190564 480023 190946 480051
rect 191024 480023 191406 480051
rect 191866 480023 192156 480051
rect 190564 462126 190592 480023
rect 191024 466454 191052 480023
rect 192128 473006 192156 480023
rect 192220 480023 192326 480051
rect 192404 480023 192694 480051
rect 192864 480023 193154 480051
rect 193416 480023 193614 480051
rect 193784 480023 194074 480051
rect 194152 480023 194534 480051
rect 192116 473000 192168 473006
rect 192116 472942 192168 472948
rect 192024 471232 192076 471238
rect 192024 471174 192076 471180
rect 191840 471164 191892 471170
rect 191840 471106 191892 471112
rect 190656 466426 191052 466454
rect 190656 465526 190684 466426
rect 190644 465520 190696 465526
rect 190644 465462 190696 465468
rect 190552 462120 190604 462126
rect 190552 462062 190604 462068
rect 190918 461000 190974 461009
rect 190918 460935 190920 460944
rect 190972 460935 190974 460944
rect 190920 460906 190972 460912
rect 191852 459474 191880 471106
rect 192036 465662 192064 471174
rect 192024 465656 192076 465662
rect 192024 465598 192076 465604
rect 192220 463694 192248 480023
rect 192404 471170 192432 480023
rect 192668 473000 192720 473006
rect 192668 472942 192720 472948
rect 192392 471164 192444 471170
rect 192392 471106 192444 471112
rect 192680 465458 192708 472942
rect 192864 471238 192892 480023
rect 192852 471232 192904 471238
rect 192852 471174 192904 471180
rect 193220 471232 193272 471238
rect 193220 471174 193272 471180
rect 192668 465452 192720 465458
rect 192668 465394 192720 465400
rect 191944 463666 192248 463694
rect 191840 459468 191892 459474
rect 191840 459410 191892 459416
rect 190460 459400 190512 459406
rect 190460 459342 190512 459348
rect 182180 459332 182232 459338
rect 182180 459274 182232 459280
rect 176660 459196 176712 459202
rect 176660 459138 176712 459144
rect 173900 459128 173952 459134
rect 168378 459096 168434 459105
rect 173900 459070 173952 459076
rect 168378 459031 168434 459040
rect 164238 458960 164294 458969
rect 134064 458924 134116 458930
rect 134064 458866 134116 458872
rect 142160 458924 142212 458930
rect 164238 458895 164294 458904
rect 142160 458866 142212 458872
rect 109316 458798 109368 458804
rect 125690 458824 125746 458833
rect 69018 458759 69074 458768
rect 191944 458794 191972 463666
rect 193232 460494 193260 471174
rect 193312 471164 193364 471170
rect 193312 471106 193364 471112
rect 193324 462806 193352 471106
rect 193416 463622 193444 480023
rect 193784 471238 193812 480023
rect 193772 471232 193824 471238
rect 193772 471174 193824 471180
rect 194152 471170 194180 480023
rect 194888 477562 194916 480037
rect 195348 477630 195376 480037
rect 195440 480023 195822 480051
rect 195336 477624 195388 477630
rect 195336 477566 195388 477572
rect 194876 477556 194928 477562
rect 194876 477498 194928 477504
rect 194140 471164 194192 471170
rect 194140 471106 194192 471112
rect 195440 466454 195468 480023
rect 194612 466426 195468 466454
rect 193404 463616 193456 463622
rect 193404 463558 193456 463564
rect 193312 462800 193364 462806
rect 193312 462742 193364 462748
rect 193220 460488 193272 460494
rect 193220 460430 193272 460436
rect 194612 459678 194640 466426
rect 194600 459672 194652 459678
rect 194600 459614 194652 459620
rect 125690 458759 125746 458768
rect 191932 458788 191984 458794
rect 191932 458730 191984 458736
rect 60740 374944 60792 374950
rect 60740 374886 60792 374892
rect 60752 353394 60780 374886
rect 158534 374640 158590 374649
rect 158534 374575 158590 374584
rect 165986 374640 166042 374649
rect 165986 374575 165988 374584
rect 158548 374542 158576 374575
rect 166040 374575 166042 374584
rect 195886 374640 195942 374649
rect 195886 374575 195942 374584
rect 165988 374546 166040 374552
rect 158536 374536 158588 374542
rect 105450 374504 105506 374513
rect 105450 374439 105506 374448
rect 116030 374504 116086 374513
rect 116030 374439 116086 374448
rect 140962 374504 141018 374513
rect 140962 374439 141018 374448
rect 143538 374504 143594 374513
rect 143538 374439 143594 374448
rect 156510 374504 156566 374513
rect 158536 374478 158588 374484
rect 160926 374504 160982 374513
rect 156510 374439 156512 374448
rect 105464 374134 105492 374439
rect 105452 374128 105504 374134
rect 105452 374070 105504 374076
rect 116044 374066 116072 374439
rect 139214 374096 139270 374105
rect 116032 374060 116084 374066
rect 140976 374066 141004 374439
rect 143552 374202 143580 374439
rect 156564 374439 156566 374448
rect 160926 374439 160982 374448
rect 163410 374504 163466 374513
rect 163410 374439 163466 374448
rect 156512 374410 156564 374416
rect 146206 374368 146262 374377
rect 146206 374303 146262 374312
rect 148966 374368 149022 374377
rect 160940 374338 160968 374439
rect 163424 374406 163452 374439
rect 163412 374400 163464 374406
rect 163412 374342 163464 374348
rect 148966 374303 149022 374312
rect 160928 374332 160980 374338
rect 146220 374270 146248 374303
rect 146208 374264 146260 374270
rect 146208 374206 146260 374212
rect 143540 374196 143592 374202
rect 143540 374138 143592 374144
rect 148980 374134 149008 374303
rect 160928 374274 160980 374280
rect 148968 374128 149020 374134
rect 148968 374070 149020 374076
rect 139214 374031 139270 374040
rect 140964 374060 141016 374066
rect 116032 374002 116084 374008
rect 139228 373862 139256 374031
rect 140964 374002 141016 374008
rect 96068 373856 96120 373862
rect 96068 373798 96120 373804
rect 139216 373856 139268 373862
rect 139216 373798 139268 373804
rect 96080 373697 96108 373798
rect 118332 373788 118384 373794
rect 118332 373730 118384 373736
rect 136456 373788 136508 373794
rect 136456 373730 136508 373736
rect 103520 373720 103572 373726
rect 95054 373688 95110 373697
rect 95054 373623 95110 373632
rect 96066 373688 96122 373697
rect 96066 373623 96122 373632
rect 103518 373688 103520 373697
rect 118344 373697 118372 373730
rect 133696 373720 133748 373726
rect 103572 373688 103574 373697
rect 103518 373623 103574 373632
rect 107842 373688 107898 373697
rect 107842 373623 107898 373632
rect 113546 373688 113602 373697
rect 113546 373623 113548 373632
rect 93674 373416 93730 373425
rect 93674 373351 93730 373360
rect 93688 373318 93716 373351
rect 95068 373318 95096 373623
rect 107856 373590 107884 373623
rect 113600 373623 113602 373632
rect 118330 373688 118386 373697
rect 118330 373623 118386 373632
rect 121366 373688 121422 373697
rect 133696 373662 133748 373668
rect 121366 373623 121422 373632
rect 131028 373652 131080 373658
rect 113548 373594 113600 373600
rect 107844 373584 107896 373590
rect 107844 373526 107896 373532
rect 110418 373552 110474 373561
rect 110418 373487 110474 373496
rect 110432 373454 110460 373487
rect 121380 373454 121408 373623
rect 131028 373594 131080 373600
rect 124128 373584 124180 373590
rect 124126 373552 124128 373561
rect 131040 373561 131068 373594
rect 133708 373561 133736 373662
rect 136468 373561 136496 373730
rect 124180 373552 124182 373561
rect 124126 373487 124182 373496
rect 125690 373552 125746 373561
rect 125690 373487 125692 373496
rect 125744 373487 125746 373496
rect 128910 373552 128966 373561
rect 128910 373487 128912 373496
rect 125692 373458 125744 373464
rect 128964 373487 128966 373496
rect 131026 373552 131082 373561
rect 131026 373487 131082 373496
rect 133694 373552 133750 373561
rect 133694 373487 133750 373496
rect 136454 373552 136510 373561
rect 136454 373487 136510 373496
rect 151726 373552 151782 373561
rect 151726 373487 151782 373496
rect 154118 373552 154174 373561
rect 154118 373487 154174 373496
rect 128912 373458 128964 373464
rect 110420 373448 110472 373454
rect 98274 373416 98330 373425
rect 110420 373390 110472 373396
rect 121368 373448 121420 373454
rect 121368 373390 121420 373396
rect 98274 373351 98276 373360
rect 98328 373351 98330 373360
rect 99380 373380 99432 373386
rect 98276 373322 98328 373328
rect 99380 373322 99432 373328
rect 93676 373312 93728 373318
rect 88338 373280 88394 373289
rect 93676 373254 93728 373260
rect 95056 373312 95108 373318
rect 95056 373254 95108 373260
rect 95974 373280 96030 373289
rect 88338 373215 88394 373224
rect 95974 373215 96030 373224
rect 88352 373182 88380 373215
rect 88340 373176 88392 373182
rect 88340 373118 88392 373124
rect 90178 373144 90234 373153
rect 90178 373079 90180 373088
rect 90232 373079 90234 373088
rect 92386 373144 92442 373153
rect 92386 373079 92442 373088
rect 90180 373050 90232 373056
rect 62118 372736 62174 372745
rect 62118 372671 62174 372680
rect 60740 353388 60792 353394
rect 60740 353330 60792 353336
rect 62132 353326 62160 372671
rect 77206 372600 77262 372609
rect 77206 372535 77262 372544
rect 85486 372600 85542 372609
rect 85486 372535 85542 372544
rect 86590 372600 86646 372609
rect 86590 372535 86646 372544
rect 88062 372600 88118 372609
rect 88062 372535 88118 372544
rect 89350 372600 89406 372609
rect 89350 372535 89352 372544
rect 77220 372366 77248 372535
rect 78494 372464 78550 372473
rect 78494 372399 78550 372408
rect 79966 372464 80022 372473
rect 79966 372399 80022 372408
rect 85118 372464 85174 372473
rect 85118 372399 85174 372408
rect 77208 372360 77260 372366
rect 77208 372302 77260 372308
rect 77022 372192 77078 372201
rect 77022 372127 77078 372136
rect 77036 370326 77064 372127
rect 78508 372026 78536 372399
rect 78496 372020 78548 372026
rect 78496 371962 78548 371968
rect 78508 371414 78536 371962
rect 79980 371890 80008 372399
rect 80518 372328 80574 372337
rect 80518 372263 80574 372272
rect 81898 372328 81954 372337
rect 81898 372263 81954 372272
rect 79968 371884 80020 371890
rect 79968 371826 80020 371832
rect 79980 371482 80008 371826
rect 79968 371476 80020 371482
rect 79968 371418 80020 371424
rect 78496 371408 78548 371414
rect 78496 371350 78548 371356
rect 80532 371346 80560 372263
rect 81912 371550 81940 372263
rect 83830 371920 83886 371929
rect 83830 371855 83886 371864
rect 81900 371544 81952 371550
rect 81900 371486 81952 371492
rect 82452 371544 82504 371550
rect 82452 371486 82504 371492
rect 80520 371340 80572 371346
rect 80520 371282 80572 371288
rect 82464 371278 82492 371486
rect 82452 371272 82504 371278
rect 82452 371214 82504 371220
rect 77024 370320 77076 370326
rect 77024 370262 77076 370268
rect 83844 369850 83872 371855
rect 85132 371550 85160 372399
rect 85500 371890 85528 372535
rect 86604 372162 86632 372535
rect 86592 372156 86644 372162
rect 86592 372098 86644 372104
rect 85488 371884 85540 371890
rect 85488 371826 85540 371832
rect 88076 371822 88104 372535
rect 89404 372535 89406 372544
rect 90086 372600 90142 372609
rect 90086 372535 90142 372544
rect 92202 372600 92258 372609
rect 92202 372535 92258 372544
rect 89352 372506 89404 372512
rect 90100 372434 90128 372535
rect 90088 372428 90140 372434
rect 90088 372370 90140 372376
rect 88064 371816 88116 371822
rect 88064 371758 88116 371764
rect 92216 371686 92244 372535
rect 92400 372502 92428 373079
rect 95988 372638 96016 373215
rect 95976 372632 96028 372638
rect 93582 372600 93638 372609
rect 95976 372574 96028 372580
rect 93582 372535 93638 372544
rect 92388 372496 92440 372502
rect 92388 372438 92440 372444
rect 93596 371754 93624 372535
rect 99392 372366 99420 373322
rect 100850 373280 100906 373289
rect 151740 373250 151768 373487
rect 100850 373215 100852 373224
rect 100904 373215 100906 373224
rect 151728 373244 151780 373250
rect 100852 373186 100904 373192
rect 151728 373186 151780 373192
rect 154132 373182 154160 373487
rect 154120 373176 154172 373182
rect 154120 373118 154172 373124
rect 108854 372600 108910 372609
rect 108854 372535 108910 372544
rect 114006 372600 114062 372609
rect 114006 372535 114062 372544
rect 183190 372600 183246 372609
rect 183190 372535 183246 372544
rect 102782 372464 102838 372473
rect 102782 372399 102838 372408
rect 99380 372360 99432 372366
rect 99380 372302 99432 372308
rect 102046 372328 102102 372337
rect 102046 372263 102102 372272
rect 93584 371748 93636 371754
rect 93584 371690 93636 371696
rect 92204 371680 92256 371686
rect 92204 371622 92256 371628
rect 97722 371648 97778 371657
rect 97722 371583 97778 371592
rect 99286 371648 99342 371657
rect 99286 371583 99342 371592
rect 100114 371648 100170 371657
rect 100114 371583 100170 371592
rect 85120 371544 85172 371550
rect 85120 371486 85172 371492
rect 83832 369844 83884 369850
rect 83832 369786 83884 369792
rect 97736 369170 97764 371583
rect 99300 369238 99328 371583
rect 100128 369306 100156 371583
rect 101034 371512 101090 371521
rect 101034 371447 101090 371456
rect 100116 369300 100168 369306
rect 100116 369242 100168 369248
rect 99288 369232 99340 369238
rect 99288 369174 99340 369180
rect 97724 369164 97776 369170
rect 97724 369106 97776 369112
rect 101048 368830 101076 371447
rect 102060 370530 102088 372263
rect 102796 371006 102824 372399
rect 108868 371958 108896 372535
rect 108856 371952 108908 371958
rect 104622 371920 104678 371929
rect 108856 371894 108908 371900
rect 114020 371890 114048 372535
rect 117962 372328 118018 372337
rect 117962 372263 118018 372272
rect 117976 372065 118004 372263
rect 117962 372056 118018 372065
rect 117962 371991 118018 372000
rect 104622 371855 104678 371864
rect 106188 371884 106240 371890
rect 102784 371000 102836 371006
rect 102784 370942 102836 370948
rect 102048 370524 102100 370530
rect 102048 370466 102100 370472
rect 104636 369753 104664 371855
rect 106188 371826 106240 371832
rect 114008 371884 114060 371890
rect 114008 371826 114060 371832
rect 105910 371784 105966 371793
rect 105910 371719 105966 371728
rect 104622 369744 104678 369753
rect 104622 369679 104678 369688
rect 105924 369617 105952 371719
rect 105910 369608 105966 369617
rect 105910 369543 105966 369552
rect 106200 369034 106228 371826
rect 182822 371512 182878 371521
rect 182822 371447 182878 371456
rect 107566 371376 107622 371385
rect 107566 371311 107622 371320
rect 106188 369028 106240 369034
rect 106188 368970 106240 368976
rect 101036 368824 101088 368830
rect 101036 368766 101088 368772
rect 107580 367810 107608 371311
rect 182836 371142 182864 371447
rect 183204 371210 183232 372535
rect 183192 371204 183244 371210
rect 183192 371146 183244 371152
rect 182824 371136 182876 371142
rect 182824 371078 182876 371084
rect 107568 367804 107620 367810
rect 107568 367746 107620 367752
rect 182836 356726 182864 371078
rect 182824 356720 182876 356726
rect 182824 356662 182876 356668
rect 191380 356040 191432 356046
rect 191380 355982 191432 355988
rect 179788 355972 179840 355978
rect 179788 355914 179840 355920
rect 179800 355337 179828 355914
rect 191392 355337 191420 355982
rect 195900 355978 195928 374575
rect 196636 370666 196664 480066
rect 248420 480072 248472 480078
rect 196742 480023 196848 480051
rect 196716 471300 196768 471306
rect 196716 471242 196768 471248
rect 196728 370802 196756 471242
rect 196716 370796 196768 370802
rect 196716 370738 196768 370744
rect 196820 370734 196848 480023
rect 196912 480023 197110 480051
rect 196912 471306 196940 480023
rect 197360 478372 197412 478378
rect 197360 478314 197412 478320
rect 197372 477737 197400 478314
rect 197358 477728 197414 477737
rect 197358 477663 197414 477672
rect 196992 477556 197044 477562
rect 196992 477498 197044 477504
rect 196900 471300 196952 471306
rect 196900 471242 196952 471248
rect 196898 465760 196954 465769
rect 196898 465695 196954 465704
rect 196808 370728 196860 370734
rect 196808 370670 196860 370676
rect 196624 370660 196676 370666
rect 196624 370602 196676 370608
rect 195888 355972 195940 355978
rect 195888 355914 195940 355920
rect 179786 355328 179842 355337
rect 179786 355263 179842 355272
rect 191378 355328 191434 355337
rect 191378 355263 191434 355272
rect 195900 355230 195928 355914
rect 195888 355224 195940 355230
rect 195888 355166 195940 355172
rect 178590 354784 178646 354793
rect 178590 354719 178592 354728
rect 178644 354719 178646 354728
rect 178592 354690 178644 354696
rect 62120 353320 62172 353326
rect 62120 353262 62172 353268
rect 110970 269920 111026 269929
rect 110970 269855 111026 269864
rect 148506 269920 148562 269929
rect 148506 269855 148562 269864
rect 60096 269680 60148 269686
rect 60096 269622 60148 269628
rect 83094 269648 83150 269657
rect 60108 268734 60136 269622
rect 83094 269583 83150 269592
rect 91282 269648 91338 269657
rect 91282 269583 91338 269592
rect 93582 269648 93638 269657
rect 93582 269583 93638 269592
rect 94502 269648 94558 269657
rect 110984 269618 111012 269855
rect 133418 269784 133474 269793
rect 133418 269719 133474 269728
rect 135902 269784 135958 269793
rect 135902 269719 135958 269728
rect 138478 269784 138534 269793
rect 138478 269719 138534 269728
rect 140870 269784 140926 269793
rect 148520 269754 148548 269855
rect 140870 269719 140926 269728
rect 148508 269748 148560 269754
rect 94502 269583 94558 269592
rect 110972 269612 111024 269618
rect 62120 269000 62172 269006
rect 62120 268942 62172 268948
rect 60096 268728 60148 268734
rect 60096 268670 60148 268676
rect 62132 249014 62160 268942
rect 76010 268832 76066 268841
rect 76010 268767 76066 268776
rect 77114 268832 77170 268841
rect 77114 268767 77170 268776
rect 66260 268184 66312 268190
rect 66260 268126 66312 268132
rect 66272 267073 66300 268126
rect 76024 268122 76052 268767
rect 77128 268258 77156 268767
rect 77116 268252 77168 268258
rect 77116 268194 77168 268200
rect 76012 268116 76064 268122
rect 76012 268058 76064 268064
rect 79324 268116 79376 268122
rect 79324 268058 79376 268064
rect 66258 267064 66314 267073
rect 66258 266999 66314 267008
rect 77298 267064 77354 267073
rect 77298 266999 77354 267008
rect 78678 267064 78734 267073
rect 78678 266999 78734 267008
rect 77312 266830 77340 266999
rect 78692 266898 78720 266999
rect 78680 266892 78732 266898
rect 78680 266834 78732 266840
rect 77300 266824 77352 266830
rect 77300 266766 77352 266772
rect 62212 266144 62264 266150
rect 62212 266086 62264 266092
rect 62224 264790 62252 266086
rect 62212 264784 62264 264790
rect 62212 264726 62264 264732
rect 79336 250578 79364 268058
rect 83108 268054 83136 269583
rect 91296 269142 91324 269583
rect 91284 269136 91336 269142
rect 91284 269078 91336 269084
rect 90730 268832 90786 268841
rect 90730 268767 90786 268776
rect 90744 268598 90772 268767
rect 93596 268666 93624 269583
rect 94516 268734 94544 269583
rect 110972 269554 111024 269560
rect 133432 269550 133460 269719
rect 133420 269544 133472 269550
rect 133420 269486 133472 269492
rect 135916 269482 135944 269719
rect 135904 269476 135956 269482
rect 135904 269418 135956 269424
rect 138492 269414 138520 269719
rect 138480 269408 138532 269414
rect 138480 269350 138532 269356
rect 140884 269346 140912 269719
rect 148508 269690 148560 269696
rect 143538 269648 143594 269657
rect 143538 269583 143594 269592
rect 145930 269648 145986 269657
rect 145930 269583 145986 269592
rect 140872 269340 140924 269346
rect 140872 269282 140924 269288
rect 143552 269278 143580 269583
rect 143540 269272 143592 269278
rect 143540 269214 143592 269220
rect 145944 269210 145972 269583
rect 145932 269204 145984 269210
rect 145932 269146 145984 269152
rect 196624 269068 196676 269074
rect 196624 269010 196676 269016
rect 95882 268832 95938 268841
rect 95882 268767 95938 268776
rect 96066 268832 96122 268841
rect 96066 268767 96122 268776
rect 98458 268832 98514 268841
rect 98458 268767 98514 268776
rect 99378 268832 99434 268841
rect 99378 268767 99434 268776
rect 100758 268832 100814 268841
rect 100758 268767 100814 268776
rect 106370 268832 106426 268841
rect 106370 268767 106426 268776
rect 94504 268728 94556 268734
rect 94504 268670 94556 268676
rect 93584 268660 93636 268666
rect 93584 268602 93636 268608
rect 90732 268592 90784 268598
rect 90732 268534 90784 268540
rect 95896 268190 95924 268767
rect 96080 268462 96108 268767
rect 98472 268530 98500 268767
rect 98460 268524 98512 268530
rect 98460 268466 98512 268472
rect 96068 268456 96120 268462
rect 96068 268398 96120 268404
rect 95884 268184 95936 268190
rect 85394 268152 85450 268161
rect 85394 268087 85450 268096
rect 92386 268152 92442 268161
rect 95884 268126 95936 268132
rect 92386 268087 92442 268096
rect 83096 268048 83148 268054
rect 83096 267990 83148 267996
rect 84198 267744 84254 267753
rect 84198 267679 84254 267688
rect 80060 266416 80112 266422
rect 80060 266358 80112 266364
rect 80072 264246 80100 266358
rect 84212 266082 84240 267679
rect 84200 266076 84252 266082
rect 84200 266018 84252 266024
rect 85408 265878 85436 268087
rect 88338 267064 88394 267073
rect 88338 266999 88394 267008
rect 88352 266966 88380 266999
rect 88340 266960 88392 266966
rect 88340 266902 88392 266908
rect 85578 266384 85634 266393
rect 85578 266319 85634 266328
rect 86958 266384 87014 266393
rect 86958 266319 87014 266328
rect 88338 266384 88394 266393
rect 88338 266319 88394 266328
rect 89718 266384 89774 266393
rect 92400 266354 92428 268087
rect 96988 267980 97040 267986
rect 96988 267922 97040 267928
rect 97000 267753 97028 267922
rect 99392 267850 99420 268767
rect 100772 268394 100800 268767
rect 100760 268388 100812 268394
rect 100760 268330 100812 268336
rect 103518 268152 103574 268161
rect 106384 268122 106412 268767
rect 113546 268152 113602 268161
rect 103518 268087 103574 268096
rect 106372 268116 106424 268122
rect 102692 267912 102744 267918
rect 102692 267854 102744 267860
rect 99380 267844 99432 267850
rect 99380 267786 99432 267792
rect 98000 267776 98052 267782
rect 96986 267744 97042 267753
rect 96986 267679 97042 267688
rect 97998 267744 98000 267753
rect 102704 267753 102732 267854
rect 98052 267744 98054 267753
rect 97998 267679 98054 267688
rect 102690 267744 102746 267753
rect 102690 267679 102746 267688
rect 103532 267102 103560 268087
rect 113546 268087 113602 268096
rect 128358 268152 128414 268161
rect 128358 268087 128414 268096
rect 106372 268058 106424 268064
rect 106924 267912 106976 267918
rect 106924 267854 106976 267860
rect 104898 267200 104954 267209
rect 104898 267135 104900 267144
rect 104952 267135 104954 267144
rect 104900 267106 104952 267112
rect 103520 267096 103572 267102
rect 100758 267064 100814 267073
rect 103520 267038 103572 267044
rect 100758 266999 100760 267008
rect 100812 266999 100814 267008
rect 100760 266970 100812 266976
rect 104898 266520 104954 266529
rect 104898 266455 104954 266464
rect 104912 266422 104940 266455
rect 104900 266416 104952 266422
rect 92478 266384 92534 266393
rect 89718 266319 89774 266328
rect 92388 266348 92440 266354
rect 85592 265946 85620 266319
rect 85580 265940 85632 265946
rect 85580 265882 85632 265888
rect 85396 265872 85448 265878
rect 85396 265814 85448 265820
rect 86972 265742 87000 266319
rect 88352 265810 88380 266319
rect 89732 266014 89760 266319
rect 104900 266358 104952 266364
rect 106278 266384 106334 266393
rect 92478 266319 92534 266328
rect 106278 266319 106334 266328
rect 92388 266290 92440 266296
rect 92492 266150 92520 266319
rect 92480 266144 92532 266150
rect 92480 266086 92532 266092
rect 89720 266008 89772 266014
rect 89720 265950 89772 265956
rect 88340 265804 88392 265810
rect 88340 265746 88392 265752
rect 86960 265736 87012 265742
rect 86960 265678 87012 265684
rect 88248 265736 88300 265742
rect 88248 265678 88300 265684
rect 88260 264926 88288 265678
rect 88248 264920 88300 264926
rect 88248 264862 88300 264868
rect 80060 264240 80112 264246
rect 80060 264182 80112 264188
rect 79324 250572 79376 250578
rect 79324 250514 79376 250520
rect 85856 250572 85908 250578
rect 85856 250514 85908 250520
rect 85868 249121 85896 250514
rect 106292 250510 106320 266319
rect 106936 250578 106964 267854
rect 112352 267844 112404 267850
rect 112352 267786 112404 267792
rect 111248 267776 111300 267782
rect 111246 267744 111248 267753
rect 112364 267753 112392 267786
rect 111300 267744 111302 267753
rect 111246 267679 111302 267688
rect 112350 267744 112406 267753
rect 112350 267679 112406 267688
rect 107658 267336 107714 267345
rect 113560 267306 113588 268087
rect 119068 267912 119120 267918
rect 119068 267854 119120 267860
rect 119080 267753 119108 267854
rect 119066 267744 119122 267753
rect 119066 267679 119122 267688
rect 120078 267744 120134 267753
rect 120078 267679 120134 267688
rect 125598 267744 125654 267753
rect 128372 267714 128400 268087
rect 196636 267782 196664 269010
rect 196624 267776 196676 267782
rect 150990 267744 151046 267753
rect 125598 267679 125654 267688
rect 128360 267708 128412 267714
rect 120092 267578 120120 267679
rect 125612 267646 125640 267679
rect 150990 267679 151046 267688
rect 158534 267744 158590 267753
rect 158534 267679 158536 267688
rect 128360 267650 128412 267656
rect 151004 267646 151032 267679
rect 158588 267679 158590 267688
rect 163502 267744 163558 267753
rect 196912 267734 196940 465695
rect 197004 370462 197032 477498
rect 197360 471300 197412 471306
rect 197360 471242 197412 471248
rect 197084 465996 197136 466002
rect 197084 465938 197136 465944
rect 197096 374134 197124 465938
rect 197176 375352 197228 375358
rect 197176 375294 197228 375300
rect 197084 374128 197136 374134
rect 197084 374070 197136 374076
rect 196992 370456 197044 370462
rect 196992 370398 197044 370404
rect 197188 269074 197216 375294
rect 197372 371074 197400 471242
rect 197556 466454 197584 480037
rect 197648 480023 198030 480051
rect 197648 471306 197676 480023
rect 197728 478984 197780 478990
rect 197728 478926 197780 478932
rect 197636 471300 197688 471306
rect 197636 471242 197688 471248
rect 197464 466426 197584 466454
rect 197360 371068 197412 371074
rect 197360 371010 197412 371016
rect 197464 370870 197492 466426
rect 197544 459060 197596 459066
rect 197544 459002 197596 459008
rect 197452 370864 197504 370870
rect 197452 370806 197504 370812
rect 197360 355224 197412 355230
rect 197360 355166 197412 355172
rect 197176 269068 197228 269074
rect 197176 269010 197228 269016
rect 196624 267718 196676 267724
rect 163502 267679 163558 267688
rect 158536 267650 158588 267656
rect 125600 267640 125652 267646
rect 150992 267640 151044 267646
rect 125600 267582 125652 267588
rect 129738 267608 129794 267617
rect 120080 267572 120132 267578
rect 150992 267582 151044 267588
rect 155958 267608 156014 267617
rect 129738 267543 129794 267552
rect 155958 267543 156014 267552
rect 160926 267608 160982 267617
rect 160926 267543 160982 267552
rect 120080 267514 120132 267520
rect 129752 267510 129780 267543
rect 129740 267504 129792 267510
rect 115938 267472 115994 267481
rect 115938 267407 115994 267416
rect 117318 267472 117374 267481
rect 129740 267446 129792 267452
rect 155972 267442 156000 267543
rect 117318 267407 117320 267416
rect 115952 267374 115980 267407
rect 117372 267407 117374 267416
rect 155960 267436 156012 267442
rect 117320 267378 117372 267384
rect 155960 267378 156012 267384
rect 160940 267374 160968 267543
rect 163516 267510 163544 267679
rect 163504 267504 163556 267510
rect 163504 267446 163556 267452
rect 115940 267368 115992 267374
rect 115940 267310 115992 267316
rect 160928 267368 160980 267374
rect 160928 267310 160980 267316
rect 183282 267336 183338 267345
rect 107658 267271 107714 267280
rect 113548 267300 113600 267306
rect 107672 267238 107700 267271
rect 183282 267271 183338 267280
rect 113548 267242 113600 267248
rect 107660 267232 107712 267238
rect 107660 267174 107712 267180
rect 109958 267064 110014 267073
rect 183296 267034 183324 267271
rect 183466 267064 183522 267073
rect 109958 266999 110014 267008
rect 183284 267028 183336 267034
rect 107658 266384 107714 266393
rect 109972 266354 110000 266999
rect 183466 266999 183522 267008
rect 183284 266970 183336 266976
rect 114374 266656 114430 266665
rect 114374 266591 114430 266600
rect 117318 266656 117374 266665
rect 117318 266591 117374 266600
rect 113730 266384 113786 266393
rect 107658 266319 107714 266328
rect 109960 266348 110012 266354
rect 107672 265674 107700 266319
rect 113730 266319 113786 266328
rect 109960 266290 110012 266296
rect 113744 265742 113772 266319
rect 113732 265736 113784 265742
rect 113732 265678 113784 265684
rect 114388 265674 114416 266591
rect 117332 266286 117360 266591
rect 183480 266422 183508 266999
rect 183468 266416 183520 266422
rect 183468 266358 183520 266364
rect 117320 266280 117372 266286
rect 117320 266222 117372 266228
rect 107660 265668 107712 265674
rect 107660 265610 107712 265616
rect 114376 265668 114428 265674
rect 114376 265610 114428 265616
rect 106924 250572 106976 250578
rect 106924 250514 106976 250520
rect 179788 250572 179840 250578
rect 179788 250514 179840 250520
rect 106280 250504 106332 250510
rect 106280 250446 106332 250452
rect 179328 250504 179380 250510
rect 179328 250446 179380 250452
rect 179340 249937 179368 250446
rect 179800 249937 179828 250514
rect 179326 249928 179382 249937
rect 179326 249863 179382 249872
rect 179786 249928 179842 249937
rect 179786 249863 179842 249872
rect 190918 249928 190974 249937
rect 190918 249863 190974 249872
rect 190932 249830 190960 249863
rect 190920 249824 190972 249830
rect 190920 249766 190972 249772
rect 85854 249112 85910 249121
rect 85854 249047 85910 249056
rect 62120 249008 62172 249014
rect 62120 248950 62172 248956
rect 96066 164928 96122 164937
rect 96066 164863 96122 164872
rect 115754 164928 115810 164937
rect 115754 164863 115810 164872
rect 96080 164694 96108 164863
rect 96068 164688 96120 164694
rect 84106 164656 84162 164665
rect 96068 164630 96120 164636
rect 103518 164656 103574 164665
rect 84106 164591 84162 164600
rect 103518 164591 103574 164600
rect 105910 164656 105966 164665
rect 105910 164591 105966 164600
rect 114374 164656 114430 164665
rect 115768 164626 115796 164863
rect 138478 164792 138534 164801
rect 138478 164727 138534 164736
rect 140870 164792 140926 164801
rect 140870 164727 140926 164736
rect 143538 164792 143594 164801
rect 143538 164727 143594 164736
rect 163318 164792 163374 164801
rect 163318 164727 163374 164736
rect 118054 164656 118110 164665
rect 114374 164591 114430 164600
rect 115756 164620 115808 164626
rect 60004 163532 60056 163538
rect 60004 163474 60056 163480
rect 76010 162752 76066 162761
rect 76010 162687 76066 162696
rect 77298 162752 77354 162761
rect 77298 162687 77354 162696
rect 78678 162752 78734 162761
rect 78678 162687 78734 162696
rect 80058 162752 80114 162761
rect 80058 162687 80114 162696
rect 81438 162752 81494 162761
rect 81438 162687 81494 162696
rect 82818 162752 82874 162761
rect 82818 162687 82874 162696
rect 75918 162208 75974 162217
rect 75918 162143 75974 162152
rect 60004 160812 60056 160818
rect 60004 160754 60056 160760
rect 60016 160614 60044 160754
rect 60004 160608 60056 160614
rect 60004 160550 60056 160556
rect 59820 146260 59872 146266
rect 59820 146202 59872 146208
rect 59452 146124 59504 146130
rect 59740 146118 59952 146146
rect 59452 146066 59504 146072
rect 59464 145314 59492 146066
rect 59820 145580 59872 145586
rect 59820 145522 59872 145528
rect 59452 145308 59504 145314
rect 59452 145250 59504 145256
rect 59358 140856 59414 140865
rect 59358 140791 59414 140800
rect 59832 59294 59860 145522
rect 59820 59288 59872 59294
rect 59820 59230 59872 59236
rect 59268 57316 59320 57322
rect 59268 57258 59320 57264
rect 59924 56438 59952 146118
rect 59912 56432 59964 56438
rect 59912 56374 59964 56380
rect 59176 56364 59228 56370
rect 59176 56306 59228 56312
rect 60016 56302 60044 160550
rect 75932 145450 75960 162143
rect 75920 145444 75972 145450
rect 75920 145386 75972 145392
rect 76024 145382 76052 162687
rect 77312 145518 77340 162687
rect 78692 148714 78720 162687
rect 78680 148708 78732 148714
rect 78680 148650 78732 148656
rect 80072 148646 80100 162687
rect 80060 148640 80112 148646
rect 80060 148582 80112 148588
rect 81452 148578 81480 162687
rect 81440 148572 81492 148578
rect 81440 148514 81492 148520
rect 82832 145790 82860 162687
rect 84120 161673 84148 164591
rect 98458 164248 98514 164257
rect 98458 164183 98514 164192
rect 101034 164248 101090 164257
rect 101034 164183 101090 164192
rect 98472 164014 98500 164183
rect 101048 164082 101076 164183
rect 101036 164076 101088 164082
rect 101036 164018 101088 164024
rect 98460 164008 98512 164014
rect 98460 163950 98512 163956
rect 103532 163946 103560 164591
rect 103520 163940 103572 163946
rect 103520 163882 103572 163888
rect 105924 163878 105952 164591
rect 108210 164248 108266 164257
rect 108210 164183 108266 164192
rect 105912 163872 105964 163878
rect 105912 163814 105964 163820
rect 108224 163742 108252 164183
rect 111154 163976 111210 163985
rect 111154 163911 111210 163920
rect 111168 163878 111196 163911
rect 110788 163872 110840 163878
rect 110788 163814 110840 163820
rect 111156 163872 111208 163878
rect 111156 163814 111208 163820
rect 108212 163736 108264 163742
rect 108212 163678 108264 163684
rect 110512 163736 110564 163742
rect 110512 163678 110564 163684
rect 99378 163160 99434 163169
rect 99378 163095 99434 163104
rect 84198 162752 84254 162761
rect 84198 162687 84254 162696
rect 85578 162752 85634 162761
rect 85578 162687 85634 162696
rect 86958 162752 87014 162761
rect 86958 162687 87014 162696
rect 88430 162752 88486 162761
rect 88430 162687 88486 162696
rect 89810 162752 89866 162761
rect 89810 162687 89866 162696
rect 90730 162752 90786 162761
rect 90730 162687 90786 162696
rect 91190 162752 91246 162761
rect 91190 162687 91246 162696
rect 92478 162752 92534 162761
rect 92478 162687 92534 162696
rect 93858 162752 93914 162761
rect 93858 162687 93914 162696
rect 95238 162752 95294 162761
rect 95238 162687 95294 162696
rect 96618 162752 96674 162761
rect 96618 162687 96674 162696
rect 97998 162752 98054 162761
rect 97998 162687 98054 162696
rect 84106 161664 84162 161673
rect 84106 161599 84162 161608
rect 84212 145858 84240 162687
rect 84290 161664 84346 161673
rect 84290 161599 84346 161608
rect 84304 145926 84332 161599
rect 85592 145994 85620 162687
rect 86972 146198 87000 162687
rect 88338 162208 88394 162217
rect 88338 162143 88394 162152
rect 88352 161974 88380 162143
rect 88340 161968 88392 161974
rect 88340 161910 88392 161916
rect 86960 146192 87012 146198
rect 86960 146134 87012 146140
rect 88444 146130 88472 162687
rect 88432 146124 88484 146130
rect 88432 146066 88484 146072
rect 89824 146062 89852 162687
rect 90744 162042 90772 162687
rect 90914 162480 90970 162489
rect 90914 162415 90970 162424
rect 91098 162480 91154 162489
rect 91098 162415 91154 162424
rect 90928 162217 90956 162415
rect 90914 162208 90970 162217
rect 90914 162143 90970 162152
rect 90732 162036 90784 162042
rect 90732 161978 90784 161984
rect 89812 146056 89864 146062
rect 89812 145998 89864 146004
rect 85580 145988 85632 145994
rect 85580 145930 85632 145936
rect 84292 145920 84344 145926
rect 84292 145862 84344 145868
rect 84200 145852 84252 145858
rect 84200 145794 84252 145800
rect 82820 145784 82872 145790
rect 82820 145726 82872 145732
rect 91112 145654 91140 162415
rect 91204 145722 91232 162687
rect 92492 146033 92520 162687
rect 92478 146024 92534 146033
rect 92478 145959 92534 145968
rect 91192 145716 91244 145722
rect 91192 145658 91244 145664
rect 91100 145648 91152 145654
rect 91100 145590 91152 145596
rect 93872 145586 93900 162687
rect 95252 161022 95280 162687
rect 95240 161016 95292 161022
rect 95240 160958 95292 160964
rect 96632 160954 96660 162687
rect 96620 160948 96672 160954
rect 96620 160890 96672 160896
rect 98012 160886 98040 162687
rect 98644 161492 98696 161498
rect 98644 161434 98696 161440
rect 98000 160880 98052 160886
rect 98000 160822 98052 160828
rect 98656 145897 98684 161434
rect 99392 161294 99420 163095
rect 110524 162761 110552 163678
rect 100758 162752 100814 162761
rect 100758 162687 100814 162696
rect 102138 162752 102194 162761
rect 102138 162687 102194 162696
rect 103794 162752 103850 162761
rect 103794 162687 103850 162696
rect 104898 162752 104954 162761
rect 104898 162687 104954 162696
rect 106278 162752 106334 162761
rect 106278 162687 106334 162696
rect 107658 162752 107714 162761
rect 107658 162687 107714 162696
rect 110510 162752 110566 162761
rect 110510 162687 110566 162696
rect 100772 162178 100800 162687
rect 100024 162172 100076 162178
rect 100024 162114 100076 162120
rect 100760 162172 100812 162178
rect 100760 162114 100812 162120
rect 99380 161288 99432 161294
rect 99380 161230 99432 161236
rect 98642 145888 98698 145897
rect 98642 145823 98698 145832
rect 100036 145761 100064 162114
rect 100758 162072 100814 162081
rect 100758 162007 100814 162016
rect 100022 145752 100078 145761
rect 100022 145687 100078 145696
rect 100772 145625 100800 162007
rect 102152 146266 102180 162687
rect 103808 161498 103836 162687
rect 103796 161492 103848 161498
rect 103796 161434 103848 161440
rect 104912 147558 104940 162687
rect 106292 160818 106320 162687
rect 106370 162480 106426 162489
rect 106370 162415 106426 162424
rect 106384 161362 106412 162415
rect 106372 161356 106424 161362
rect 106372 161298 106424 161304
rect 106280 160812 106332 160818
rect 106280 160754 106332 160760
rect 107672 147626 107700 162687
rect 110524 148374 110552 162687
rect 110800 148510 110828 163814
rect 113454 163704 113510 163713
rect 113454 163639 113510 163648
rect 113468 163062 113496 163639
rect 113456 163056 113508 163062
rect 113456 162998 113508 163004
rect 114388 162994 114416 164591
rect 118054 164591 118110 164600
rect 115756 164562 115808 164568
rect 114376 162988 114428 162994
rect 114376 162930 114428 162936
rect 118068 162926 118096 164591
rect 138492 164490 138520 164727
rect 140884 164558 140912 164727
rect 140872 164552 140924 164558
rect 140872 164494 140924 164500
rect 138480 164484 138532 164490
rect 138480 164426 138532 164432
rect 143552 164422 143580 164727
rect 153382 164656 153438 164665
rect 153382 164591 153438 164600
rect 143540 164416 143592 164422
rect 143540 164358 143592 164364
rect 122746 164248 122802 164257
rect 122746 164183 122802 164192
rect 145930 164248 145986 164257
rect 145930 164183 145986 164192
rect 148506 164248 148562 164257
rect 148506 164183 148562 164192
rect 150898 164248 150954 164257
rect 150898 164183 150954 164192
rect 118056 162920 118108 162926
rect 118056 162862 118108 162868
rect 110970 162752 111026 162761
rect 110970 162687 111026 162696
rect 113178 162752 113234 162761
rect 113178 162687 113234 162696
rect 115938 162752 115994 162761
rect 115938 162687 115994 162696
rect 118330 162752 118386 162761
rect 118330 162687 118386 162696
rect 118698 162752 118754 162761
rect 118698 162687 118754 162696
rect 120722 162752 120778 162761
rect 120722 162687 120778 162696
rect 110984 162110 111012 162687
rect 112810 162208 112866 162217
rect 112810 162143 112812 162152
rect 112864 162143 112866 162152
rect 113088 162172 113140 162178
rect 112812 162114 112864 162120
rect 113088 162114 113140 162120
rect 110972 162104 111024 162110
rect 110972 162046 111024 162052
rect 113100 161514 113128 162114
rect 113192 161906 113220 162687
rect 113180 161900 113232 161906
rect 113180 161842 113232 161848
rect 113100 161486 113220 161514
rect 110788 148504 110840 148510
rect 110788 148446 110840 148452
rect 113192 148442 113220 161486
rect 115952 161430 115980 162687
rect 116030 162480 116086 162489
rect 116030 162415 116086 162424
rect 116044 162314 116072 162415
rect 116032 162308 116084 162314
rect 116032 162250 116084 162256
rect 118344 162246 118372 162687
rect 118332 162240 118384 162246
rect 118332 162182 118384 162188
rect 115940 161424 115992 161430
rect 115940 161366 115992 161372
rect 118712 160750 118740 162687
rect 120736 162382 120764 162687
rect 122760 162518 122788 164183
rect 145944 163810 145972 164183
rect 145932 163804 145984 163810
rect 145932 163746 145984 163752
rect 148520 163674 148548 164183
rect 148508 163668 148560 163674
rect 148508 163610 148560 163616
rect 150912 163606 150940 164183
rect 150900 163600 150952 163606
rect 150900 163542 150952 163548
rect 153396 163538 153424 164591
rect 163332 164354 163360 164727
rect 165894 164656 165950 164665
rect 165894 164591 165950 164600
rect 163320 164348 163372 164354
rect 163320 164290 163372 164296
rect 165908 164286 165936 164591
rect 165896 164280 165948 164286
rect 165896 164222 165948 164228
rect 196636 163878 196664 267718
rect 196820 267706 196940 267734
rect 196820 266354 196848 267706
rect 196808 266348 196860 266354
rect 196808 266290 196860 266296
rect 196716 266008 196768 266014
rect 196716 265950 196768 265956
rect 196728 265674 196756 265950
rect 196716 265668 196768 265674
rect 196716 265610 196768 265616
rect 196624 163872 196676 163878
rect 196624 163814 196676 163820
rect 153384 163532 153436 163538
rect 153384 163474 153436 163480
rect 128358 163160 128414 163169
rect 128358 163095 128414 163104
rect 123024 163056 123076 163062
rect 123024 162998 123076 163004
rect 123036 162518 123064 162998
rect 125874 162752 125930 162761
rect 125874 162687 125930 162696
rect 122748 162512 122800 162518
rect 122748 162454 122800 162460
rect 123024 162512 123076 162518
rect 123024 162454 123076 162460
rect 125888 162450 125916 162687
rect 128372 162586 128400 163095
rect 155960 162852 156012 162858
rect 155960 162794 156012 162800
rect 135996 162784 136048 162790
rect 130842 162752 130898 162761
rect 130842 162687 130898 162696
rect 133418 162752 133474 162761
rect 133418 162687 133420 162696
rect 130856 162654 130884 162687
rect 133472 162687 133474 162696
rect 135994 162752 135996 162761
rect 155972 162761 156000 162794
rect 136048 162752 136050 162761
rect 135994 162687 136050 162696
rect 155958 162752 156014 162761
rect 155958 162687 156014 162696
rect 183466 162752 183522 162761
rect 183466 162687 183522 162696
rect 133420 162658 133472 162664
rect 130844 162648 130896 162654
rect 130844 162590 130896 162596
rect 183190 162616 183246 162625
rect 128360 162580 128412 162586
rect 183190 162551 183246 162560
rect 128360 162522 128412 162528
rect 125876 162444 125928 162450
rect 125876 162386 125928 162392
rect 120724 162376 120776 162382
rect 120724 162318 120776 162324
rect 183204 162246 183232 162551
rect 183480 162382 183508 162687
rect 196728 162518 196756 265610
rect 196820 163742 196848 266290
rect 197372 251122 197400 355166
rect 197452 266416 197504 266422
rect 197452 266358 197504 266364
rect 197360 251116 197412 251122
rect 197360 251058 197412 251064
rect 197464 171134 197492 266358
rect 197556 266014 197584 459002
rect 197636 458856 197688 458862
rect 197636 458798 197688 458804
rect 197648 267510 197676 458798
rect 197740 373250 197768 478926
rect 198476 478174 198504 480037
rect 198858 480023 198964 480051
rect 198464 478168 198516 478174
rect 198464 478110 198516 478116
rect 198004 478032 198056 478038
rect 198004 477974 198056 477980
rect 197820 475516 197872 475522
rect 197820 475458 197872 475464
rect 197832 373590 197860 475458
rect 197820 373584 197872 373590
rect 197820 373526 197872 373532
rect 197728 373244 197780 373250
rect 197728 373186 197780 373192
rect 197728 354748 197780 354754
rect 197728 354690 197780 354696
rect 197636 267504 197688 267510
rect 197636 267446 197688 267452
rect 197544 266008 197596 266014
rect 197544 265950 197596 265956
rect 197740 258074 197768 354690
rect 198016 268394 198044 477974
rect 198096 475720 198148 475726
rect 198096 475662 198148 475668
rect 198108 410582 198136 475662
rect 198188 475244 198240 475250
rect 198188 475186 198240 475192
rect 198096 410576 198148 410582
rect 198096 410518 198148 410524
rect 198094 394632 198150 394641
rect 198094 394567 198150 394576
rect 198004 268388 198056 268394
rect 198004 268330 198056 268336
rect 197912 267844 197964 267850
rect 197912 267786 197964 267792
rect 197924 258074 197952 267786
rect 198108 267646 198136 394567
rect 198200 393446 198228 475186
rect 198936 471510 198964 480023
rect 199028 480023 199318 480051
rect 199488 480023 199778 480051
rect 198924 471504 198976 471510
rect 198924 471446 198976 471452
rect 198740 471300 198792 471306
rect 198740 471242 198792 471248
rect 198280 461644 198332 461650
rect 198280 461586 198332 461592
rect 198188 393440 198240 393446
rect 198188 393382 198240 393388
rect 198292 392057 198320 461586
rect 198372 393372 198424 393378
rect 198372 393314 198424 393320
rect 198278 392048 198334 392057
rect 198278 391983 198334 391992
rect 198186 390688 198242 390697
rect 198186 390623 198242 390632
rect 198200 375358 198228 390623
rect 198188 375352 198240 375358
rect 198188 375294 198240 375300
rect 198384 373182 198412 393314
rect 198372 373176 198424 373182
rect 198372 373118 198424 373124
rect 198752 370394 198780 471242
rect 199028 468466 199056 480023
rect 199384 477624 199436 477630
rect 199384 477566 199436 477572
rect 199108 471504 199160 471510
rect 199108 471446 199160 471452
rect 198844 468438 199056 468466
rect 198844 371142 198872 468438
rect 199120 463694 199148 471446
rect 199200 471232 199252 471238
rect 199200 471174 199252 471180
rect 198936 463666 199148 463694
rect 198832 371136 198884 371142
rect 198832 371078 198884 371084
rect 198936 370938 198964 463666
rect 199016 460216 199068 460222
rect 199016 460158 199068 460164
rect 199028 458386 199056 460158
rect 199108 458992 199160 458998
rect 199108 458934 199160 458940
rect 199016 458380 199068 458386
rect 199016 458322 199068 458328
rect 199028 454753 199056 458322
rect 199014 454744 199070 454753
rect 199014 454679 199070 454688
rect 198924 370932 198976 370938
rect 198924 370874 198976 370880
rect 198740 370388 198792 370394
rect 198740 370330 198792 370336
rect 199028 349625 199056 454679
rect 199120 373658 199148 458934
rect 199212 390833 199240 471174
rect 199292 410576 199344 410582
rect 199292 410518 199344 410524
rect 199198 390824 199254 390833
rect 199198 390759 199254 390768
rect 199304 373726 199332 410518
rect 199292 373720 199344 373726
rect 199292 373662 199344 373668
rect 199108 373652 199160 373658
rect 199108 373594 199160 373600
rect 199396 370598 199424 477566
rect 199488 471306 199516 480023
rect 200224 478310 200252 480037
rect 200316 480023 200698 480051
rect 200776 480023 201066 480051
rect 201526 480023 201632 480051
rect 200120 478304 200172 478310
rect 200118 478272 200120 478281
rect 200212 478304 200264 478310
rect 200172 478272 200174 478281
rect 200212 478246 200264 478252
rect 200118 478207 200174 478216
rect 200316 476114 200344 480023
rect 200672 478440 200724 478446
rect 200672 478382 200724 478388
rect 200684 477737 200712 478382
rect 200670 477728 200726 477737
rect 200670 477663 200726 477672
rect 200224 476086 200344 476114
rect 199660 475448 199712 475454
rect 199660 475390 199712 475396
rect 199476 471300 199528 471306
rect 199476 471242 199528 471248
rect 199568 465656 199620 465662
rect 199568 465598 199620 465604
rect 199476 459672 199528 459678
rect 199476 459614 199528 459620
rect 199488 374134 199516 459614
rect 199580 391270 199608 465598
rect 199672 411942 199700 475390
rect 199660 411936 199712 411942
rect 199660 411878 199712 411884
rect 199658 394088 199714 394097
rect 199658 394023 199714 394032
rect 199672 393990 199700 394023
rect 199660 393984 199712 393990
rect 199660 393926 199712 393932
rect 199568 391264 199620 391270
rect 199568 391206 199620 391212
rect 199566 390824 199622 390833
rect 199566 390759 199622 390768
rect 199476 374128 199528 374134
rect 199476 374070 199528 374076
rect 199474 372736 199530 372745
rect 199474 372671 199530 372680
rect 199384 370592 199436 370598
rect 199384 370534 199436 370540
rect 199384 366376 199436 366382
rect 199384 366318 199436 366324
rect 198738 349616 198794 349625
rect 198738 349551 198794 349560
rect 199014 349616 199070 349625
rect 199014 349551 199070 349560
rect 198096 267640 198148 267646
rect 198096 267582 198148 267588
rect 198280 267096 198332 267102
rect 198280 267038 198332 267044
rect 198292 266422 198320 267038
rect 198280 266416 198332 266422
rect 198280 266358 198332 266364
rect 197556 258046 197768 258074
rect 197832 258046 197952 258074
rect 197556 250510 197584 258046
rect 197636 251116 197688 251122
rect 197636 251058 197688 251064
rect 197648 250578 197676 251058
rect 197636 250572 197688 250578
rect 197636 250514 197688 250520
rect 197544 250504 197596 250510
rect 197544 250446 197596 250452
rect 197372 171106 197492 171134
rect 196808 163736 196860 163742
rect 196808 163678 196860 163684
rect 196716 162512 196768 162518
rect 196716 162454 196768 162460
rect 197372 162382 197400 171106
rect 197452 162920 197504 162926
rect 197452 162862 197504 162868
rect 183468 162376 183520 162382
rect 183468 162318 183520 162324
rect 197360 162376 197412 162382
rect 197360 162318 197412 162324
rect 183192 162240 183244 162246
rect 183192 162182 183244 162188
rect 118700 160744 118752 160750
rect 118700 160686 118752 160692
rect 113180 148436 113232 148442
rect 113180 148378 113232 148384
rect 110512 148368 110564 148374
rect 110512 148310 110564 148316
rect 107660 147620 107712 147626
rect 107660 147562 107712 147568
rect 104900 147552 104952 147558
rect 104900 147494 104952 147500
rect 102140 146260 102192 146266
rect 102140 146202 102192 146208
rect 179052 146260 179104 146266
rect 179052 146202 179104 146208
rect 100758 145616 100814 145625
rect 93860 145580 93912 145586
rect 100758 145551 100814 145560
rect 93860 145522 93912 145528
rect 77300 145512 77352 145518
rect 77300 145454 77352 145460
rect 76012 145376 76064 145382
rect 76012 145318 76064 145324
rect 179064 144945 179092 146202
rect 179696 146192 179748 146198
rect 179696 146134 179748 146140
rect 179708 144945 179736 146134
rect 191748 145580 191800 145586
rect 191748 145522 191800 145528
rect 191760 145489 191788 145522
rect 191746 145480 191802 145489
rect 191746 145415 191802 145424
rect 179050 144936 179106 144945
rect 179050 144871 179106 144880
rect 179694 144936 179750 144945
rect 179694 144871 179750 144880
rect 77114 59800 77170 59809
rect 77114 59735 77170 59744
rect 83094 59800 83150 59809
rect 83094 59735 83150 59744
rect 99470 59800 99526 59809
rect 99470 59735 99526 59744
rect 113546 59800 113602 59809
rect 113546 59735 113602 59744
rect 77128 59634 77156 59735
rect 77116 59628 77168 59634
rect 77116 59570 77168 59576
rect 83108 59566 83136 59735
rect 94502 59664 94558 59673
rect 94502 59599 94558 59608
rect 95698 59664 95754 59673
rect 95698 59599 95754 59608
rect 83096 59560 83148 59566
rect 83096 59502 83148 59508
rect 84200 59356 84252 59362
rect 84200 59298 84252 59304
rect 84212 58041 84240 59298
rect 94516 59294 94544 59599
rect 95712 59401 95740 59599
rect 99484 59498 99512 59735
rect 102782 59664 102838 59673
rect 102782 59599 102838 59608
rect 103886 59664 103942 59673
rect 103886 59599 103942 59608
rect 99472 59492 99524 59498
rect 99472 59434 99524 59440
rect 95698 59392 95754 59401
rect 95698 59327 95754 59336
rect 95882 59392 95938 59401
rect 95882 59327 95938 59336
rect 96986 59392 97042 59401
rect 96986 59327 97042 59336
rect 101770 59392 101826 59401
rect 101770 59327 101826 59336
rect 94504 59288 94556 59294
rect 94504 59230 94556 59236
rect 95896 59226 95924 59327
rect 95884 59220 95936 59226
rect 95884 59162 95936 59168
rect 97000 59158 97028 59327
rect 96988 59152 97040 59158
rect 96988 59094 97040 59100
rect 101784 59022 101812 59327
rect 102796 59090 102824 59599
rect 102784 59084 102836 59090
rect 102784 59026 102836 59032
rect 101772 59016 101824 59022
rect 101772 58958 101824 58964
rect 103900 58954 103928 59599
rect 113560 59430 113588 59735
rect 113548 59424 113600 59430
rect 111154 59392 111210 59401
rect 113548 59366 113600 59372
rect 115938 59392 115994 59401
rect 111154 59327 111210 59336
rect 115938 59327 115994 59336
rect 103888 58948 103940 58954
rect 103888 58890 103940 58896
rect 111168 58886 111196 59327
rect 111156 58880 111208 58886
rect 111156 58822 111208 58828
rect 115952 58818 115980 59327
rect 148506 59256 148562 59265
rect 148506 59191 148562 59200
rect 150898 59256 150954 59265
rect 150898 59191 150954 59200
rect 115940 58812 115992 58818
rect 115940 58754 115992 58760
rect 148520 58750 148548 59191
rect 148508 58744 148560 58750
rect 148508 58686 148560 58692
rect 150912 58682 150940 59191
rect 150900 58676 150952 58682
rect 150900 58618 150952 58624
rect 84198 58032 84254 58041
rect 84198 57967 84254 57976
rect 76010 57896 76066 57905
rect 76010 57831 76066 57840
rect 78218 57896 78274 57905
rect 78218 57831 78274 57840
rect 79506 57896 79562 57905
rect 79506 57831 79562 57840
rect 80058 57896 80114 57905
rect 80058 57831 80114 57840
rect 81806 57896 81862 57905
rect 81806 57831 81862 57840
rect 85394 57896 85450 57905
rect 85394 57831 85450 57840
rect 86498 57896 86554 57905
rect 86498 57831 86554 57840
rect 86958 57896 87014 57905
rect 86958 57831 87014 57840
rect 88338 57896 88394 57905
rect 88338 57831 88394 57840
rect 88706 57896 88762 57905
rect 88706 57831 88762 57840
rect 89718 57896 89774 57905
rect 89718 57831 89774 57840
rect 90730 57896 90786 57905
rect 90730 57831 90786 57840
rect 91190 57896 91246 57905
rect 91190 57831 91246 57840
rect 92110 57896 92166 57905
rect 92110 57831 92166 57840
rect 92478 57896 92534 57905
rect 92478 57831 92534 57840
rect 93674 57896 93730 57905
rect 93674 57831 93730 57840
rect 98090 57896 98146 57905
rect 98090 57831 98146 57840
rect 106370 57896 106426 57905
rect 106370 57831 106426 57840
rect 107382 57896 107438 57905
rect 107382 57831 107438 57840
rect 108026 57896 108082 57905
rect 108026 57831 108082 57840
rect 112074 57896 112130 57905
rect 112074 57831 112130 57840
rect 113178 57896 113234 57905
rect 113178 57831 113234 57840
rect 123482 57896 123538 57905
rect 123482 57831 123538 57840
rect 130842 57896 130898 57905
rect 130842 57831 130898 57840
rect 133234 57896 133290 57905
rect 133234 57831 133290 57840
rect 145562 57896 145618 57905
rect 145562 57831 145564 57840
rect 76024 57186 76052 57831
rect 78232 57254 78260 57831
rect 78220 57248 78272 57254
rect 78220 57190 78272 57196
rect 76012 57180 76064 57186
rect 76012 57122 76064 57128
rect 60004 56296 60056 56302
rect 60004 56238 60056 56244
rect 79520 55962 79548 57831
rect 79508 55956 79560 55962
rect 79508 55898 79560 55904
rect 58992 54732 59044 54738
rect 58992 54674 59044 54680
rect 80072 54670 80100 57831
rect 81820 56030 81848 57831
rect 85408 56574 85436 57831
rect 85396 56568 85448 56574
rect 85396 56510 85448 56516
rect 86512 56098 86540 57831
rect 86500 56092 86552 56098
rect 86500 56034 86552 56040
rect 81808 56024 81860 56030
rect 81808 55966 81860 55972
rect 86972 54942 87000 57831
rect 88352 57390 88380 57831
rect 88340 57384 88392 57390
rect 88340 57326 88392 57332
rect 88720 56166 88748 57831
rect 88708 56160 88760 56166
rect 88708 56102 88760 56108
rect 86960 54936 87012 54942
rect 86960 54878 87012 54884
rect 89732 54806 89760 57831
rect 90744 57526 90772 57831
rect 90732 57520 90784 57526
rect 90732 57462 90784 57468
rect 89720 54800 89772 54806
rect 89720 54742 89772 54748
rect 91204 54738 91232 57831
rect 92124 56234 92152 57831
rect 92112 56228 92164 56234
rect 92112 56170 92164 56176
rect 92492 54874 92520 57831
rect 93688 57322 93716 57831
rect 98104 57458 98132 57831
rect 98642 57488 98698 57497
rect 98092 57452 98144 57458
rect 98642 57423 98698 57432
rect 98092 57394 98144 57400
rect 93676 57316 93728 57322
rect 93676 57258 93728 57264
rect 98656 57089 98684 57423
rect 98642 57080 98698 57089
rect 98642 57015 98698 57024
rect 106384 56302 106412 57831
rect 107396 56370 107424 57831
rect 108040 56438 108068 57831
rect 109038 57624 109094 57633
rect 112088 57594 112116 57831
rect 109038 57559 109094 57568
rect 112076 57588 112128 57594
rect 108028 56432 108080 56438
rect 108028 56374 108080 56380
rect 107384 56364 107436 56370
rect 107384 56306 107436 56312
rect 106372 56296 106424 56302
rect 106372 56238 106424 56244
rect 109052 55010 109080 57559
rect 112076 57530 112128 57536
rect 113192 56506 113220 57831
rect 123496 57798 123524 57831
rect 123484 57792 123536 57798
rect 123484 57734 123536 57740
rect 130856 57730 130884 57831
rect 130844 57724 130896 57730
rect 130844 57666 130896 57672
rect 133248 57662 133276 57831
rect 145616 57831 145618 57840
rect 153290 57896 153346 57905
rect 153290 57831 153346 57840
rect 157430 57896 157486 57905
rect 157430 57831 157486 57840
rect 183282 57896 183338 57905
rect 183282 57831 183284 57840
rect 145564 57802 145616 57808
rect 133236 57656 133288 57662
rect 113270 57624 113326 57633
rect 113270 57559 113326 57568
rect 114558 57624 114614 57633
rect 114558 57559 114614 57568
rect 116122 57624 116178 57633
rect 116122 57559 116178 57568
rect 117318 57624 117374 57633
rect 117318 57559 117374 57568
rect 118698 57624 118754 57633
rect 133236 57598 133288 57604
rect 118698 57559 118754 57568
rect 113180 56500 113232 56506
rect 113180 56442 113232 56448
rect 113284 55146 113312 57559
rect 113272 55140 113324 55146
rect 113272 55082 113324 55088
rect 114572 55078 114600 57559
rect 114560 55072 114612 55078
rect 114560 55014 114612 55020
rect 109040 55004 109092 55010
rect 109040 54946 109092 54952
rect 92480 54868 92532 54874
rect 92480 54810 92532 54816
rect 91192 54732 91244 54738
rect 91192 54674 91244 54680
rect 80060 54664 80112 54670
rect 116136 54641 116164 57559
rect 117332 55214 117360 57559
rect 117320 55208 117372 55214
rect 117320 55150 117372 55156
rect 118712 54777 118740 57559
rect 153304 56409 153332 57831
rect 155958 57624 156014 57633
rect 155958 57559 156014 57568
rect 153290 56400 153346 56409
rect 153290 56335 153346 56344
rect 155972 54913 156000 57559
rect 157444 55894 157472 57831
rect 183336 57831 183338 57840
rect 183284 57802 183336 57808
rect 197372 57798 197400 162318
rect 197464 162246 197492 162862
rect 197452 162240 197504 162246
rect 197452 162182 197504 162188
rect 197464 57866 197492 162182
rect 197556 146266 197584 250446
rect 197544 146260 197596 146266
rect 197544 146202 197596 146208
rect 197648 146198 197676 250514
rect 197832 162178 197860 258046
rect 198752 244225 198780 349551
rect 199014 289776 199070 289785
rect 199014 289711 199070 289720
rect 198830 288416 198886 288425
rect 198830 288351 198886 288360
rect 198844 287745 198872 288351
rect 198830 287736 198886 287745
rect 198830 287671 198886 287680
rect 198738 244216 198794 244225
rect 198738 244151 198794 244160
rect 198844 183569 198872 287671
rect 198922 283112 198978 283121
rect 198922 283047 198978 283056
rect 198830 183560 198886 183569
rect 198830 183495 198886 183504
rect 198830 182064 198886 182073
rect 198830 181999 198886 182008
rect 198844 181393 198872 181999
rect 198830 181384 198886 181393
rect 198830 181319 198886 181328
rect 198738 179480 198794 179489
rect 198738 179415 198794 179424
rect 198004 173188 198056 173194
rect 198004 173130 198056 173136
rect 197820 162172 197872 162178
rect 197820 162114 197872 162120
rect 197636 146192 197688 146198
rect 197636 146134 197688 146140
rect 198016 145586 198044 173130
rect 198004 145580 198056 145586
rect 198004 145522 198056 145528
rect 198752 74905 198780 179415
rect 198844 76401 198872 181319
rect 198936 178673 198964 283047
rect 199028 184385 199056 289711
rect 199396 288425 199424 366318
rect 199488 362234 199516 372671
rect 199476 362228 199528 362234
rect 199476 362170 199528 362176
rect 199382 288416 199438 288425
rect 199382 288351 199438 288360
rect 199488 287054 199516 362170
rect 199580 358086 199608 390759
rect 199658 388512 199714 388521
rect 199658 388447 199714 388456
rect 199568 358080 199620 358086
rect 199568 358022 199620 358028
rect 199120 287026 199516 287054
rect 199120 284889 199148 287026
rect 199580 286385 199608 358022
rect 199672 354006 199700 388447
rect 200224 374814 200252 476086
rect 200396 475652 200448 475658
rect 200396 475594 200448 475600
rect 200304 475584 200356 475590
rect 200304 475526 200356 475532
rect 200212 374808 200264 374814
rect 200212 374750 200264 374756
rect 199750 373824 199806 373833
rect 200316 373794 200344 475526
rect 200408 373862 200436 475594
rect 200776 466454 200804 480023
rect 201500 478236 201552 478242
rect 201500 478178 201552 478184
rect 201512 478009 201540 478178
rect 201498 478000 201554 478009
rect 201498 477935 201554 477944
rect 201500 471300 201552 471306
rect 201500 471242 201552 471248
rect 200684 466426 200804 466454
rect 200580 465928 200632 465934
rect 200580 465870 200632 465876
rect 200488 463208 200540 463214
rect 200488 463150 200540 463156
rect 200500 374610 200528 463150
rect 200592 393378 200620 465870
rect 200580 393372 200632 393378
rect 200580 393314 200632 393320
rect 200580 393236 200632 393242
rect 200580 393178 200632 393184
rect 200488 374604 200540 374610
rect 200488 374546 200540 374552
rect 200396 373856 200448 373862
rect 200396 373798 200448 373804
rect 199750 373759 199806 373768
rect 200304 373788 200356 373794
rect 199764 366382 199792 373759
rect 200304 373730 200356 373736
rect 200592 373454 200620 393178
rect 200684 374746 200712 466426
rect 200764 466336 200816 466342
rect 200764 466278 200816 466284
rect 200672 374740 200724 374746
rect 200672 374682 200724 374688
rect 200580 373448 200632 373454
rect 200580 373390 200632 373396
rect 199752 366376 199804 366382
rect 199752 366318 199804 366324
rect 199752 359508 199804 359514
rect 199752 359450 199804 359456
rect 199660 354000 199712 354006
rect 199660 353942 199712 353948
rect 199566 286376 199622 286385
rect 199566 286311 199622 286320
rect 199106 284880 199162 284889
rect 199106 284815 199162 284824
rect 199014 184376 199070 184385
rect 199014 184311 199070 184320
rect 198922 178664 198978 178673
rect 198922 178599 198978 178608
rect 198830 76392 198886 76401
rect 198830 76327 198886 76336
rect 198738 74896 198794 74905
rect 198738 74831 198794 74840
rect 198936 73681 198964 178599
rect 199028 79393 199056 184311
rect 199120 179489 199148 284815
rect 199580 277394 199608 286311
rect 199672 283121 199700 353942
rect 199764 289785 199792 359450
rect 199750 289776 199806 289785
rect 199750 289711 199806 289720
rect 199658 283112 199714 283121
rect 199658 283047 199714 283056
rect 199304 277366 199608 277394
rect 199198 244216 199254 244225
rect 199198 244151 199254 244160
rect 199106 179480 199162 179489
rect 199106 179415 199162 179424
rect 199212 139233 199240 244151
rect 199304 182073 199332 277366
rect 200776 268530 200804 466278
rect 201040 465452 201092 465458
rect 201040 465394 201092 465400
rect 200856 463684 200908 463690
rect 200856 463626 200908 463632
rect 200764 268524 200816 268530
rect 200764 268466 200816 268472
rect 200868 267510 200896 463626
rect 200948 459536 201000 459542
rect 200948 459478 201000 459484
rect 200960 280158 200988 459478
rect 201052 383654 201080 465394
rect 201052 383626 201172 383654
rect 201040 371204 201092 371210
rect 201040 371146 201092 371152
rect 201052 364342 201080 371146
rect 201144 369442 201172 383626
rect 201406 375320 201462 375329
rect 201406 375255 201462 375264
rect 201132 369436 201184 369442
rect 201132 369378 201184 369384
rect 201040 364336 201092 364342
rect 201040 364278 201092 364284
rect 200948 280152 201000 280158
rect 200948 280094 201000 280100
rect 200856 267504 200908 267510
rect 200856 267446 200908 267452
rect 201052 267034 201080 364278
rect 200120 267028 200172 267034
rect 200120 266970 200172 266976
rect 201040 267028 201092 267034
rect 201040 266970 201092 266976
rect 199382 183560 199438 183569
rect 199382 183495 199438 183504
rect 199396 182753 199424 183495
rect 199382 182744 199438 182753
rect 199382 182679 199438 182688
rect 199290 182064 199346 182073
rect 199290 181999 199346 182008
rect 199198 139224 199254 139233
rect 199198 139159 199254 139168
rect 199014 79384 199070 79393
rect 199014 79319 199070 79328
rect 199396 77761 199424 182679
rect 200132 162926 200160 266970
rect 200120 162920 200172 162926
rect 200120 162862 200172 162868
rect 199382 77752 199438 77761
rect 199382 77687 199438 77696
rect 198922 73672 198978 73681
rect 198922 73607 198978 73616
rect 201420 58818 201448 375255
rect 201512 371210 201540 471242
rect 201604 466454 201632 480023
rect 201696 480023 201986 480051
rect 202064 480023 202446 480051
rect 202906 480023 203012 480051
rect 201696 471306 201724 480023
rect 201684 471300 201736 471306
rect 201684 471242 201736 471248
rect 202064 466454 202092 480023
rect 202984 476114 203012 480023
rect 202892 476086 203012 476114
rect 203076 480023 203274 480051
rect 203076 476114 203104 480023
rect 203076 476086 203196 476114
rect 202892 471594 202920 476086
rect 202800 471566 202920 471594
rect 202800 471322 202828 471566
rect 202800 471294 203012 471322
rect 202880 471232 202932 471238
rect 202880 471174 202932 471180
rect 202144 467220 202196 467226
rect 202144 467162 202196 467168
rect 201604 466426 201724 466454
rect 201592 465724 201644 465730
rect 201592 465666 201644 465672
rect 201500 371204 201552 371210
rect 201500 371146 201552 371152
rect 201604 267850 201632 465666
rect 201696 374678 201724 466426
rect 201788 466426 202092 466454
rect 201684 374672 201736 374678
rect 201684 374614 201736 374620
rect 201788 374610 201816 466426
rect 201868 463072 201920 463078
rect 201868 463014 201920 463020
rect 201776 374604 201828 374610
rect 201776 374546 201828 374552
rect 201592 267844 201644 267850
rect 201592 267786 201644 267792
rect 201880 267442 201908 463014
rect 201960 461032 202012 461038
rect 201960 460974 202012 460980
rect 201972 354754 202000 460974
rect 201960 354748 202012 354754
rect 201960 354690 202012 354696
rect 201868 267436 201920 267442
rect 201868 267378 201920 267384
rect 202156 162314 202184 467162
rect 202328 462868 202380 462874
rect 202328 462810 202380 462816
rect 202236 462052 202288 462058
rect 202236 461994 202288 462000
rect 202248 267442 202276 461994
rect 202340 268734 202368 462810
rect 202420 458788 202472 458794
rect 202420 458730 202472 458736
rect 202432 369510 202460 458730
rect 202786 375320 202842 375329
rect 202786 375255 202842 375264
rect 202420 369504 202472 369510
rect 202420 369446 202472 369452
rect 202328 268728 202380 268734
rect 202328 268670 202380 268676
rect 202236 267436 202288 267442
rect 202236 267378 202288 267384
rect 202144 162308 202196 162314
rect 202144 162250 202196 162256
rect 201408 58812 201460 58818
rect 201408 58754 201460 58760
rect 202800 58750 202828 375255
rect 202892 369782 202920 471174
rect 202880 369776 202932 369782
rect 202880 369718 202932 369724
rect 202984 369714 203012 471294
rect 203064 471300 203116 471306
rect 203064 471242 203116 471248
rect 203076 372706 203104 471242
rect 203168 471238 203196 476086
rect 203524 475992 203576 475998
rect 203524 475934 203576 475940
rect 203156 471232 203208 471238
rect 203156 471174 203208 471180
rect 203156 465860 203208 465866
rect 203156 465802 203208 465808
rect 203168 374474 203196 465802
rect 203248 462188 203300 462194
rect 203248 462130 203300 462136
rect 203156 374468 203208 374474
rect 203156 374410 203208 374416
rect 203260 374066 203288 462130
rect 203248 374060 203300 374066
rect 203248 374002 203300 374008
rect 203064 372700 203116 372706
rect 203064 372642 203116 372648
rect 203076 370326 203104 372642
rect 203064 370320 203116 370326
rect 203064 370262 203116 370268
rect 202972 369708 203024 369714
rect 202972 369650 203024 369656
rect 202880 356720 202932 356726
rect 202880 356662 202932 356668
rect 202892 267102 202920 356662
rect 203536 267578 203564 475934
rect 203720 475318 203748 480037
rect 203904 480023 204194 480051
rect 204272 480023 204654 480051
rect 203708 475312 203760 475318
rect 203708 475254 203760 475260
rect 203904 471306 203932 480023
rect 203892 471300 203944 471306
rect 203892 471242 203944 471248
rect 203708 467152 203760 467158
rect 203708 467094 203760 467100
rect 203616 460352 203668 460358
rect 203616 460294 203668 460300
rect 203524 267572 203576 267578
rect 203524 267514 203576 267520
rect 202880 267096 202932 267102
rect 202880 267038 202932 267044
rect 203524 250504 203576 250510
rect 203524 250446 203576 250452
rect 203536 249830 203564 250446
rect 203524 249824 203576 249830
rect 203524 249766 203576 249772
rect 203536 173874 203564 249766
rect 203524 173868 203576 173874
rect 203524 173810 203576 173816
rect 203628 164286 203656 460294
rect 203720 267617 203748 467094
rect 203892 465656 203944 465662
rect 203892 465598 203944 465604
rect 203800 460692 203852 460698
rect 203800 460634 203852 460640
rect 203812 268666 203840 460634
rect 203904 369374 203932 465598
rect 204272 373658 204300 480023
rect 204352 478576 204404 478582
rect 204350 478544 204352 478553
rect 204404 478544 204406 478553
rect 204350 478479 204406 478488
rect 204904 478100 204956 478106
rect 204904 478042 204956 478048
rect 204352 471300 204404 471306
rect 204352 471242 204404 471248
rect 204364 457502 204392 471242
rect 204444 465792 204496 465798
rect 204444 465734 204496 465740
rect 204352 457496 204404 457502
rect 204352 457438 204404 457444
rect 204456 374542 204484 465734
rect 204444 374536 204496 374542
rect 204444 374478 204496 374484
rect 204260 373652 204312 373658
rect 204260 373594 204312 373600
rect 204272 373386 204300 373594
rect 204260 373380 204312 373386
rect 204260 373322 204312 373328
rect 204168 371952 204220 371958
rect 204168 371894 204220 371900
rect 203892 369368 203944 369374
rect 203892 369310 203944 369316
rect 203800 268660 203852 268666
rect 203800 268602 203852 268608
rect 203706 267608 203762 267617
rect 203706 267543 203762 267552
rect 204180 250646 204208 371894
rect 204168 250640 204220 250646
rect 204168 250582 204220 250588
rect 204168 173868 204220 173874
rect 204168 173810 204220 173816
rect 204180 173194 204208 173810
rect 204168 173188 204220 173194
rect 204168 173130 204220 173136
rect 203616 164280 203668 164286
rect 203616 164222 203668 164228
rect 204916 163878 204944 478042
rect 205008 471238 205036 480037
rect 205192 480023 205482 480051
rect 205192 471306 205220 480023
rect 205640 478712 205692 478718
rect 205638 478680 205640 478689
rect 205692 478680 205694 478689
rect 205638 478615 205694 478624
rect 205640 478508 205692 478514
rect 205640 478450 205692 478456
rect 205652 478417 205680 478450
rect 205638 478408 205694 478417
rect 205638 478343 205694 478352
rect 205456 478236 205508 478242
rect 205456 478178 205508 478184
rect 205180 471300 205232 471306
rect 205180 471242 205232 471248
rect 204996 471232 205048 471238
rect 204996 471174 205048 471180
rect 205088 467288 205140 467294
rect 205088 467230 205140 467236
rect 204996 463344 205048 463350
rect 204996 463286 205048 463292
rect 204904 163872 204956 163878
rect 204904 163814 204956 163820
rect 205008 162586 205036 463286
rect 205100 267170 205128 467230
rect 205180 466268 205232 466274
rect 205180 466210 205232 466216
rect 205192 268598 205220 466210
rect 205272 460556 205324 460562
rect 205272 460498 205324 460504
rect 205284 269278 205312 460498
rect 205364 459468 205416 459474
rect 205364 459410 205416 459416
rect 205376 369646 205404 459410
rect 205468 373969 205496 478178
rect 205732 475380 205784 475386
rect 205732 475322 205784 475328
rect 205640 463004 205692 463010
rect 205640 462946 205692 462952
rect 205546 456920 205602 456929
rect 205546 456855 205602 456864
rect 205454 373960 205510 373969
rect 205454 373895 205510 373904
rect 205468 373697 205496 373895
rect 205454 373688 205510 373697
rect 205454 373623 205510 373632
rect 205364 369640 205416 369646
rect 205364 369582 205416 369588
rect 205272 269272 205324 269278
rect 205272 269214 205324 269220
rect 205180 268592 205232 268598
rect 205180 268534 205232 268540
rect 205088 267164 205140 267170
rect 205088 267106 205140 267112
rect 204996 162580 205048 162586
rect 204996 162522 205048 162528
rect 204904 145580 204956 145586
rect 204904 145522 204956 145528
rect 204916 67658 204944 145522
rect 204904 67652 204956 67658
rect 204904 67594 204956 67600
rect 202788 58744 202840 58750
rect 202788 58686 202840 58692
rect 204916 57934 204944 67594
rect 205560 59090 205588 456855
rect 205652 267714 205680 462946
rect 205744 409154 205772 475322
rect 205928 474162 205956 480037
rect 206020 480023 206402 480051
rect 206480 480023 206862 480051
rect 207230 480023 207336 480051
rect 205916 474156 205968 474162
rect 205916 474098 205968 474104
rect 206020 470594 206048 480023
rect 206480 475386 206508 480023
rect 207112 478916 207164 478922
rect 207112 478858 207164 478864
rect 206468 475380 206520 475386
rect 206468 475322 206520 475328
rect 206560 474088 206612 474094
rect 206560 474030 206612 474036
rect 205836 470566 206048 470594
rect 205836 413982 205864 470566
rect 205916 468716 205968 468722
rect 205916 468658 205968 468664
rect 205824 413976 205876 413982
rect 205824 413918 205876 413924
rect 205824 411936 205876 411942
rect 205824 411878 205876 411884
rect 205732 409148 205784 409154
rect 205732 409090 205784 409096
rect 205836 373522 205864 411878
rect 205928 374202 205956 468658
rect 206284 466404 206336 466410
rect 206284 466346 206336 466352
rect 205916 374196 205968 374202
rect 205916 374138 205968 374144
rect 205824 373516 205876 373522
rect 205824 373458 205876 373464
rect 206296 369102 206324 466346
rect 206468 461712 206520 461718
rect 206468 461654 206520 461660
rect 206376 460420 206428 460426
rect 206376 460362 206428 460368
rect 206284 369096 206336 369102
rect 206284 369038 206336 369044
rect 205640 267708 205692 267714
rect 205640 267650 205692 267656
rect 206388 163742 206416 460362
rect 206480 173806 206508 461654
rect 206572 266966 206600 474030
rect 206652 463548 206704 463554
rect 206652 463490 206704 463496
rect 206664 269210 206692 463490
rect 207020 460964 207072 460970
rect 207020 460906 207072 460912
rect 206744 459264 206796 459270
rect 206744 459206 206796 459212
rect 206756 278730 206784 459206
rect 207032 383654 207060 460906
rect 206940 383648 207072 383654
rect 206940 383626 207020 383648
rect 206834 375320 206890 375329
rect 206834 375255 206890 375264
rect 206744 278724 206796 278730
rect 206744 278666 206796 278672
rect 206652 269204 206704 269210
rect 206652 269146 206704 269152
rect 206560 266960 206612 266966
rect 206560 266902 206612 266908
rect 206468 173800 206520 173806
rect 206468 173742 206520 173748
rect 206376 163736 206428 163742
rect 206376 163678 206428 163684
rect 205548 59084 205600 59090
rect 205548 59026 205600 59032
rect 206848 58886 206876 375255
rect 206940 356114 206968 383626
rect 207020 383590 207072 383596
rect 206928 356108 206980 356114
rect 206928 356050 206980 356056
rect 207124 267374 207152 478858
rect 207204 475380 207256 475386
rect 207204 475322 207256 475328
rect 207216 373182 207244 475322
rect 207308 467158 207336 480023
rect 207400 480023 207690 480051
rect 207768 480023 208150 480051
rect 208412 480023 208610 480051
rect 208688 480023 209070 480051
rect 207296 467152 207348 467158
rect 207296 467094 207348 467100
rect 207400 458250 207428 480023
rect 207768 475386 207796 480023
rect 207756 475380 207808 475386
rect 207756 475322 207808 475328
rect 207664 469872 207716 469878
rect 207664 469814 207716 469820
rect 207480 468580 207532 468586
rect 207480 468522 207532 468528
rect 207388 458244 207440 458250
rect 207388 458186 207440 458192
rect 207296 413976 207348 413982
rect 207296 413918 207348 413924
rect 207308 407794 207336 413918
rect 207296 407788 207348 407794
rect 207296 407730 207348 407736
rect 207492 374270 207520 468522
rect 207480 374264 207532 374270
rect 207480 374206 207532 374212
rect 207204 373176 207256 373182
rect 207204 373118 207256 373124
rect 207216 369850 207244 373118
rect 207204 369844 207256 369850
rect 207204 369786 207256 369792
rect 207112 267368 207164 267374
rect 207112 267310 207164 267316
rect 207676 70378 207704 469814
rect 207848 468784 207900 468790
rect 207848 468726 207900 468732
rect 207754 459368 207810 459377
rect 207754 459303 207810 459312
rect 207768 163674 207796 459303
rect 207860 266898 207888 468726
rect 208032 459400 208084 459406
rect 208032 459342 208084 459348
rect 207940 459332 207992 459338
rect 207940 459274 207992 459280
rect 207952 269142 207980 459274
rect 208044 368966 208072 459342
rect 208124 458244 208176 458250
rect 208124 458186 208176 458192
rect 208136 413302 208164 458186
rect 208124 413296 208176 413302
rect 208124 413238 208176 413244
rect 208306 407824 208362 407833
rect 208306 407759 208362 407768
rect 208216 371408 208268 371414
rect 208216 371350 208268 371356
rect 208032 368960 208084 368966
rect 208032 368902 208084 368908
rect 207940 269136 207992 269142
rect 207940 269078 207992 269084
rect 207848 266892 207900 266898
rect 207848 266834 207900 266840
rect 208228 265577 208256 371350
rect 208214 265568 208270 265577
rect 208214 265503 208270 265512
rect 207756 163668 207808 163674
rect 207756 163610 207808 163616
rect 207664 70372 207716 70378
rect 207664 70314 207716 70320
rect 206836 58880 206888 58886
rect 206836 58822 206888 58828
rect 204904 57928 204956 57934
rect 204904 57870 204956 57876
rect 197452 57860 197504 57866
rect 197452 57802 197504 57808
rect 183468 57792 183520 57798
rect 183466 57760 183468 57769
rect 197360 57792 197412 57798
rect 183520 57760 183522 57769
rect 197360 57734 197412 57740
rect 208320 57730 208348 407759
rect 208412 374270 208440 480023
rect 208492 478644 208544 478650
rect 208492 478586 208544 478592
rect 208504 478553 208532 478586
rect 208490 478544 208546 478553
rect 208490 478479 208546 478488
rect 208688 470594 208716 480023
rect 209424 477562 209452 480037
rect 209898 480023 210004 480051
rect 209412 477556 209464 477562
rect 209412 477498 209464 477504
rect 209976 475522 210004 480023
rect 210068 480023 210358 480051
rect 210528 480023 210818 480051
rect 211186 480023 211292 480051
rect 209964 475516 210016 475522
rect 209964 475458 210016 475464
rect 210068 475402 210096 480023
rect 210332 477556 210384 477562
rect 210332 477498 210384 477504
rect 210240 476944 210292 476950
rect 210240 476886 210292 476892
rect 210148 475516 210200 475522
rect 210148 475458 210200 475464
rect 209780 475380 209832 475386
rect 209780 475322 209832 475328
rect 209884 475374 210096 475402
rect 209504 475312 209556 475318
rect 209504 475254 209556 475260
rect 209228 471436 209280 471442
rect 209228 471378 209280 471384
rect 208504 470566 208716 470594
rect 208504 374474 208532 470566
rect 209042 466032 209098 466041
rect 209042 465967 209098 465976
rect 208584 463140 208636 463146
rect 208584 463082 208636 463088
rect 208492 374468 208544 374474
rect 208492 374410 208544 374416
rect 208596 374338 208624 463082
rect 208952 462120 209004 462126
rect 208952 462062 209004 462068
rect 208584 374332 208636 374338
rect 208584 374274 208636 374280
rect 208400 374264 208452 374270
rect 208400 374206 208452 374212
rect 208412 369034 208440 374206
rect 208964 373994 208992 462062
rect 208872 373966 208992 373994
rect 208400 369028 208452 369034
rect 208400 368970 208452 368976
rect 208872 368898 208900 373966
rect 208950 369200 209006 369209
rect 208950 369135 209006 369144
rect 208860 368892 208912 368898
rect 208860 368834 208912 368840
rect 208400 360188 208452 360194
rect 208400 360130 208452 360136
rect 208412 359514 208440 360130
rect 208400 359508 208452 359514
rect 208400 359450 208452 359456
rect 208964 59022 208992 369135
rect 209056 162178 209084 465967
rect 209136 463412 209188 463418
rect 209136 463354 209188 463360
rect 209148 163606 209176 463354
rect 209240 267646 209268 471378
rect 209320 466200 209372 466206
rect 209320 466142 209372 466148
rect 209332 268802 209360 466142
rect 209412 460624 209464 460630
rect 209412 460566 209464 460572
rect 209320 268796 209372 268802
rect 209320 268738 209372 268744
rect 209228 267640 209280 267646
rect 209228 267582 209280 267588
rect 209424 266801 209452 460566
rect 209516 385014 209544 475254
rect 209504 385008 209556 385014
rect 209504 384950 209556 384956
rect 209688 373516 209740 373522
rect 209688 373458 209740 373464
rect 209596 371476 209648 371482
rect 209596 371418 209648 371424
rect 209504 370524 209556 370530
rect 209504 370466 209556 370472
rect 209516 268462 209544 370466
rect 209504 268456 209556 268462
rect 209504 268398 209556 268404
rect 209410 266792 209466 266801
rect 209410 266727 209466 266736
rect 209608 265713 209636 371418
rect 209700 360194 209728 373458
rect 209792 372298 209820 475322
rect 209884 372570 209912 475374
rect 210160 475266 210188 475458
rect 209976 475238 210188 475266
rect 209976 374066 210004 475238
rect 210252 475130 210280 476886
rect 210344 475250 210372 477498
rect 210424 475788 210476 475794
rect 210424 475730 210476 475736
rect 210436 475266 210464 475730
rect 210528 475386 210556 480023
rect 211264 475522 211292 480023
rect 211356 480023 211646 480051
rect 211252 475516 211304 475522
rect 211252 475458 211304 475464
rect 211356 475402 211384 480023
rect 212092 477562 212120 480037
rect 212566 480023 212672 480051
rect 212540 478848 212592 478854
rect 212540 478790 212592 478796
rect 212552 478145 212580 478790
rect 212538 478136 212594 478145
rect 212538 478071 212594 478080
rect 212080 477556 212132 477562
rect 212080 477498 212132 477504
rect 212080 475924 212132 475930
rect 212080 475866 212132 475872
rect 211804 475856 211856 475862
rect 211804 475798 211856 475804
rect 210516 475380 210568 475386
rect 210516 475322 210568 475328
rect 211172 475374 211384 475402
rect 210332 475244 210384 475250
rect 210436 475238 210556 475266
rect 210332 475186 210384 475192
rect 210252 475102 210464 475130
rect 210332 475040 210384 475046
rect 210332 474982 210384 474988
rect 210240 374468 210292 374474
rect 210240 374410 210292 374416
rect 209964 374060 210016 374066
rect 209964 374002 210016 374008
rect 210148 372768 210200 372774
rect 210148 372710 210200 372716
rect 209872 372564 209924 372570
rect 209872 372506 209924 372512
rect 209780 372292 209832 372298
rect 209780 372234 209832 372240
rect 210160 372162 210188 372710
rect 210148 372156 210200 372162
rect 210148 372098 210200 372104
rect 210054 371920 210110 371929
rect 210054 371855 210110 371864
rect 210068 371657 210096 371855
rect 210054 371648 210110 371657
rect 210054 371583 210110 371592
rect 210252 371550 210280 374410
rect 210344 372774 210372 474982
rect 210332 372768 210384 372774
rect 210332 372710 210384 372716
rect 210332 372564 210384 372570
rect 210332 372506 210384 372512
rect 210344 372094 210372 372506
rect 210332 372088 210384 372094
rect 210332 372030 210384 372036
rect 210330 371920 210386 371929
rect 210330 371855 210386 371864
rect 210240 371544 210292 371550
rect 210344 371521 210372 371855
rect 210240 371486 210292 371492
rect 210330 371512 210386 371521
rect 210330 371447 210386 371456
rect 210240 369164 210292 369170
rect 210240 369106 210292 369112
rect 209688 360188 209740 360194
rect 209688 360130 209740 360136
rect 209594 265704 209650 265713
rect 209594 265639 209650 265648
rect 209594 265568 209650 265577
rect 209594 265503 209650 265512
rect 209136 163600 209188 163606
rect 209136 163542 209188 163548
rect 209044 162172 209096 162178
rect 209044 162114 209096 162120
rect 209608 144906 209636 265503
rect 210252 264314 210280 369106
rect 210240 264308 210292 264314
rect 210240 264250 210292 264256
rect 210344 263702 210372 371447
rect 210332 263696 210384 263702
rect 210332 263638 210384 263644
rect 210436 162450 210464 475102
rect 210424 162444 210476 162450
rect 210424 162386 210476 162392
rect 210528 162110 210556 475238
rect 210608 472728 210660 472734
rect 210608 472670 210660 472676
rect 210620 162858 210648 472670
rect 210792 466064 210844 466070
rect 210792 466006 210844 466012
rect 210700 463276 210752 463282
rect 210700 463218 210752 463224
rect 210712 164354 210740 463218
rect 210804 269346 210832 466006
rect 210884 459196 210936 459202
rect 210884 459138 210936 459144
rect 210792 269340 210844 269346
rect 210792 269282 210844 269288
rect 210896 267102 210924 459138
rect 211066 375320 211122 375329
rect 211066 375255 211122 375264
rect 210974 372736 211030 372745
rect 210974 372671 211030 372680
rect 210884 267096 210936 267102
rect 210884 267038 210936 267044
rect 210700 164348 210752 164354
rect 210700 164290 210752 164296
rect 210608 162852 210660 162858
rect 210608 162794 210660 162800
rect 210516 162104 210568 162110
rect 210516 162046 210568 162052
rect 209596 144900 209648 144906
rect 209596 144842 209648 144848
rect 208952 59016 209004 59022
rect 208952 58958 209004 58964
rect 210988 57934 211016 372671
rect 210976 57928 211028 57934
rect 210976 57870 211028 57876
rect 183466 57695 183522 57704
rect 208308 57724 208360 57730
rect 208308 57666 208360 57672
rect 160098 57624 160154 57633
rect 160098 57559 160154 57568
rect 165618 57624 165674 57633
rect 165618 57559 165674 57568
rect 157432 55888 157484 55894
rect 157432 55830 157484 55836
rect 160112 55049 160140 57559
rect 165632 55185 165660 57559
rect 211080 57526 211108 375255
rect 211172 372366 211200 475374
rect 211252 475312 211304 475318
rect 211252 475254 211304 475260
rect 211160 372360 211212 372366
rect 211160 372302 211212 372308
rect 211264 371686 211292 475254
rect 211344 458924 211396 458930
rect 211344 458866 211396 458872
rect 211356 374406 211384 458866
rect 211528 391264 211580 391270
rect 211528 391206 211580 391212
rect 211344 374400 211396 374406
rect 211344 374342 211396 374348
rect 211252 371680 211304 371686
rect 211252 371622 211304 371628
rect 211540 369578 211568 391206
rect 211712 374332 211764 374338
rect 211712 374274 211764 374280
rect 211724 374066 211752 374274
rect 211712 374060 211764 374066
rect 211712 374002 211764 374008
rect 211724 372570 211752 374002
rect 211712 372564 211764 372570
rect 211712 372506 211764 372512
rect 211618 372192 211674 372201
rect 211618 372127 211674 372136
rect 211632 369594 211660 372127
rect 211724 371822 211752 372506
rect 211712 371816 211764 371822
rect 211712 371758 211764 371764
rect 211528 369572 211580 369578
rect 211632 369566 211752 369594
rect 211528 369514 211580 369520
rect 211620 369232 211672 369238
rect 211620 369174 211672 369180
rect 211632 269006 211660 369174
rect 211620 269000 211672 269006
rect 211620 268942 211672 268948
rect 211724 264858 211752 369566
rect 211712 264852 211764 264858
rect 211712 264794 211764 264800
rect 211724 263634 211752 264794
rect 211712 263628 211764 263634
rect 211712 263570 211764 263576
rect 211816 162722 211844 475798
rect 211896 471368 211948 471374
rect 211896 471310 211948 471316
rect 211804 162716 211856 162722
rect 211804 162658 211856 162664
rect 211908 162246 211936 471310
rect 211986 465896 212042 465905
rect 211986 465831 212042 465840
rect 212000 163946 212028 465831
rect 212092 267481 212120 475866
rect 212540 475312 212592 475318
rect 212540 475254 212592 475260
rect 212264 462936 212316 462942
rect 212264 462878 212316 462884
rect 212172 461916 212224 461922
rect 212172 461858 212224 461864
rect 212184 268870 212212 461858
rect 212276 383382 212304 462878
rect 212264 383376 212316 383382
rect 212264 383318 212316 383324
rect 212446 382392 212502 382401
rect 212446 382327 212502 382336
rect 212354 375320 212410 375329
rect 212354 375255 212410 375264
rect 212262 371784 212318 371793
rect 212262 371719 212318 371728
rect 212172 268864 212224 268870
rect 212172 268806 212224 268812
rect 212276 267734 212304 371719
rect 212184 267706 212304 267734
rect 212078 267472 212134 267481
rect 212078 267407 212134 267416
rect 212184 264926 212212 267706
rect 212172 264920 212224 264926
rect 212172 264862 212224 264868
rect 212080 263628 212132 263634
rect 212080 263570 212132 263576
rect 211988 163940 212040 163946
rect 211988 163882 212040 163888
rect 211896 162240 211948 162246
rect 211896 162182 211948 162188
rect 212092 144634 212120 263570
rect 212184 160478 212212 264862
rect 212172 160472 212224 160478
rect 212172 160414 212224 160420
rect 212080 144628 212132 144634
rect 212080 144570 212132 144576
rect 212368 57866 212396 375255
rect 212356 57860 212408 57866
rect 212356 57802 212408 57808
rect 211068 57520 211120 57526
rect 211068 57462 211120 57468
rect 212460 57390 212488 382327
rect 212552 372774 212580 475254
rect 212644 379846 212672 480023
rect 212828 480023 213026 480051
rect 213104 480023 213394 480051
rect 213472 480023 213854 480051
rect 214024 480023 214314 480051
rect 214392 480023 214774 480051
rect 214944 480023 215234 480051
rect 212724 475380 212776 475386
rect 212724 475322 212776 475328
rect 212632 379840 212684 379846
rect 212632 379782 212684 379788
rect 212736 373994 212764 475322
rect 212644 373966 212764 373994
rect 212828 373994 212856 480023
rect 213104 475386 213132 480023
rect 213092 475380 213144 475386
rect 213092 475322 213144 475328
rect 213472 475318 213500 480023
rect 213920 478780 213972 478786
rect 213920 478722 213972 478728
rect 213932 478689 213960 478722
rect 213918 478680 213974 478689
rect 213918 478615 213974 478624
rect 213920 475380 213972 475386
rect 213920 475322 213972 475328
rect 213460 475312 213512 475318
rect 213460 475254 213512 475260
rect 213092 462800 213144 462806
rect 213092 462742 213144 462748
rect 212908 461780 212960 461786
rect 212908 461722 212960 461728
rect 212920 460970 212948 461722
rect 212908 460964 212960 460970
rect 212908 460906 212960 460912
rect 212920 374649 212948 460906
rect 212906 374640 212962 374649
rect 212906 374575 212962 374584
rect 212828 373966 212948 373994
rect 212644 372978 212672 373966
rect 212920 373046 212948 373966
rect 212908 373040 212960 373046
rect 212908 372982 212960 372988
rect 212632 372972 212684 372978
rect 212632 372914 212684 372920
rect 212540 372768 212592 372774
rect 212540 372710 212592 372716
rect 212552 369238 212580 372710
rect 212540 369232 212592 369238
rect 212540 369174 212592 369180
rect 212644 369170 212672 372914
rect 212920 372638 212948 372982
rect 212908 372632 212960 372638
rect 212908 372574 212960 372580
rect 212920 370326 212948 372574
rect 212908 370320 212960 370326
rect 212908 370262 212960 370268
rect 212632 369164 212684 369170
rect 212632 369106 212684 369112
rect 213104 369034 213132 462742
rect 213276 461984 213328 461990
rect 213276 461926 213328 461932
rect 213182 459096 213238 459105
rect 213182 459031 213238 459040
rect 213092 369028 213144 369034
rect 213092 368970 213144 368976
rect 213196 163810 213224 459031
rect 213288 267345 213316 461926
rect 213368 461848 213420 461854
rect 213368 461790 213420 461796
rect 213274 267336 213330 267345
rect 213274 267271 213330 267280
rect 213380 266762 213408 461790
rect 213460 379840 213512 379846
rect 213460 379782 213512 379788
rect 213472 373318 213500 379782
rect 213460 373312 213512 373318
rect 213460 373254 213512 373260
rect 213932 373250 213960 475322
rect 213920 373244 213972 373250
rect 213920 373186 213972 373192
rect 213552 373176 213604 373182
rect 213552 373118 213604 373124
rect 213460 372020 213512 372026
rect 213460 371962 213512 371968
rect 213472 371686 213500 371962
rect 213460 371680 213512 371686
rect 213460 371622 213512 371628
rect 213460 370320 213512 370326
rect 213460 370262 213512 370268
rect 213472 268938 213500 370262
rect 213564 269074 213592 373118
rect 213736 372564 213788 372570
rect 213736 372506 213788 372512
rect 213642 371648 213698 371657
rect 213642 371583 213698 371592
rect 213552 269068 213604 269074
rect 213552 269010 213604 269016
rect 213460 268932 213512 268938
rect 213460 268874 213512 268880
rect 213656 267734 213684 371583
rect 213472 267706 213684 267734
rect 213368 266756 213420 266762
rect 213368 266698 213420 266704
rect 213472 266257 213500 267706
rect 213748 266286 213776 372506
rect 213932 370530 213960 373186
rect 214024 372910 214052 480023
rect 214392 470594 214420 480023
rect 214564 477012 214616 477018
rect 214564 476954 214616 476960
rect 214116 470566 214420 470594
rect 214116 373114 214144 470566
rect 214196 468512 214248 468518
rect 214196 468454 214248 468460
rect 214208 393990 214236 468454
rect 214196 393984 214248 393990
rect 214196 393926 214248 393932
rect 214208 373522 214236 393926
rect 214196 373516 214248 373522
rect 214196 373458 214248 373464
rect 214104 373108 214156 373114
rect 214104 373050 214156 373056
rect 214012 372904 214064 372910
rect 214012 372846 214064 372852
rect 213920 370524 213972 370530
rect 213920 370466 213972 370472
rect 214024 369306 214052 372846
rect 214012 369300 214064 369306
rect 214012 369242 214064 369248
rect 213826 369200 213882 369209
rect 213826 369135 213882 369144
rect 213736 266280 213788 266286
rect 213458 266248 213514 266257
rect 213736 266222 213788 266228
rect 213458 266183 213514 266192
rect 213366 265160 213422 265169
rect 213366 265095 213422 265104
rect 213184 163804 213236 163810
rect 213184 163746 213236 163752
rect 213276 160744 213328 160750
rect 213276 160686 213328 160692
rect 213288 160478 213316 160686
rect 213276 160472 213328 160478
rect 213276 160414 213328 160420
rect 213184 147688 213236 147694
rect 213184 147630 213236 147636
rect 212448 57384 212500 57390
rect 212448 57326 212500 57332
rect 213196 55758 213224 147630
rect 213184 55752 213236 55758
rect 213184 55694 213236 55700
rect 165618 55176 165674 55185
rect 165618 55111 165674 55120
rect 160098 55040 160154 55049
rect 160098 54975 160154 54984
rect 155958 54904 156014 54913
rect 155958 54839 156014 54848
rect 118698 54768 118754 54777
rect 118698 54703 118754 54712
rect 80060 54606 80112 54612
rect 116122 54632 116178 54641
rect 116122 54567 116178 54576
rect 213288 54466 213316 160414
rect 213380 148986 213408 265095
rect 213368 148980 213420 148986
rect 213368 148922 213420 148928
rect 213276 54460 213328 54466
rect 213276 54402 213328 54408
rect 213380 54398 213408 148922
rect 213472 148374 213500 266183
rect 213644 265124 213696 265130
rect 213644 265066 213696 265072
rect 213552 264240 213604 264246
rect 213552 264182 213604 264188
rect 213564 263702 213592 264182
rect 213552 263696 213604 263702
rect 213552 263638 213604 263644
rect 213460 148368 213512 148374
rect 213460 148310 213512 148316
rect 213460 146328 213512 146334
rect 213460 146270 213512 146276
rect 213472 55894 213500 146270
rect 213564 144702 213592 263638
rect 213656 144770 213684 265066
rect 213748 144838 213776 266222
rect 213736 144832 213788 144838
rect 213736 144774 213788 144780
rect 213644 144764 213696 144770
rect 213644 144706 213696 144712
rect 213552 144696 213604 144702
rect 213552 144638 213604 144644
rect 213840 57594 213868 369135
rect 214116 368830 214144 373050
rect 214472 372564 214524 372570
rect 214472 372506 214524 372512
rect 214484 371890 214512 372506
rect 214472 371884 214524 371890
rect 214472 371826 214524 371832
rect 214380 369300 214432 369306
rect 214380 369242 214432 369248
rect 214104 368824 214156 368830
rect 214104 368766 214156 368772
rect 214392 277394 214420 369242
rect 214472 368824 214524 368830
rect 214472 368766 214524 368772
rect 214300 277366 214420 277394
rect 214300 264994 214328 277366
rect 214484 272626 214512 368766
rect 214392 272598 214512 272626
rect 214392 265062 214420 272598
rect 214472 268456 214524 268462
rect 214472 268398 214524 268404
rect 214484 267782 214512 268398
rect 214472 267776 214524 267782
rect 214472 267718 214524 267724
rect 214380 265056 214432 265062
rect 214380 264998 214432 265004
rect 214288 264988 214340 264994
rect 214288 264930 214340 264936
rect 214392 263022 214420 264998
rect 214380 263016 214432 263022
rect 214380 262958 214432 262964
rect 214484 262834 214512 267718
rect 214300 262806 214512 262834
rect 214300 161294 214328 262806
rect 214472 262744 214524 262750
rect 214472 262686 214524 262692
rect 214484 161474 214512 262686
rect 214576 162790 214604 476954
rect 214656 476876 214708 476882
rect 214656 476818 214708 476824
rect 214564 162784 214616 162790
rect 214564 162726 214616 162732
rect 214668 162518 214696 476818
rect 214944 475386 214972 480023
rect 214932 475380 214984 475386
rect 214932 475322 214984 475328
rect 215392 475380 215444 475386
rect 215392 475322 215444 475328
rect 215300 475312 215352 475318
rect 215300 475254 215352 475260
rect 214840 469940 214892 469946
rect 214840 469882 214892 469888
rect 214746 459232 214802 459241
rect 214746 459167 214802 459176
rect 214760 163538 214788 459167
rect 214852 267374 214880 469882
rect 214930 466304 214986 466313
rect 214930 466239 214986 466248
rect 214944 268462 214972 466239
rect 215312 373522 215340 475254
rect 215404 373862 215432 475322
rect 215588 470594 215616 480037
rect 215680 480023 216062 480051
rect 216232 480023 216522 480051
rect 215680 475318 215708 480023
rect 215944 477556 215996 477562
rect 215944 477498 215996 477504
rect 215668 475312 215720 475318
rect 215668 475254 215720 475260
rect 215496 470566 215616 470594
rect 215496 374377 215524 470566
rect 215760 459672 215812 459678
rect 215760 459614 215812 459620
rect 215482 374368 215538 374377
rect 215482 374303 215538 374312
rect 215392 373856 215444 373862
rect 215392 373798 215444 373804
rect 215300 373516 215352 373522
rect 215300 373458 215352 373464
rect 215312 372638 215340 373458
rect 215300 372632 215352 372638
rect 215300 372574 215352 372580
rect 215024 371884 215076 371890
rect 215024 371826 215076 371832
rect 214932 268456 214984 268462
rect 214932 268398 214984 268404
rect 214840 267368 214892 267374
rect 214840 267310 214892 267316
rect 215036 267034 215064 371826
rect 215300 371612 215352 371618
rect 215300 371554 215352 371560
rect 215116 371544 215168 371550
rect 215116 371486 215168 371492
rect 215024 267028 215076 267034
rect 215024 266970 215076 266976
rect 214930 265024 214986 265033
rect 214930 264959 214986 264968
rect 214748 163532 214800 163538
rect 214748 163474 214800 163480
rect 214656 162512 214708 162518
rect 214656 162454 214708 162460
rect 214484 161446 214880 161474
rect 214288 161288 214340 161294
rect 214288 161230 214340 161236
rect 214300 160138 214328 161230
rect 214288 160132 214340 160138
rect 214288 160074 214340 160080
rect 214748 160132 214800 160138
rect 214748 160074 214800 160080
rect 214562 145888 214618 145897
rect 214562 145823 214618 145832
rect 214576 144906 214604 145823
rect 214656 145580 214708 145586
rect 214656 145522 214708 145528
rect 214564 144900 214616 144906
rect 214564 144842 214616 144848
rect 213828 57588 213880 57594
rect 213828 57530 213880 57536
rect 213460 55888 213512 55894
rect 213460 55830 213512 55836
rect 213368 54392 213420 54398
rect 213368 54334 213420 54340
rect 214576 54330 214604 144842
rect 214668 144770 214696 145522
rect 214656 144764 214708 144770
rect 214656 144706 214708 144712
rect 214668 54602 214696 144706
rect 214760 59430 214788 160074
rect 214852 160070 214880 161446
rect 214840 160064 214892 160070
rect 214840 160006 214892 160012
rect 214748 59424 214800 59430
rect 214748 59366 214800 59372
rect 214852 59226 214880 160006
rect 214944 148918 214972 264959
rect 215036 149054 215064 266970
rect 215128 266014 215156 371486
rect 215312 371346 215340 371554
rect 215300 371340 215352 371346
rect 215300 371282 215352 371288
rect 215206 369880 215262 369889
rect 215206 369815 215262 369824
rect 215116 266008 215168 266014
rect 215116 265950 215168 265956
rect 215116 264580 215168 264586
rect 215116 264522 215168 264528
rect 215024 149048 215076 149054
rect 215024 148990 215076 148996
rect 214932 148912 214984 148918
rect 214932 148854 214984 148860
rect 214840 59220 214892 59226
rect 214840 59162 214892 59168
rect 214944 56574 214972 148854
rect 215036 147694 215064 148990
rect 215024 147688 215076 147694
rect 215024 147630 215076 147636
rect 215128 145790 215156 264522
rect 215116 145784 215168 145790
rect 215116 145726 215168 145732
rect 215022 145480 215078 145489
rect 215022 145415 215078 145424
rect 215036 144634 215064 145415
rect 215024 144628 215076 144634
rect 215024 144570 215076 144576
rect 214932 56568 214984 56574
rect 214932 56510 214984 56516
rect 215036 56370 215064 144570
rect 215024 56364 215076 56370
rect 215024 56306 215076 56312
rect 214656 54596 214708 54602
rect 214656 54538 214708 54544
rect 215128 54534 215156 145726
rect 215220 58954 215248 369815
rect 215404 369617 215432 373798
rect 215496 371006 215524 374303
rect 215668 372632 215720 372638
rect 215668 372574 215720 372580
rect 215576 371612 215628 371618
rect 215576 371554 215628 371560
rect 215484 371000 215536 371006
rect 215484 370942 215536 370948
rect 215390 369608 215446 369617
rect 215390 369543 215446 369552
rect 215300 368484 215352 368490
rect 215300 368426 215352 368432
rect 215312 367810 215340 368426
rect 215300 367804 215352 367810
rect 215300 367746 215352 367752
rect 215392 269068 215444 269074
rect 215392 269010 215444 269016
rect 215404 267918 215432 269010
rect 215392 267912 215444 267918
rect 215392 267854 215444 267860
rect 215298 266384 215354 266393
rect 215298 266319 215354 266328
rect 215208 58948 215260 58954
rect 215208 58890 215260 58896
rect 215312 57322 215340 266319
rect 215404 145518 215432 267854
rect 215496 265742 215524 370942
rect 215588 266121 215616 371554
rect 215680 370326 215708 372574
rect 215772 372337 215800 459614
rect 215956 374542 215984 477498
rect 216232 475386 216260 480023
rect 216968 477601 216996 480037
rect 217324 478168 217376 478174
rect 217324 478110 217376 478116
rect 216954 477592 217010 477601
rect 216954 477527 217010 477536
rect 217336 477442 217364 478110
rect 217428 477562 217456 480037
rect 217508 478304 217560 478310
rect 217508 478246 217560 478252
rect 217416 477556 217468 477562
rect 217416 477498 217468 477504
rect 217336 477414 217456 477442
rect 216220 475380 216272 475386
rect 216220 475322 216272 475328
rect 217324 474156 217376 474162
rect 217324 474098 217376 474104
rect 216036 474020 216088 474026
rect 216036 473962 216088 473968
rect 215944 374536 215996 374542
rect 215944 374478 215996 374484
rect 215758 372328 215814 372337
rect 215758 372263 215814 372272
rect 215760 372156 215812 372162
rect 215760 372098 215812 372104
rect 215668 370320 215720 370326
rect 215668 370262 215720 370268
rect 215680 369753 215708 370262
rect 215666 369744 215722 369753
rect 215666 369679 215722 369688
rect 215772 354674 215800 372098
rect 215944 356108 215996 356114
rect 215944 356050 215996 356056
rect 215680 354646 215800 354674
rect 215574 266112 215630 266121
rect 215680 266082 215708 354646
rect 215956 278322 215984 356050
rect 215944 278316 215996 278322
rect 215944 278258 215996 278264
rect 215574 266047 215630 266056
rect 215668 266076 215720 266082
rect 215484 265736 215536 265742
rect 215484 265678 215536 265684
rect 215588 265169 215616 266047
rect 215668 266018 215720 266024
rect 215574 265160 215630 265169
rect 215680 265130 215708 266018
rect 215850 265704 215906 265713
rect 215850 265639 215906 265648
rect 215574 265095 215630 265104
rect 215668 265124 215720 265130
rect 215668 265066 215720 265072
rect 215760 264988 215812 264994
rect 215760 264930 215812 264936
rect 215772 159594 215800 264930
rect 215760 159588 215812 159594
rect 215760 159530 215812 159536
rect 215864 151814 215892 265639
rect 215956 250510 215984 278258
rect 215944 250504 215996 250510
rect 215944 250446 215996 250452
rect 216048 162042 216076 473962
rect 216404 466132 216456 466138
rect 216404 466074 216456 466080
rect 216128 463480 216180 463486
rect 216128 463422 216180 463428
rect 216140 267238 216168 463422
rect 216220 459128 216272 459134
rect 216220 459070 216272 459076
rect 216128 267232 216180 267238
rect 216128 267174 216180 267180
rect 216232 266830 216260 459070
rect 216312 372700 216364 372706
rect 216312 372642 216364 372648
rect 216324 267073 216352 372642
rect 216416 369850 216444 466074
rect 217336 422294 217364 474098
rect 216876 422266 217364 422294
rect 216680 409148 216732 409154
rect 216680 409090 216732 409096
rect 216692 408785 216720 409090
rect 216678 408776 216734 408785
rect 216734 408734 216812 408762
rect 216678 408711 216734 408720
rect 216678 407824 216734 407833
rect 216678 407759 216680 407768
rect 216732 407759 216734 407768
rect 216680 407730 216732 407736
rect 216692 388498 216720 407730
rect 216784 388618 216812 408734
rect 216876 406065 216904 422266
rect 216956 413296 217008 413302
rect 216956 413238 217008 413244
rect 216968 411369 216996 413238
rect 216954 411360 217010 411369
rect 216954 411295 217010 411304
rect 217046 410000 217102 410009
rect 217046 409935 217102 409944
rect 216862 406056 216918 406065
rect 216862 405991 216918 406000
rect 216772 388612 216824 388618
rect 216772 388554 216824 388560
rect 216692 388470 216812 388498
rect 216680 385008 216732 385014
rect 216678 384976 216680 384985
rect 216732 384976 216734 384985
rect 216678 384911 216734 384920
rect 216680 383648 216732 383654
rect 216680 383590 216732 383596
rect 216692 383353 216720 383590
rect 216678 383344 216734 383353
rect 216678 383279 216734 383288
rect 216784 378842 216812 388470
rect 216876 383518 216904 405991
rect 216956 388612 217008 388618
rect 216956 388554 217008 388560
rect 216864 383512 216916 383518
rect 216864 383454 216916 383460
rect 216864 383376 216916 383382
rect 216864 383318 216916 383324
rect 216876 383081 216904 383318
rect 216862 383072 216918 383081
rect 216862 383007 216918 383016
rect 216784 378814 216904 378842
rect 216770 375320 216826 375329
rect 216770 375255 216826 375264
rect 216784 374921 216812 375255
rect 216770 374912 216826 374921
rect 216770 374847 216826 374856
rect 216404 369844 216456 369850
rect 216404 369786 216456 369792
rect 216588 368484 216640 368490
rect 216588 368426 216640 368432
rect 216310 267064 216366 267073
rect 216310 266999 216366 267008
rect 216220 266824 216272 266830
rect 216220 266766 216272 266772
rect 216220 266348 216272 266354
rect 216220 266290 216272 266296
rect 216128 266008 216180 266014
rect 216128 265950 216180 265956
rect 216140 265606 216168 265950
rect 216232 265742 216260 266290
rect 216220 265736 216272 265742
rect 216220 265678 216272 265684
rect 216128 265600 216180 265606
rect 216128 265542 216180 265548
rect 216036 162036 216088 162042
rect 216036 161978 216088 161984
rect 215680 151786 215892 151814
rect 215680 148850 215708 151786
rect 215668 148844 215720 148850
rect 215668 148786 215720 148792
rect 215392 145512 215444 145518
rect 215392 145454 215444 145460
rect 215404 145042 215432 145454
rect 215392 145036 215444 145042
rect 215392 144978 215444 144984
rect 215300 57316 215352 57322
rect 215300 57258 215352 57264
rect 215680 56506 215708 148786
rect 215944 148368 215996 148374
rect 215944 148310 215996 148316
rect 215758 146024 215814 146033
rect 215758 145959 215814 145968
rect 215772 59158 215800 145959
rect 215852 144968 215904 144974
rect 215852 144910 215904 144916
rect 215760 59152 215812 59158
rect 215760 59094 215812 59100
rect 215668 56500 215720 56506
rect 215668 56442 215720 56448
rect 215864 55962 215892 144910
rect 215852 55956 215904 55962
rect 215852 55898 215904 55904
rect 215956 55146 215984 148310
rect 216140 145722 216168 265542
rect 216232 146305 216260 265678
rect 216218 146296 216274 146305
rect 216218 146231 216274 146240
rect 216232 146033 216260 146231
rect 216218 146024 216274 146033
rect 216218 145959 216274 145968
rect 216324 145874 216352 266999
rect 216494 266520 216550 266529
rect 216494 266455 216550 266464
rect 216404 159996 216456 160002
rect 216404 159938 216456 159944
rect 216416 159594 216444 159938
rect 216404 159588 216456 159594
rect 216404 159530 216456 159536
rect 216232 145846 216352 145874
rect 216128 145716 216180 145722
rect 216128 145658 216180 145664
rect 216140 144974 216168 145658
rect 216232 145382 216260 145846
rect 216310 145752 216366 145761
rect 216310 145687 216366 145696
rect 216220 145376 216272 145382
rect 216220 145318 216272 145324
rect 216220 145036 216272 145042
rect 216220 144978 216272 144984
rect 216128 144968 216180 144974
rect 216128 144910 216180 144916
rect 216036 144832 216088 144838
rect 216036 144774 216088 144780
rect 215944 55140 215996 55146
rect 215944 55082 215996 55088
rect 216048 54670 216076 144774
rect 216128 144696 216180 144702
rect 216128 144638 216180 144644
rect 216140 55078 216168 144638
rect 216232 55214 216260 144978
rect 216324 144702 216352 145687
rect 216312 144696 216364 144702
rect 216312 144638 216364 144644
rect 216416 58614 216444 159530
rect 216404 58608 216456 58614
rect 216404 58550 216456 58556
rect 216508 57662 216536 266455
rect 216600 265674 216628 368426
rect 216784 299441 216812 374847
rect 216876 373930 216904 378814
rect 216968 375057 216996 388554
rect 216954 375048 217010 375057
rect 216954 374983 217010 374992
rect 216864 373924 216916 373930
rect 216864 373866 216916 373872
rect 216876 302841 216904 373866
rect 216968 303793 216996 374983
rect 217060 373998 217088 409935
rect 217324 383512 217376 383518
rect 217324 383454 217376 383460
rect 217232 375352 217284 375358
rect 217232 375294 217284 375300
rect 217244 375086 217272 375294
rect 217232 375080 217284 375086
rect 217232 375022 217284 375028
rect 217048 373992 217100 373998
rect 217048 373934 217100 373940
rect 217060 372842 217088 373934
rect 217048 372836 217100 372842
rect 217048 372778 217100 372784
rect 217046 372736 217102 372745
rect 217046 372671 217102 372680
rect 217060 371958 217088 372671
rect 217048 371952 217100 371958
rect 217048 371894 217100 371900
rect 217140 370320 217192 370326
rect 217140 370262 217192 370268
rect 216954 303784 217010 303793
rect 216954 303719 217010 303728
rect 216862 302832 216918 302841
rect 216862 302767 216918 302776
rect 217046 301064 217102 301073
rect 217046 300999 217102 301008
rect 216770 299432 216826 299441
rect 216770 299367 216826 299376
rect 216680 280152 216732 280158
rect 216680 280094 216732 280100
rect 216692 279993 216720 280094
rect 216678 279984 216734 279993
rect 216678 279919 216734 279928
rect 216680 278724 216732 278730
rect 216680 278666 216732 278672
rect 216692 278089 216720 278666
rect 216954 278352 217010 278361
rect 216954 278287 216956 278296
rect 217008 278287 217010 278296
rect 216956 278258 217008 278264
rect 216678 278080 216734 278089
rect 216678 278015 216734 278024
rect 216956 269000 217008 269006
rect 216956 268942 217008 268948
rect 216968 268841 216996 268942
rect 216954 268832 217010 268841
rect 216954 268767 217010 268776
rect 216956 266212 217008 266218
rect 216956 266154 217008 266160
rect 216588 265668 216640 265674
rect 216588 265610 216640 265616
rect 216678 201920 216734 201929
rect 216678 201855 216734 201864
rect 216692 174026 216720 201855
rect 216770 201376 216826 201385
rect 216770 201311 216826 201320
rect 216600 173998 216720 174026
rect 216600 173210 216628 173998
rect 216680 173868 216732 173874
rect 216680 173810 216732 173816
rect 216692 173369 216720 173810
rect 216678 173360 216734 173369
rect 216678 173295 216734 173304
rect 216600 173182 216720 173210
rect 216588 145648 216640 145654
rect 216588 145590 216640 145596
rect 216600 144838 216628 145590
rect 216588 144832 216640 144838
rect 216588 144774 216640 144780
rect 216692 96937 216720 173182
rect 216678 96928 216734 96937
rect 216678 96863 216734 96872
rect 216784 95985 216812 201311
rect 216862 197432 216918 197441
rect 216862 197367 216918 197376
rect 216770 95976 216826 95985
rect 216770 95911 216826 95920
rect 216876 92857 216904 197367
rect 216968 147674 216996 266154
rect 217060 196081 217088 300999
rect 217152 265810 217180 370262
rect 217244 299985 217272 375022
rect 217336 375018 217364 383454
rect 217324 375012 217376 375018
rect 217324 374954 217376 374960
rect 217336 301073 217364 374954
rect 217428 370530 217456 477414
rect 217520 371006 217548 478246
rect 217796 477737 217824 480037
rect 218164 480023 218270 480051
rect 218440 480023 218730 480051
rect 218808 480023 219190 480051
rect 217782 477728 217838 477737
rect 217782 477663 217838 477672
rect 218060 475380 218112 475386
rect 218060 475322 218112 475328
rect 217692 471300 217744 471306
rect 217692 471242 217744 471248
rect 217600 463616 217652 463622
rect 217600 463558 217652 463564
rect 217612 374202 217640 463558
rect 217704 404297 217732 471242
rect 217784 467152 217836 467158
rect 217784 467094 217836 467100
rect 217796 410961 217824 467094
rect 217876 457496 217928 457502
rect 217876 457438 217928 457444
rect 217782 410952 217838 410961
rect 217782 410887 217838 410896
rect 217796 410009 217824 410887
rect 217782 410000 217838 410009
rect 217782 409935 217838 409944
rect 217888 404977 217916 457438
rect 217966 411904 218022 411913
rect 217966 411839 218022 411848
rect 217980 411369 218008 411839
rect 217966 411360 218022 411369
rect 217966 411295 218022 411304
rect 217874 404968 217930 404977
rect 217796 404926 217874 404954
rect 217690 404288 217746 404297
rect 217690 404223 217746 404232
rect 217796 375358 217824 404926
rect 217874 404903 217930 404912
rect 217874 404288 217930 404297
rect 217874 404223 217930 404232
rect 217888 403209 217916 404223
rect 217874 403200 217930 403209
rect 217874 403135 217930 403144
rect 217784 375352 217836 375358
rect 217888 375329 217916 403135
rect 217784 375294 217836 375300
rect 217874 375320 217930 375329
rect 217874 375255 217930 375264
rect 217600 374196 217652 374202
rect 217600 374138 217652 374144
rect 217784 373108 217836 373114
rect 217784 373050 217836 373056
rect 217796 372842 217824 373050
rect 217692 372836 217744 372842
rect 217692 372778 217744 372784
rect 217784 372836 217836 372842
rect 217784 372778 217836 372784
rect 217508 371000 217560 371006
rect 217508 370942 217560 370948
rect 217416 370524 217468 370530
rect 217416 370466 217468 370472
rect 217704 305969 217732 372778
rect 217876 353456 217928 353462
rect 217876 353398 217928 353404
rect 217782 307728 217838 307737
rect 217782 307663 217838 307672
rect 217796 306921 217824 307663
rect 217782 306912 217838 306921
rect 217782 306847 217838 306856
rect 217690 305960 217746 305969
rect 217690 305895 217746 305904
rect 217414 303784 217470 303793
rect 217414 303719 217470 303728
rect 217322 301064 217378 301073
rect 217322 300999 217378 301008
rect 217230 299976 217286 299985
rect 217230 299911 217286 299920
rect 217140 265804 217192 265810
rect 217140 265746 217192 265752
rect 217140 264308 217192 264314
rect 217140 264250 217192 264256
rect 217046 196072 217102 196081
rect 217046 196007 217102 196016
rect 217048 173800 217100 173806
rect 217048 173742 217100 173748
rect 217060 173097 217088 173742
rect 217046 173088 217102 173097
rect 217046 173023 217102 173032
rect 217152 162994 217180 264250
rect 217244 194993 217272 299911
rect 217428 198801 217456 303719
rect 217506 302832 217562 302841
rect 217506 302767 217562 302776
rect 217414 198792 217470 198801
rect 217414 198727 217470 198736
rect 217520 197849 217548 302767
rect 217598 299432 217654 299441
rect 217598 299367 217654 299376
rect 217612 298217 217640 299367
rect 217598 298208 217654 298217
rect 217598 298143 217654 298152
rect 217506 197840 217562 197849
rect 217506 197775 217562 197784
rect 217520 197441 217548 197775
rect 217506 197432 217562 197441
rect 217506 197367 217562 197376
rect 217230 194984 217286 194993
rect 217230 194919 217286 194928
rect 217140 162988 217192 162994
rect 217140 162930 217192 162936
rect 217152 156670 217180 162930
rect 217140 156664 217192 156670
rect 217140 156606 217192 156612
rect 216968 147646 217180 147674
rect 217152 145178 217180 147646
rect 217140 145172 217192 145178
rect 217140 145114 217192 145120
rect 217048 144968 217100 144974
rect 217048 144910 217100 144916
rect 216862 92848 216918 92857
rect 216862 92783 216918 92792
rect 216680 70372 216732 70378
rect 216680 70314 216732 70320
rect 216692 70009 216720 70314
rect 216678 70000 216734 70009
rect 216678 69935 216734 69944
rect 216678 68368 216734 68377
rect 216678 68303 216734 68312
rect 216692 67658 216720 68303
rect 216680 67652 216732 67658
rect 216680 67594 216732 67600
rect 216496 57656 216548 57662
rect 216496 57598 216548 57604
rect 216220 55208 216272 55214
rect 216220 55150 216272 55156
rect 216128 55072 216180 55078
rect 216128 55014 216180 55020
rect 217060 54738 217088 144910
rect 217152 54806 217180 145114
rect 217244 90001 217272 194919
rect 217612 193225 217640 298143
rect 217704 201385 217732 305895
rect 217796 201929 217824 306847
rect 217888 265849 217916 353398
rect 217980 307737 218008 411295
rect 218072 378826 218100 475322
rect 218060 378820 218112 378826
rect 218060 378762 218112 378768
rect 218060 374264 218112 374270
rect 218060 374206 218112 374212
rect 218072 374066 218100 374206
rect 218060 374060 218112 374066
rect 218060 374002 218112 374008
rect 218164 371521 218192 480023
rect 218440 470594 218468 480023
rect 218808 475386 218836 480023
rect 218796 475380 218848 475386
rect 218796 475322 218848 475328
rect 219440 475380 219492 475386
rect 219440 475322 219492 475328
rect 218704 472660 218756 472666
rect 218704 472602 218756 472608
rect 218256 470566 218468 470594
rect 218256 374241 218284 470566
rect 218612 459604 218664 459610
rect 218612 459546 218664 459552
rect 218336 378820 218388 378826
rect 218336 378762 218388 378768
rect 218242 374232 218298 374241
rect 218242 374167 218298 374176
rect 218348 371657 218376 378762
rect 218624 372473 218652 459546
rect 218610 372464 218666 372473
rect 218610 372399 218666 372408
rect 218334 371648 218390 371657
rect 218334 371583 218390 371592
rect 218150 371512 218206 371521
rect 218150 371447 218206 371456
rect 218612 353388 218664 353394
rect 218612 353330 218664 353336
rect 217966 307728 218022 307737
rect 217966 307663 218022 307672
rect 217966 268016 218022 268025
rect 217966 267951 218022 267960
rect 217980 267850 218008 267951
rect 217968 267844 218020 267850
rect 217968 267786 218020 267792
rect 218426 266928 218482 266937
rect 218426 266863 218482 266872
rect 217968 266008 218020 266014
rect 217968 265950 218020 265956
rect 217874 265840 217930 265849
rect 217874 265775 217930 265784
rect 217888 265033 217916 265775
rect 217874 265024 217930 265033
rect 217874 264959 217930 264968
rect 217782 201920 217838 201929
rect 217782 201855 217838 201864
rect 217690 201376 217746 201385
rect 217690 201311 217746 201320
rect 217704 200977 217732 201311
rect 217690 200968 217746 200977
rect 217690 200903 217746 200912
rect 217782 198792 217838 198801
rect 217782 198727 217838 198736
rect 217690 196072 217746 196081
rect 217690 196007 217746 196016
rect 217598 193216 217654 193225
rect 217598 193151 217654 193160
rect 217230 89992 217286 90001
rect 217230 89927 217286 89936
rect 217612 88233 217640 193151
rect 217704 91089 217732 196007
rect 217796 93809 217824 198727
rect 217874 161120 217930 161129
rect 217874 161055 217876 161064
rect 217928 161055 217930 161064
rect 217876 161026 217928 161032
rect 217876 156664 217928 156670
rect 217876 156606 217928 156612
rect 217782 93800 217838 93809
rect 217782 93735 217838 93744
rect 217690 91080 217746 91089
rect 217690 91015 217746 91024
rect 217598 88224 217654 88233
rect 217598 88159 217654 88168
rect 217888 59566 217916 156606
rect 217980 145926 218008 265950
rect 218334 163704 218390 163713
rect 218334 163639 218390 163648
rect 218244 160132 218296 160138
rect 218244 160074 218296 160080
rect 217968 145920 218020 145926
rect 217968 145862 218020 145868
rect 217980 144974 218008 145862
rect 217968 144968 218020 144974
rect 217968 144910 218020 144916
rect 217966 68368 218022 68377
rect 217966 68303 218022 68312
rect 217876 59560 217928 59566
rect 217876 59502 217928 59508
rect 217980 59362 218008 68303
rect 217968 59356 218020 59362
rect 217968 59298 218020 59304
rect 218256 56234 218284 160074
rect 218348 57458 218376 163639
rect 218440 147674 218468 266863
rect 218624 265878 218652 353330
rect 218612 265872 218664 265878
rect 218612 265814 218664 265820
rect 218612 265668 218664 265674
rect 218612 265610 218664 265616
rect 218520 249824 218572 249830
rect 218520 249766 218572 249772
rect 218532 161362 218560 249766
rect 218624 163470 218652 265610
rect 218612 163464 218664 163470
rect 218612 163406 218664 163412
rect 218520 161356 218572 161362
rect 218520 161298 218572 161304
rect 218532 160138 218560 161298
rect 218520 160132 218572 160138
rect 218520 160074 218572 160080
rect 218440 147646 218652 147674
rect 218624 145450 218652 147646
rect 218612 145444 218664 145450
rect 218612 145386 218664 145392
rect 218520 145104 218572 145110
rect 218520 145046 218572 145052
rect 218532 59634 218560 145046
rect 218624 59702 218652 145386
rect 218716 61010 218744 472602
rect 218796 468648 218848 468654
rect 218796 468590 218848 468596
rect 218808 162654 218836 468590
rect 218980 460828 219032 460834
rect 218980 460770 219032 460776
rect 218886 458960 218942 458969
rect 218886 458895 218942 458904
rect 218796 162648 218848 162654
rect 218796 162590 218848 162596
rect 218900 162382 218928 458895
rect 218992 267306 219020 460770
rect 219164 460488 219216 460494
rect 219164 460430 219216 460436
rect 219072 374060 219124 374066
rect 219072 374002 219124 374008
rect 218980 267300 219032 267306
rect 218980 267242 219032 267248
rect 218980 265804 219032 265810
rect 218980 265746 219032 265752
rect 218888 162376 218940 162382
rect 218888 162318 218940 162324
rect 218992 161158 219020 265746
rect 219084 264586 219112 374002
rect 219176 369306 219204 460430
rect 219348 374264 219400 374270
rect 219348 374206 219400 374212
rect 219360 373862 219388 374206
rect 219348 373856 219400 373862
rect 219348 373798 219400 373804
rect 219256 373652 219308 373658
rect 219256 373594 219308 373600
rect 219268 372706 219296 373594
rect 219256 372700 219308 372706
rect 219256 372642 219308 372648
rect 219164 369300 219216 369306
rect 219164 369242 219216 369248
rect 219164 353320 219216 353326
rect 219164 353262 219216 353268
rect 219176 266218 219204 353262
rect 219268 266937 219296 372642
rect 219254 266928 219310 266937
rect 219254 266863 219310 266872
rect 219164 266212 219216 266218
rect 219164 266154 219216 266160
rect 219256 266144 219308 266150
rect 219256 266086 219308 266092
rect 219164 265940 219216 265946
rect 219164 265882 219216 265888
rect 219072 264580 219124 264586
rect 219072 264522 219124 264528
rect 219072 250572 219124 250578
rect 219072 250514 219124 250520
rect 218980 161152 219032 161158
rect 218980 161094 219032 161100
rect 219084 146266 219112 250514
rect 219072 146260 219124 146266
rect 219072 146202 219124 146208
rect 218980 145376 219032 145382
rect 218980 145318 219032 145324
rect 218796 145036 218848 145042
rect 218796 144978 218848 144984
rect 218808 61130 218836 144978
rect 218888 144968 218940 144974
rect 218888 144910 218940 144916
rect 218796 61124 218848 61130
rect 218796 61066 218848 61072
rect 218716 60982 218836 61010
rect 218702 60616 218758 60625
rect 218702 60551 218758 60560
rect 218612 59696 218664 59702
rect 218612 59638 218664 59644
rect 218520 59628 218572 59634
rect 218520 59570 218572 59576
rect 218716 57798 218744 60551
rect 218704 57792 218756 57798
rect 218704 57734 218756 57740
rect 218336 57452 218388 57458
rect 218336 57394 218388 57400
rect 218808 57254 218836 60982
rect 218796 57248 218848 57254
rect 218796 57190 218848 57196
rect 218244 56228 218296 56234
rect 218244 56170 218296 56176
rect 218900 56098 218928 144910
rect 218992 56438 219020 145318
rect 219084 145110 219112 146202
rect 219176 145858 219204 265882
rect 219268 145994 219296 266086
rect 219360 265742 219388 373798
rect 219452 371385 219480 475322
rect 219544 372570 219572 480037
rect 219636 480023 220018 480051
rect 220096 480023 220478 480051
rect 220832 480023 220938 480051
rect 221016 480023 221398 480051
rect 219636 374105 219664 480023
rect 219716 477556 219768 477562
rect 219716 477498 219768 477504
rect 219992 477556 220044 477562
rect 219992 477498 220044 477504
rect 219622 374096 219678 374105
rect 219622 374031 219678 374040
rect 219532 372564 219584 372570
rect 219532 372506 219584 372512
rect 219532 372088 219584 372094
rect 219532 372030 219584 372036
rect 219438 371376 219494 371385
rect 219438 371311 219494 371320
rect 219544 265946 219572 372030
rect 219624 372020 219676 372026
rect 219624 371962 219676 371968
rect 219636 266150 219664 371962
rect 219728 368490 219756 477498
rect 219808 373312 219860 373318
rect 219808 373254 219860 373260
rect 219716 368484 219768 368490
rect 219716 368426 219768 368432
rect 219624 266144 219676 266150
rect 219624 266086 219676 266092
rect 219532 265940 219584 265946
rect 219532 265882 219584 265888
rect 219348 265736 219400 265742
rect 219348 265678 219400 265684
rect 219624 265736 219676 265742
rect 219624 265678 219676 265684
rect 219532 250504 219584 250510
rect 219532 250446 219584 250452
rect 219544 161430 219572 250446
rect 219532 161424 219584 161430
rect 219532 161366 219584 161372
rect 219348 161152 219400 161158
rect 219348 161094 219400 161100
rect 219256 145988 219308 145994
rect 219256 145930 219308 145936
rect 219164 145852 219216 145858
rect 219164 145794 219216 145800
rect 219072 145104 219124 145110
rect 219072 145046 219124 145052
rect 219072 61124 219124 61130
rect 219072 61066 219124 61072
rect 218980 56432 219032 56438
rect 218980 56374 219032 56380
rect 219084 56166 219112 61066
rect 219072 56160 219124 56166
rect 219072 56102 219124 56108
rect 218888 56092 218940 56098
rect 218888 56034 218940 56040
rect 219176 56030 219204 145794
rect 219268 144974 219296 145930
rect 219256 144968 219308 144974
rect 219256 144910 219308 144916
rect 219254 60616 219310 60625
rect 219254 60551 219310 60560
rect 219268 58682 219296 60551
rect 219360 59498 219388 161094
rect 219348 59492 219400 59498
rect 219348 59434 219400 59440
rect 219256 58676 219308 58682
rect 219256 58618 219308 58624
rect 219544 56302 219572 161366
rect 219636 161226 219664 265678
rect 219820 264790 219848 373254
rect 219900 371340 219952 371346
rect 219900 371282 219952 371288
rect 219912 266014 219940 371282
rect 219900 266008 219952 266014
rect 219900 265950 219952 265956
rect 219900 265872 219952 265878
rect 219900 265814 219952 265820
rect 219808 264784 219860 264790
rect 219808 264726 219860 264732
rect 219716 163464 219768 163470
rect 219716 163406 219768 163412
rect 219624 161220 219676 161226
rect 219624 161162 219676 161168
rect 219532 56296 219584 56302
rect 219532 56238 219584 56244
rect 219164 56024 219216 56030
rect 219164 55966 219216 55972
rect 219636 54942 219664 161162
rect 219728 55010 219756 163406
rect 219820 146130 219848 264726
rect 219808 146124 219860 146130
rect 219808 146066 219860 146072
rect 219716 55004 219768 55010
rect 219716 54946 219768 54952
rect 219624 54936 219676 54942
rect 219624 54878 219676 54884
rect 219820 54874 219848 146066
rect 219912 146062 219940 265814
rect 219900 146056 219952 146062
rect 219900 145998 219952 146004
rect 219912 145042 219940 145998
rect 219900 145036 219952 145042
rect 219900 144978 219952 144984
rect 220004 55826 220032 477498
rect 220096 475386 220124 480023
rect 220084 475380 220136 475386
rect 220084 475322 220136 475328
rect 220832 475250 220860 480023
rect 221016 475538 221044 480023
rect 221752 478242 221780 480037
rect 221740 478236 221792 478242
rect 221740 478178 221792 478184
rect 222212 476785 222240 480037
rect 222672 477562 222700 480037
rect 223132 477601 223160 480037
rect 223606 480023 223636 480051
rect 223608 479874 223636 480023
rect 223684 480023 223974 480051
rect 223596 479868 223648 479874
rect 223596 479810 223648 479816
rect 223118 477592 223174 477601
rect 222660 477556 222712 477562
rect 223118 477527 223174 477536
rect 222660 477498 222712 477504
rect 222198 476776 222254 476785
rect 222198 476711 222254 476720
rect 220924 475510 221044 475538
rect 220820 475244 220872 475250
rect 220820 475186 220872 475192
rect 220924 459678 220952 475510
rect 223580 475380 223632 475386
rect 223580 475322 223632 475328
rect 221004 475244 221056 475250
rect 221004 475186 221056 475192
rect 220912 459672 220964 459678
rect 220912 459614 220964 459620
rect 221016 459610 221044 475186
rect 221004 459604 221056 459610
rect 221004 459546 221056 459552
rect 223592 458833 223620 475322
rect 223684 467158 223712 480023
rect 223764 479868 223816 479874
rect 223764 479810 223816 479816
rect 223672 467152 223724 467158
rect 223672 467094 223724 467100
rect 223776 458969 223804 479810
rect 224420 478310 224448 480037
rect 224512 480023 224894 480051
rect 224408 478304 224460 478310
rect 224408 478246 224460 478252
rect 224512 475386 224540 480023
rect 225340 478174 225368 480037
rect 225708 478242 225736 480037
rect 226168 478281 226196 480037
rect 226444 480023 226642 480051
rect 226720 480023 227102 480051
rect 226154 478272 226210 478281
rect 225696 478236 225748 478242
rect 226154 478207 226210 478216
rect 225696 478178 225748 478184
rect 225328 478168 225380 478174
rect 225328 478110 225380 478116
rect 224500 475380 224552 475386
rect 224500 475322 224552 475328
rect 226340 475380 226392 475386
rect 226340 475322 226392 475328
rect 226352 465730 226380 475322
rect 226444 468518 226472 480023
rect 226720 475386 226748 480023
rect 226708 475380 226760 475386
rect 226708 475322 226760 475328
rect 227548 472666 227576 480037
rect 227720 475380 227772 475386
rect 227720 475322 227772 475328
rect 227536 472660 227588 472666
rect 227536 472602 227588 472608
rect 227732 468586 227760 475322
rect 227916 471306 227944 480037
rect 228008 480023 228390 480051
rect 228560 480023 228850 480051
rect 229204 480023 229310 480051
rect 229480 480023 229770 480051
rect 229848 480023 230138 480051
rect 227904 471300 227956 471306
rect 227904 471242 227956 471248
rect 228008 470594 228036 480023
rect 228560 475386 228588 480023
rect 228548 475380 228600 475386
rect 228548 475322 228600 475328
rect 229100 475380 229152 475386
rect 229100 475322 229152 475328
rect 227824 470566 228036 470594
rect 227824 469946 227852 470566
rect 227812 469940 227864 469946
rect 227812 469882 227864 469888
rect 227720 468580 227772 468586
rect 227720 468522 227772 468528
rect 226432 468512 226484 468518
rect 226432 468454 226484 468460
rect 229112 465769 229140 475322
rect 229204 467226 229232 480023
rect 229480 475386 229508 480023
rect 229468 475380 229520 475386
rect 229468 475322 229520 475328
rect 229848 470594 229876 480023
rect 230584 478553 230612 480037
rect 230768 480023 231058 480051
rect 230570 478544 230626 478553
rect 230570 478479 230626 478488
rect 230768 470594 230796 480023
rect 231504 478417 231532 480037
rect 231490 478408 231546 478417
rect 231490 478343 231546 478352
rect 231872 475561 231900 480037
rect 232332 478145 232360 480037
rect 232792 478378 232820 480037
rect 232780 478372 232832 478378
rect 232780 478314 232832 478320
rect 232318 478136 232374 478145
rect 232318 478071 232374 478080
rect 231858 475552 231914 475561
rect 231858 475487 231914 475496
rect 233252 474201 233280 480037
rect 233712 478281 233740 480037
rect 233698 478272 233754 478281
rect 233698 478207 233754 478216
rect 233238 474192 233294 474201
rect 233238 474127 233294 474136
rect 234080 471209 234108 480037
rect 234540 478009 234568 480037
rect 234526 478000 234582 478009
rect 234526 477935 234582 477944
rect 235000 472802 235028 480037
rect 235460 478689 235488 480037
rect 235920 478825 235948 480037
rect 236288 478854 236316 480037
rect 236472 480023 236762 480051
rect 236276 478848 236328 478854
rect 235906 478816 235962 478825
rect 236276 478790 236328 478796
rect 235906 478751 235962 478760
rect 235446 478680 235502 478689
rect 235446 478615 235502 478624
rect 234988 472796 235040 472802
rect 234988 472738 235040 472744
rect 234066 471200 234122 471209
rect 234066 471135 234122 471144
rect 236472 470594 236500 480023
rect 237208 474026 237236 480037
rect 237196 474020 237248 474026
rect 237196 473962 237248 473968
rect 237668 471442 237696 480037
rect 238128 475454 238156 480037
rect 238220 480023 238510 480051
rect 238116 475448 238168 475454
rect 238116 475390 238168 475396
rect 237656 471436 237708 471442
rect 237656 471378 237708 471384
rect 238220 470594 238248 480023
rect 238956 472734 238984 480037
rect 239416 478582 239444 480037
rect 239404 478576 239456 478582
rect 239404 478518 239456 478524
rect 239876 478446 239904 480037
rect 240244 478514 240272 480037
rect 240336 480023 240718 480051
rect 240888 480023 241178 480051
rect 241532 480023 241638 480051
rect 240232 478508 240284 478514
rect 240232 478450 240284 478456
rect 239864 478440 239916 478446
rect 239864 478382 239916 478388
rect 240140 475380 240192 475386
rect 240140 475322 240192 475328
rect 238944 472728 238996 472734
rect 238944 472670 238996 472676
rect 229296 470566 229876 470594
rect 230492 470566 230796 470594
rect 236012 470566 236500 470594
rect 237392 470566 238248 470594
rect 229296 469878 229324 470566
rect 229284 469872 229336 469878
rect 229284 469814 229336 469820
rect 230492 468489 230520 470566
rect 236012 470014 236040 470566
rect 236000 470008 236052 470014
rect 236000 469950 236052 469956
rect 230478 468480 230534 468489
rect 230478 468415 230534 468424
rect 229192 467220 229244 467226
rect 229192 467162 229244 467168
rect 229098 465760 229154 465769
rect 226340 465724 226392 465730
rect 229098 465695 229154 465704
rect 226340 465666 226392 465672
rect 237392 460222 237420 470566
rect 240152 463010 240180 475322
rect 240336 470594 240364 480023
rect 240888 475386 240916 480023
rect 240876 475380 240928 475386
rect 240876 475322 240928 475328
rect 240244 470566 240364 470594
rect 240244 465798 240272 470566
rect 241532 468654 241560 480023
rect 242084 475250 242112 480037
rect 242072 475244 242124 475250
rect 242072 475186 242124 475192
rect 242452 472938 242480 480037
rect 242912 476882 242940 480037
rect 243004 480023 243386 480051
rect 243464 480023 243846 480051
rect 244306 480023 244504 480051
rect 242900 476876 242952 476882
rect 242900 476818 242952 476824
rect 243004 475300 243032 480023
rect 242912 475272 243032 475300
rect 242440 472932 242492 472938
rect 242440 472874 242492 472880
rect 241520 468648 241572 468654
rect 241520 468590 241572 468596
rect 240232 465792 240284 465798
rect 240232 465734 240284 465740
rect 240140 463004 240192 463010
rect 240140 462946 240192 462952
rect 237380 460216 237432 460222
rect 237380 460158 237432 460164
rect 223762 458960 223818 458969
rect 242912 458930 242940 475272
rect 243464 470594 243492 480023
rect 244280 475380 244332 475386
rect 244280 475322 244332 475328
rect 243004 470566 243492 470594
rect 243004 467294 243032 470566
rect 242992 467288 243044 467294
rect 242992 467230 243044 467236
rect 244292 460426 244320 475322
rect 244372 475312 244424 475318
rect 244372 475254 244424 475260
rect 244384 468722 244412 475254
rect 244476 470082 244504 480023
rect 244568 480023 244674 480051
rect 244752 480023 245134 480051
rect 244568 475318 244596 480023
rect 244752 475386 244780 480023
rect 244740 475380 244792 475386
rect 244740 475322 244792 475328
rect 244556 475312 244608 475318
rect 244556 475254 244608 475260
rect 245580 472870 245608 480037
rect 246040 474094 246068 480037
rect 246408 475522 246436 480037
rect 246396 475516 246448 475522
rect 246396 475458 246448 475464
rect 246028 474088 246080 474094
rect 246028 474030 246080 474036
rect 245568 472864 245620 472870
rect 245568 472806 245620 472812
rect 246868 471374 246896 480037
rect 247236 480023 247342 480051
rect 247512 480023 247802 480051
rect 247880 480023 248262 480051
rect 247132 475380 247184 475386
rect 247132 475322 247184 475328
rect 247040 475312 247092 475318
rect 247040 475254 247092 475260
rect 246856 471368 246908 471374
rect 246856 471310 246908 471316
rect 244464 470076 244516 470082
rect 244464 470018 244516 470024
rect 244372 468716 244424 468722
rect 244372 468658 244424 468664
rect 244280 460420 244332 460426
rect 244280 460362 244332 460368
rect 223762 458895 223818 458904
rect 242900 458924 242952 458930
rect 242900 458866 242952 458872
rect 247052 458862 247080 475254
rect 247144 460290 247172 475322
rect 247236 460358 247264 480023
rect 247512 475386 247540 480023
rect 247500 475380 247552 475386
rect 247500 475322 247552 475328
rect 247880 475318 247908 480023
rect 248788 480072 248840 480078
rect 248420 480014 248472 480020
rect 247868 475312 247920 475318
rect 247868 475254 247920 475260
rect 248432 460562 248460 480014
rect 248616 475538 248644 480037
rect 248840 480023 249090 480051
rect 249168 480023 249550 480051
rect 249812 480023 250010 480051
rect 250088 480023 250470 480051
rect 250548 480023 250838 480051
rect 251192 480023 251298 480051
rect 251376 480023 251758 480051
rect 248788 480014 248840 480020
rect 248616 475510 248736 475538
rect 248512 475312 248564 475318
rect 248512 475254 248564 475260
rect 248420 460556 248472 460562
rect 248420 460498 248472 460504
rect 248524 460494 248552 475254
rect 248708 470594 248736 475510
rect 249168 475318 249196 480023
rect 249156 475312 249208 475318
rect 249156 475254 249208 475260
rect 248616 470566 248736 470594
rect 248616 460630 248644 470566
rect 249812 463078 249840 480023
rect 250088 475402 250116 480023
rect 249904 475374 250116 475402
rect 249904 463146 249932 475374
rect 250548 470594 250576 480023
rect 249996 470566 250576 470594
rect 249996 465934 250024 470566
rect 249984 465928 250036 465934
rect 249984 465870 250036 465876
rect 251192 465866 251220 480023
rect 251376 470594 251404 480023
rect 252204 471578 252232 480037
rect 252586 480023 252616 480051
rect 252588 479890 252616 480023
rect 252848 480023 253046 480051
rect 253124 480023 253506 480051
rect 252588 479862 252784 479890
rect 252756 474337 252784 479862
rect 252742 474328 252798 474337
rect 252742 474263 252798 474272
rect 252848 474178 252876 480023
rect 252572 474150 252876 474178
rect 252192 471572 252244 471578
rect 252192 471514 252244 471520
rect 251284 470566 251404 470594
rect 251284 468790 251312 470566
rect 251272 468784 251324 468790
rect 251272 468726 251324 468732
rect 251180 465860 251232 465866
rect 251180 465802 251232 465808
rect 249892 463140 249944 463146
rect 249892 463082 249944 463088
rect 249800 463072 249852 463078
rect 249800 463014 249852 463020
rect 252572 461718 252600 474150
rect 253124 470594 253152 480023
rect 252664 470566 253152 470594
rect 252560 461712 252612 461718
rect 252560 461654 252612 461660
rect 252664 461650 252692 470566
rect 253952 461854 253980 480037
rect 254412 474298 254440 480037
rect 254780 477290 254808 480037
rect 254768 477284 254820 477290
rect 254768 477226 254820 477232
rect 255240 476921 255268 480037
rect 255700 477154 255728 480037
rect 255688 477148 255740 477154
rect 255688 477090 255740 477096
rect 255226 476912 255282 476921
rect 255226 476847 255282 476856
rect 254400 474292 254452 474298
rect 254400 474234 254452 474240
rect 256160 472569 256188 480037
rect 256620 476950 256648 480037
rect 256712 480023 257002 480051
rect 257080 480023 257462 480051
rect 257540 480023 257922 480051
rect 256608 476944 256660 476950
rect 256608 476886 256660 476892
rect 256146 472560 256202 472569
rect 256146 472495 256202 472504
rect 256712 467430 256740 480023
rect 257080 475402 257108 480023
rect 256804 475374 257108 475402
rect 256804 468858 256832 475374
rect 257540 470594 257568 480023
rect 258080 472116 258132 472122
rect 258080 472058 258132 472064
rect 256896 470566 257568 470594
rect 256896 470150 256924 470566
rect 256884 470144 256936 470150
rect 256884 470086 256936 470092
rect 256792 468852 256844 468858
rect 256792 468794 256844 468800
rect 256700 467424 256752 467430
rect 256700 467366 256752 467372
rect 253940 461848 253992 461854
rect 253940 461790 253992 461796
rect 252652 461644 252704 461650
rect 252652 461586 252704 461592
rect 248604 460624 248656 460630
rect 248604 460566 248656 460572
rect 248512 460488 248564 460494
rect 248512 460430 248564 460436
rect 247224 460352 247276 460358
rect 247224 460294 247276 460300
rect 247132 460284 247184 460290
rect 247132 460226 247184 460232
rect 258092 458998 258120 472058
rect 258368 471782 258396 480037
rect 258460 480023 258842 480051
rect 258920 480023 259210 480051
rect 259472 480023 259670 480051
rect 258356 471776 258408 471782
rect 258356 471718 258408 471724
rect 258460 470594 258488 480023
rect 258920 472122 258948 480023
rect 258908 472116 258960 472122
rect 258908 472058 258960 472064
rect 258184 470566 258488 470594
rect 258184 460766 258212 470566
rect 259472 468926 259500 480023
rect 260116 474162 260144 480037
rect 260576 477018 260604 480037
rect 260564 477012 260616 477018
rect 260564 476954 260616 476960
rect 260944 475590 260972 480037
rect 261036 480023 261418 480051
rect 260932 475584 260984 475590
rect 260932 475526 260984 475532
rect 260104 474156 260156 474162
rect 260104 474098 260156 474104
rect 261036 470594 261064 480023
rect 261864 473006 261892 480037
rect 262220 475312 262272 475318
rect 262220 475254 262272 475260
rect 261852 473000 261904 473006
rect 261852 472942 261904 472948
rect 260852 470566 261064 470594
rect 259460 468920 259512 468926
rect 259460 468862 259512 468868
rect 260852 461786 260880 470566
rect 260840 461780 260892 461786
rect 260840 461722 260892 461728
rect 262232 460834 262260 475254
rect 262324 467362 262352 480037
rect 262416 480023 262798 480051
rect 262416 475318 262444 480023
rect 262404 475312 262456 475318
rect 262404 475254 262456 475260
rect 263152 471510 263180 480037
rect 263626 480023 263656 480051
rect 263628 479890 263656 480023
rect 263888 480023 264086 480051
rect 264256 480023 264546 480051
rect 265006 480023 265296 480051
rect 263628 479862 263824 479890
rect 263600 475312 263652 475318
rect 263600 475254 263652 475260
rect 263140 471504 263192 471510
rect 263140 471446 263192 471452
rect 262312 467356 262364 467362
rect 262312 467298 262364 467304
rect 262220 460828 262272 460834
rect 262220 460770 262272 460776
rect 258172 460760 258224 460766
rect 258172 460702 258224 460708
rect 263612 459066 263640 475254
rect 263796 471850 263824 479862
rect 263784 471844 263836 471850
rect 263784 471786 263836 471792
rect 263888 470594 263916 480023
rect 264256 475318 264284 480023
rect 264244 475312 264296 475318
rect 264244 475254 264296 475260
rect 264980 475312 265032 475318
rect 264980 475254 265032 475260
rect 263704 470566 263916 470594
rect 263704 469849 263732 470566
rect 263690 469840 263746 469849
rect 263690 469775 263746 469784
rect 264992 469130 265020 475254
rect 265268 474366 265296 480023
rect 265256 474360 265308 474366
rect 265256 474302 265308 474308
rect 265360 474230 265388 480037
rect 265452 480023 265834 480051
rect 265912 480023 266294 480051
rect 266372 480023 266754 480051
rect 266832 480023 267122 480051
rect 265348 474224 265400 474230
rect 265348 474166 265400 474172
rect 265452 470594 265480 480023
rect 265912 475318 265940 480023
rect 265900 475312 265952 475318
rect 265900 475254 265952 475260
rect 265084 470566 265480 470594
rect 265084 470218 265112 470566
rect 265072 470212 265124 470218
rect 265072 470154 265124 470160
rect 264980 469124 265032 469130
rect 264980 469066 265032 469072
rect 266372 461553 266400 480023
rect 266832 470594 266860 480023
rect 267568 477222 267596 480037
rect 267752 480023 268042 480051
rect 268120 480023 268502 480051
rect 268672 480023 268962 480051
rect 267556 477216 267608 477222
rect 267556 477158 267608 477164
rect 266464 470566 266860 470594
rect 266464 467566 266492 470566
rect 266452 467560 266504 467566
rect 266452 467502 266504 467508
rect 266358 461544 266414 461553
rect 266358 461479 266414 461488
rect 267752 460698 267780 480023
rect 268120 475402 268148 480023
rect 267844 475374 268148 475402
rect 267844 463282 267872 475374
rect 268672 470594 268700 480023
rect 269316 471918 269344 480037
rect 269776 477086 269804 480037
rect 269764 477080 269816 477086
rect 269764 477022 269816 477028
rect 270236 475658 270264 480037
rect 270224 475652 270276 475658
rect 270224 475594 270276 475600
rect 269304 471912 269356 471918
rect 269304 471854 269356 471860
rect 270696 471646 270724 480037
rect 270880 480023 271170 480051
rect 270684 471640 270736 471646
rect 270684 471582 270736 471588
rect 270880 470594 270908 480023
rect 271524 475726 271552 480037
rect 271892 480023 271998 480051
rect 271512 475720 271564 475726
rect 271512 475662 271564 475668
rect 267936 470566 268700 470594
rect 270512 470566 270908 470594
rect 267936 467498 267964 470566
rect 270512 468994 270540 470566
rect 270500 468988 270552 468994
rect 270500 468930 270552 468936
rect 267924 467492 267976 467498
rect 267924 467434 267976 467440
rect 267832 463276 267884 463282
rect 267832 463218 267884 463224
rect 267740 460692 267792 460698
rect 267740 460634 267792 460640
rect 271892 459134 271920 480023
rect 272444 475794 272472 480037
rect 272432 475788 272484 475794
rect 272432 475730 272484 475736
rect 272904 474502 272932 480037
rect 272892 474496 272944 474502
rect 272892 474438 272944 474444
rect 273272 469062 273300 480037
rect 273732 471714 273760 480037
rect 274192 473074 274220 480037
rect 274180 473068 274232 473074
rect 274180 473010 274232 473016
rect 273720 471708 273772 471714
rect 273720 471650 273772 471656
rect 273260 469056 273312 469062
rect 273260 468998 273312 469004
rect 274652 467770 274680 480037
rect 274744 480023 275126 480051
rect 275204 480023 275494 480051
rect 274744 470354 274772 480023
rect 275204 470422 275232 480023
rect 275940 477358 275968 480037
rect 276032 480023 276414 480051
rect 276492 480023 276874 480051
rect 276952 480023 277334 480051
rect 277504 480023 277702 480051
rect 277872 480023 278162 480051
rect 278240 480023 278622 480051
rect 278884 480023 279082 480051
rect 279160 480023 279542 480051
rect 279620 480023 279910 480051
rect 280264 480023 280370 480051
rect 280448 480023 280830 480051
rect 280908 480023 281290 480051
rect 281552 480023 281658 480051
rect 275928 477352 275980 477358
rect 275928 477294 275980 477300
rect 275192 470416 275244 470422
rect 275192 470358 275244 470364
rect 274732 470348 274784 470354
rect 274732 470290 274784 470296
rect 274640 467764 274692 467770
rect 274640 467706 274692 467712
rect 276032 459202 276060 480023
rect 276492 476114 276520 480023
rect 276124 476086 276520 476114
rect 276124 463486 276152 476086
rect 276952 466454 276980 480023
rect 277400 471232 277452 471238
rect 277400 471174 277452 471180
rect 276216 466426 276980 466454
rect 276216 463554 276244 466426
rect 276204 463548 276256 463554
rect 276204 463490 276256 463496
rect 276112 463480 276164 463486
rect 276112 463422 276164 463428
rect 277412 461922 277440 471174
rect 277504 463622 277532 480023
rect 277872 471238 277900 480023
rect 277860 471232 277912 471238
rect 277860 471174 277912 471180
rect 278240 466454 278268 480023
rect 278780 471232 278832 471238
rect 278780 471174 278832 471180
rect 277596 466426 278268 466454
rect 277492 463616 277544 463622
rect 277492 463558 277544 463564
rect 277596 463350 277624 466426
rect 277584 463344 277636 463350
rect 277584 463286 277636 463292
rect 277400 461916 277452 461922
rect 277400 461858 277452 461864
rect 278792 460193 278820 471174
rect 278884 461990 278912 480023
rect 279160 471238 279188 480023
rect 279148 471232 279200 471238
rect 279148 471174 279200 471180
rect 279620 466454 279648 480023
rect 280264 471986 280292 480023
rect 280448 476114 280476 480023
rect 280356 476086 280476 476114
rect 280252 471980 280304 471986
rect 280252 471922 280304 471928
rect 280356 468058 280384 476086
rect 280436 471980 280488 471986
rect 280436 471922 280488 471928
rect 278976 466426 279648 466454
rect 280172 468030 280384 468058
rect 278976 463214 279004 466426
rect 278964 463208 279016 463214
rect 278964 463150 279016 463156
rect 278872 461984 278924 461990
rect 278872 461926 278924 461932
rect 278778 460184 278834 460193
rect 278778 460119 278834 460128
rect 280172 459270 280200 468030
rect 280448 463694 280476 471922
rect 280908 469198 280936 480023
rect 280896 469192 280948 469198
rect 280896 469134 280948 469140
rect 280264 463666 280476 463694
rect 280264 463418 280292 463666
rect 280252 463412 280304 463418
rect 280252 463354 280304 463360
rect 281552 459338 281580 480023
rect 282104 474434 282132 480037
rect 282564 474570 282592 480037
rect 283024 477494 283052 480037
rect 283208 480023 283498 480051
rect 283012 477488 283064 477494
rect 283012 477430 283064 477436
rect 282552 474564 282604 474570
rect 282552 474506 282604 474512
rect 282092 474428 282144 474434
rect 282092 474370 282144 474376
rect 283208 466454 283236 480023
rect 283852 475930 283880 480037
rect 283840 475924 283892 475930
rect 283840 475866 283892 475872
rect 282932 466426 283236 466454
rect 282932 462126 282960 466426
rect 284312 462942 284340 480037
rect 284772 473210 284800 480037
rect 284864 480023 285246 480051
rect 284760 473204 284812 473210
rect 284760 473146 284812 473152
rect 284864 466454 284892 480023
rect 284404 466426 284892 466454
rect 284404 464710 284432 466426
rect 284392 464704 284444 464710
rect 284392 464646 284444 464652
rect 285692 464642 285720 480037
rect 286060 470286 286088 480037
rect 286152 480023 286534 480051
rect 286704 480023 286994 480051
rect 286048 470280 286100 470286
rect 286048 470222 286100 470228
rect 285772 467628 285824 467634
rect 285772 467570 285824 467576
rect 285680 464636 285732 464642
rect 285680 464578 285732 464584
rect 285784 464370 285812 467570
rect 286152 466454 286180 480023
rect 286704 467634 286732 480023
rect 287060 471232 287112 471238
rect 287060 471174 287112 471180
rect 286692 467628 286744 467634
rect 286692 467570 286744 467576
rect 285876 466426 286180 466454
rect 285876 464438 285904 466426
rect 285864 464432 285916 464438
rect 285864 464374 285916 464380
rect 285772 464364 285824 464370
rect 285772 464306 285824 464312
rect 284300 462936 284352 462942
rect 284300 462878 284352 462884
rect 282920 462120 282972 462126
rect 282920 462062 282972 462068
rect 287072 460902 287100 471174
rect 287440 471170 287468 480037
rect 287532 480023 287822 480051
rect 287992 480023 288282 480051
rect 288452 480023 288742 480051
rect 288820 480023 289202 480051
rect 289280 480023 289662 480051
rect 289832 480023 290030 480051
rect 290200 480023 290490 480051
rect 290568 480023 290950 480051
rect 291212 480023 291410 480051
rect 291488 480023 291870 480051
rect 287428 471164 287480 471170
rect 287428 471106 287480 471112
rect 287532 466454 287560 480023
rect 287992 471238 288020 480023
rect 287980 471232 288032 471238
rect 287980 471174 288032 471180
rect 287164 466426 287560 466454
rect 287164 463690 287192 466426
rect 288452 464982 288480 480023
rect 288820 476114 288848 480023
rect 288544 476086 288848 476114
rect 288544 466002 288572 476086
rect 289280 466454 289308 480023
rect 288636 466426 289308 466454
rect 288636 466070 288664 466426
rect 289832 466138 289860 480023
rect 290200 467702 290228 480023
rect 290188 467696 290240 467702
rect 290188 467638 290240 467644
rect 290568 467634 290596 480023
rect 290556 467628 290608 467634
rect 290556 467570 290608 467576
rect 289820 466132 289872 466138
rect 289820 466074 289872 466080
rect 288624 466064 288676 466070
rect 288624 466006 288676 466012
rect 288532 465996 288584 466002
rect 288532 465938 288584 465944
rect 288440 464976 288492 464982
rect 288440 464918 288492 464924
rect 291212 464574 291240 480023
rect 291488 468450 291516 480023
rect 292224 471986 292252 480037
rect 292580 475312 292632 475318
rect 292580 475254 292632 475260
rect 292212 471980 292264 471986
rect 292212 471922 292264 471928
rect 291476 468444 291528 468450
rect 291476 468386 291528 468392
rect 292592 464778 292620 475254
rect 292684 464914 292712 480037
rect 292776 480023 293158 480051
rect 293328 480023 293618 480051
rect 292672 464908 292724 464914
rect 292672 464850 292724 464856
rect 292776 464846 292804 480023
rect 293328 475318 293356 480023
rect 293316 475312 293368 475318
rect 293316 475254 293368 475260
rect 292764 464840 292816 464846
rect 292764 464782 292816 464788
rect 292580 464772 292632 464778
rect 292580 464714 292632 464720
rect 291200 464568 291252 464574
rect 291200 464510 291252 464516
rect 293972 464506 294000 480037
rect 294432 477426 294460 480037
rect 294420 477420 294472 477426
rect 294420 477362 294472 477368
rect 294892 475862 294920 480037
rect 295366 480023 295396 480051
rect 295368 479874 295396 480023
rect 295444 480023 295826 480051
rect 295904 480023 296194 480051
rect 296272 480023 296654 480051
rect 295356 479868 295408 479874
rect 295356 479810 295408 479816
rect 294880 475856 294932 475862
rect 294880 475798 294932 475804
rect 295444 475538 295472 480023
rect 295352 475510 295472 475538
rect 293960 464500 294012 464506
rect 293960 464442 294012 464448
rect 287152 463684 287204 463690
rect 287152 463626 287204 463632
rect 287060 460896 287112 460902
rect 287060 460838 287112 460844
rect 295352 459474 295380 475510
rect 295904 475402 295932 480023
rect 295984 479868 296036 479874
rect 295984 479810 296036 479816
rect 295444 475374 295932 475402
rect 295444 460329 295472 475374
rect 295996 473142 296024 479810
rect 295984 473136 296036 473142
rect 295984 473078 296036 473084
rect 296272 470594 296300 480023
rect 296720 475312 296772 475318
rect 296720 475254 296772 475260
rect 295536 470566 296300 470594
rect 295536 462913 295564 470566
rect 295522 462904 295578 462913
rect 295522 462839 295578 462848
rect 296732 462058 296760 475254
rect 297100 474638 297128 480037
rect 297192 480023 297574 480051
rect 297744 480023 298034 480051
rect 298112 480023 298402 480051
rect 298480 480023 298862 480051
rect 298940 480023 299322 480051
rect 297088 474632 297140 474638
rect 297088 474574 297140 474580
rect 297192 470594 297220 480023
rect 297744 475318 297772 480023
rect 297732 475312 297784 475318
rect 297732 475254 297784 475260
rect 296824 470566 297220 470594
rect 296824 465905 296852 470566
rect 296810 465896 296866 465905
rect 296810 465831 296866 465840
rect 296720 462052 296772 462058
rect 296720 461994 296772 462000
rect 295430 460320 295486 460329
rect 295430 460255 295486 460264
rect 295340 459468 295392 459474
rect 295340 459410 295392 459416
rect 298112 459406 298140 480023
rect 298480 475402 298508 480023
rect 298204 475374 298508 475402
rect 298204 466342 298232 475374
rect 298940 470594 298968 480023
rect 299860 470594 299888 480134
rect 357440 478848 357492 478854
rect 357440 478790 357492 478796
rect 356704 478576 356756 478582
rect 356704 478518 356756 478524
rect 298296 470566 298968 470594
rect 299492 470566 299888 470594
rect 298192 466336 298244 466342
rect 298192 466278 298244 466284
rect 298296 466274 298324 470566
rect 298284 466268 298336 466274
rect 298284 466210 298336 466216
rect 299492 466206 299520 470566
rect 299480 466200 299532 466206
rect 299480 466142 299532 466148
rect 339776 461100 339828 461106
rect 339776 461042 339828 461048
rect 338304 461032 338356 461038
rect 338302 461000 338304 461009
rect 339788 461009 339816 461042
rect 338356 461000 338358 461009
rect 338302 460935 338358 460944
rect 339774 461000 339830 461009
rect 339774 460935 339776 460944
rect 339828 460935 339830 460944
rect 350998 461000 351054 461009
rect 350998 460935 351000 460944
rect 339776 460906 339828 460912
rect 351052 460935 351054 460944
rect 351000 460906 351052 460912
rect 298100 459400 298152 459406
rect 298100 459342 298152 459348
rect 281540 459332 281592 459338
rect 281540 459274 281592 459280
rect 280160 459264 280212 459270
rect 280160 459206 280212 459212
rect 276020 459196 276072 459202
rect 276020 459138 276072 459144
rect 271880 459128 271932 459134
rect 271880 459070 271932 459076
rect 263600 459060 263652 459066
rect 263600 459002 263652 459008
rect 258080 458992 258132 458998
rect 258080 458934 258132 458940
rect 247040 458856 247092 458862
rect 223578 458824 223634 458833
rect 247040 458798 247092 458804
rect 223578 458759 223634 458768
rect 356612 456136 356664 456142
rect 356612 456078 356664 456084
rect 244738 375048 244794 375057
rect 244738 374983 244794 374992
rect 270498 375048 270554 375057
rect 270498 374983 270554 374992
rect 283010 375048 283066 375057
rect 283010 374983 283066 374992
rect 311806 375048 311862 375057
rect 311806 374983 311862 374992
rect 220912 374536 220964 374542
rect 220912 374478 220964 374484
rect 244278 374504 244334 374513
rect 220728 373312 220780 373318
rect 220728 373254 220780 373260
rect 220740 373114 220768 373254
rect 220728 373108 220780 373114
rect 220728 373050 220780 373056
rect 220728 372428 220780 372434
rect 220728 372370 220780 372376
rect 220084 372292 220136 372298
rect 220084 372234 220136 372240
rect 220096 371346 220124 372234
rect 220740 372094 220768 372370
rect 220728 372088 220780 372094
rect 220728 372030 220780 372036
rect 220924 371890 220952 374478
rect 221556 374468 221608 374474
rect 244278 374439 244334 374448
rect 221556 374410 221608 374416
rect 221004 372360 221056 372366
rect 221004 372302 221056 372308
rect 220912 371884 220964 371890
rect 220912 371826 220964 371832
rect 220726 371784 220782 371793
rect 220726 371719 220782 371728
rect 220740 371385 220768 371719
rect 220726 371376 220782 371385
rect 220084 371340 220136 371346
rect 220726 371311 220782 371320
rect 220084 371282 220136 371288
rect 220820 371272 220872 371278
rect 220820 371214 220872 371220
rect 220832 353462 220860 371214
rect 220820 353456 220872 353462
rect 220820 353398 220872 353404
rect 220924 353394 220952 371826
rect 220912 353388 220964 353394
rect 220912 353330 220964 353336
rect 221016 353326 221044 372302
rect 221568 372230 221596 374410
rect 244292 374406 244320 374439
rect 240692 374400 240744 374406
rect 240692 374342 240744 374348
rect 244280 374400 244332 374406
rect 244280 374342 244332 374348
rect 221648 374332 221700 374338
rect 221648 374274 221700 374280
rect 221556 372224 221608 372230
rect 221556 372166 221608 372172
rect 221660 372026 221688 374274
rect 222106 374232 222162 374241
rect 222106 374167 222162 374176
rect 222014 374096 222070 374105
rect 222014 374031 222070 374040
rect 221924 372360 221976 372366
rect 221924 372302 221976 372308
rect 221648 372020 221700 372026
rect 221648 371962 221700 371968
rect 221936 371550 221964 372302
rect 222028 372065 222056 374031
rect 222120 372201 222148 374167
rect 240704 374066 240732 374342
rect 240784 374332 240836 374338
rect 240784 374274 240836 374280
rect 240692 374060 240744 374066
rect 240692 374002 240744 374008
rect 235998 373144 236054 373153
rect 235998 373079 236054 373088
rect 224316 372904 224368 372910
rect 224144 372852 224316 372858
rect 224144 372846 224368 372852
rect 224144 372842 224356 372846
rect 224132 372836 224356 372842
rect 224184 372830 224356 372836
rect 224132 372778 224184 372784
rect 236012 372638 236040 373079
rect 236092 372700 236144 372706
rect 236092 372642 236144 372648
rect 236000 372632 236052 372638
rect 236104 372609 236132 372642
rect 236000 372574 236052 372580
rect 236090 372600 236146 372609
rect 236090 372535 236146 372544
rect 238114 372600 238170 372609
rect 238114 372535 238170 372544
rect 239310 372600 239366 372609
rect 239310 372535 239366 372544
rect 240414 372600 240470 372609
rect 240414 372535 240470 372544
rect 222106 372192 222162 372201
rect 222106 372127 222162 372136
rect 222014 372056 222070 372065
rect 222014 371991 222070 372000
rect 222108 371816 222160 371822
rect 222108 371758 222160 371764
rect 221924 371544 221976 371550
rect 221924 371486 221976 371492
rect 222120 371278 222148 371758
rect 238128 371550 238156 372535
rect 223120 371544 223172 371550
rect 223120 371486 223172 371492
rect 237380 371544 237432 371550
rect 237380 371486 237432 371492
rect 238116 371544 238168 371550
rect 238116 371486 238168 371492
rect 223132 371278 223160 371486
rect 237392 371414 237420 371486
rect 239324 371482 239352 372535
rect 240428 371618 240456 372535
rect 240796 372026 240824 374274
rect 244752 374066 244780 374983
rect 247590 374504 247646 374513
rect 247590 374439 247646 374448
rect 253478 374504 253534 374513
rect 253478 374439 253534 374448
rect 265254 374504 265310 374513
rect 265254 374439 265310 374448
rect 247604 374338 247632 374439
rect 247592 374332 247644 374338
rect 247592 374274 247644 374280
rect 253492 374066 253520 374439
rect 265268 374270 265296 374439
rect 265256 374264 265308 374270
rect 265256 374206 265308 374212
rect 270314 374232 270370 374241
rect 270512 374202 270540 374983
rect 270314 374167 270370 374176
rect 270500 374196 270552 374202
rect 270222 374096 270278 374105
rect 240876 374060 240928 374066
rect 240876 374002 240928 374008
rect 244740 374060 244792 374066
rect 244740 374002 244792 374008
rect 250628 374060 250680 374066
rect 250628 374002 250680 374008
rect 253480 374060 253532 374066
rect 270222 374031 270278 374040
rect 253480 374002 253532 374008
rect 240888 372230 240916 374002
rect 242898 373280 242954 373289
rect 242898 373215 242954 373224
rect 242912 373182 242940 373215
rect 242900 373176 242952 373182
rect 242900 373118 242952 373124
rect 241518 372600 241574 372609
rect 241518 372535 241574 372544
rect 245658 372600 245714 372609
rect 245658 372535 245714 372544
rect 248418 372600 248474 372609
rect 248418 372535 248474 372544
rect 240876 372224 240928 372230
rect 240876 372166 240928 372172
rect 240784 372020 240836 372026
rect 240784 371962 240836 371968
rect 241532 371822 241560 372535
rect 245672 372162 245700 372535
rect 248432 372434 248460 372535
rect 248420 372428 248472 372434
rect 248420 372370 248472 372376
rect 245660 372156 245712 372162
rect 245660 372098 245712 372104
rect 250640 371890 250668 374002
rect 258078 373824 258134 373833
rect 258078 373759 258134 373768
rect 262862 373824 262918 373833
rect 262862 373759 262918 373768
rect 253938 373144 253994 373153
rect 253938 373079 253940 373088
rect 253992 373079 253994 373088
rect 255410 373144 255466 373153
rect 255410 373079 255466 373088
rect 253940 373050 253992 373056
rect 255424 373046 255452 373079
rect 255412 373040 255464 373046
rect 255412 372982 255464 372988
rect 256700 372972 256752 372978
rect 256700 372914 256752 372920
rect 256712 372609 256740 372914
rect 258092 372774 258120 373759
rect 262772 373380 262824 373386
rect 262772 373322 262824 373328
rect 261298 373280 261354 373289
rect 261298 373215 261300 373224
rect 261352 373215 261354 373224
rect 261300 373186 261352 373192
rect 259644 372904 259696 372910
rect 259644 372846 259696 372852
rect 259460 372836 259512 372842
rect 259460 372778 259512 372784
rect 258080 372768 258132 372774
rect 258080 372710 258132 372716
rect 259472 372609 259500 372778
rect 259656 372609 259684 372846
rect 251178 372600 251234 372609
rect 251178 372535 251234 372544
rect 256698 372600 256754 372609
rect 256698 372535 256754 372544
rect 259458 372600 259514 372609
rect 259458 372535 259514 372544
rect 259642 372600 259698 372609
rect 259642 372535 259698 372544
rect 251192 372094 251220 372535
rect 251180 372088 251232 372094
rect 251180 372030 251232 372036
rect 250628 371884 250680 371890
rect 250628 371826 250680 371832
rect 241520 371816 241572 371822
rect 241520 371758 241572 371764
rect 247038 371648 247094 371657
rect 240416 371612 240468 371618
rect 240416 371554 240468 371560
rect 241428 371612 241480 371618
rect 247038 371583 247094 371592
rect 249890 371648 249946 371657
rect 249890 371583 249946 371592
rect 251178 371648 251234 371657
rect 251178 371583 251234 371592
rect 241428 371554 241480 371560
rect 239312 371476 239364 371482
rect 239312 371418 239364 371424
rect 241440 371414 241468 371554
rect 237380 371408 237432 371414
rect 237380 371350 237432 371356
rect 241428 371408 241480 371414
rect 241428 371350 241480 371356
rect 222108 371272 222160 371278
rect 222108 371214 222160 371220
rect 223120 371272 223172 371278
rect 223120 371214 223172 371220
rect 247052 369850 247080 371583
rect 249798 371376 249854 371385
rect 249798 371311 249800 371320
rect 249852 371311 249854 371320
rect 249800 371282 249852 371288
rect 247040 369844 247092 369850
rect 247040 369786 247092 369792
rect 249904 369102 249932 371583
rect 251192 371278 251220 371583
rect 262784 371521 262812 373322
rect 262876 371958 262904 373759
rect 263690 373552 263746 373561
rect 263690 373487 263692 373496
rect 263744 373487 263746 373496
rect 263692 373458 263744 373464
rect 269210 373416 269266 373425
rect 269210 373351 269212 373360
rect 269264 373351 269266 373360
rect 269212 373322 269264 373328
rect 270236 372201 270264 374031
rect 270222 372192 270278 372201
rect 270222 372127 270278 372136
rect 270328 372065 270356 374167
rect 270500 374138 270552 374144
rect 283024 374134 283052 374983
rect 304264 374808 304316 374814
rect 304264 374750 304316 374756
rect 283012 374128 283064 374134
rect 283012 374070 283064 374076
rect 271970 373144 272026 373153
rect 271970 373079 272026 373088
rect 300858 373144 300914 373153
rect 300858 373079 300914 373088
rect 270314 372056 270370 372065
rect 270314 371991 270370 372000
rect 262864 371952 262916 371958
rect 271984 371929 272012 373079
rect 273258 372600 273314 372609
rect 273258 372535 273260 372544
rect 273312 372535 273314 372544
rect 273260 372506 273312 372512
rect 276294 372464 276350 372473
rect 276294 372399 276350 372408
rect 262864 371894 262916 371900
rect 271970 371920 272026 371929
rect 271970 371855 272026 371864
rect 275376 371884 275428 371890
rect 275376 371826 275428 371832
rect 275388 371793 275416 371826
rect 276308 371822 276336 372399
rect 278686 372328 278742 372337
rect 278686 372263 278742 372272
rect 276296 371816 276348 371822
rect 275374 371784 275430 371793
rect 273260 371748 273312 371754
rect 276296 371758 276348 371764
rect 275374 371719 275430 371728
rect 273260 371690 273312 371696
rect 262770 371512 262826 371521
rect 262770 371447 262826 371456
rect 264978 371512 265034 371521
rect 264978 371447 265034 371456
rect 252558 371376 252614 371385
rect 252558 371311 252614 371320
rect 255318 371376 255374 371385
rect 255318 371311 255374 371320
rect 258170 371376 258226 371385
rect 258170 371311 258226 371320
rect 260838 371376 260894 371385
rect 260838 371311 260894 371320
rect 263598 371376 263654 371385
rect 263598 371311 263654 371320
rect 251180 371272 251232 371278
rect 251180 371214 251232 371220
rect 249892 369096 249944 369102
rect 249892 369038 249944 369044
rect 252572 368966 252600 371311
rect 252560 368960 252612 368966
rect 252560 368902 252612 368908
rect 255332 368898 255360 371311
rect 258184 369374 258212 371311
rect 260852 369442 260880 371311
rect 263612 369510 263640 371311
rect 264992 369646 265020 371447
rect 266358 371376 266414 371385
rect 266358 371311 266414 371320
rect 267738 371376 267794 371385
rect 267738 371311 267794 371320
rect 264980 369640 265032 369646
rect 264980 369582 265032 369588
rect 263600 369504 263652 369510
rect 263600 369446 263652 369452
rect 260840 369436 260892 369442
rect 260840 369378 260892 369384
rect 258172 369368 258224 369374
rect 258172 369310 258224 369316
rect 255320 368892 255372 368898
rect 255320 368834 255372 368840
rect 266372 368490 266400 371311
rect 267752 369578 267780 371311
rect 273272 370394 273300 371690
rect 278700 371686 278728 372263
rect 278688 371680 278740 371686
rect 278688 371622 278740 371628
rect 273350 371512 273406 371521
rect 273350 371447 273406 371456
rect 273260 370388 273312 370394
rect 273260 370330 273312 370336
rect 267740 369572 267792 369578
rect 267740 369514 267792 369520
rect 273364 369306 273392 371447
rect 276018 371376 276074 371385
rect 276018 371311 276074 371320
rect 277766 371376 277822 371385
rect 277766 371311 277822 371320
rect 280158 371376 280214 371385
rect 280158 371311 280214 371320
rect 285678 371376 285734 371385
rect 285678 371311 285734 371320
rect 287242 371376 287298 371385
rect 287242 371311 287298 371320
rect 289818 371376 289874 371385
rect 289818 371311 289874 371320
rect 292578 371376 292634 371385
rect 292578 371311 292634 371320
rect 295338 371376 295394 371385
rect 295338 371311 295394 371320
rect 298098 371376 298154 371385
rect 298098 371311 298154 371320
rect 273352 369300 273404 369306
rect 273352 369242 273404 369248
rect 276032 369034 276060 371311
rect 277780 370462 277808 371311
rect 280172 370598 280200 371311
rect 285692 370666 285720 371311
rect 287256 370734 287284 371311
rect 289832 370802 289860 371311
rect 292592 370870 292620 371311
rect 295352 371074 295380 371311
rect 295340 371068 295392 371074
rect 295340 371010 295392 371016
rect 292580 370864 292632 370870
rect 292580 370806 292632 370812
rect 289820 370796 289872 370802
rect 289820 370738 289872 370744
rect 287244 370728 287296 370734
rect 287244 370670 287296 370676
rect 285680 370660 285732 370666
rect 285680 370602 285732 370608
rect 280160 370592 280212 370598
rect 280160 370534 280212 370540
rect 298112 370530 298140 371311
rect 300872 370938 300900 373079
rect 304276 372502 304304 374750
rect 305000 374740 305052 374746
rect 305000 374682 305052 374688
rect 305012 372570 305040 374682
rect 311820 374678 311848 374983
rect 311808 374672 311860 374678
rect 311808 374614 311860 374620
rect 320914 374640 320970 374649
rect 320914 374575 320916 374584
rect 320968 374575 320970 374584
rect 320916 374546 320968 374552
rect 310518 372600 310574 372609
rect 305000 372564 305052 372570
rect 310518 372535 310574 372544
rect 313278 372600 313334 372609
rect 313278 372535 313280 372544
rect 305000 372506 305052 372512
rect 310532 372502 310560 372535
rect 313332 372535 313334 372544
rect 313280 372506 313332 372512
rect 304264 372496 304316 372502
rect 310520 372496 310572 372502
rect 304264 372438 304316 372444
rect 304998 372464 305054 372473
rect 310520 372438 310572 372444
rect 304998 372399 305054 372408
rect 305012 371754 305040 372399
rect 317418 371784 317474 371793
rect 305000 371748 305052 371754
rect 317418 371719 317474 371728
rect 305000 371690 305052 371696
rect 302238 371376 302294 371385
rect 302238 371311 302294 371320
rect 307758 371376 307814 371385
rect 307758 371311 307814 371320
rect 302252 371142 302280 371311
rect 302240 371136 302292 371142
rect 302240 371078 302292 371084
rect 307772 371006 307800 371311
rect 317432 371210 317460 371719
rect 325882 371648 325938 371657
rect 325882 371583 325938 371592
rect 322938 371376 322994 371385
rect 322938 371311 322994 371320
rect 317420 371204 317472 371210
rect 317420 371146 317472 371152
rect 307760 371000 307812 371006
rect 307760 370942 307812 370948
rect 300860 370932 300912 370938
rect 300860 370874 300912 370880
rect 298100 370524 298152 370530
rect 298100 370466 298152 370472
rect 277768 370456 277820 370462
rect 277768 370398 277820 370404
rect 322952 369714 322980 371311
rect 325896 369782 325924 371583
rect 343086 371376 343142 371385
rect 342904 371340 342956 371346
rect 343086 371311 343142 371320
rect 343454 371376 343510 371385
rect 343454 371311 343456 371320
rect 342904 371282 342956 371288
rect 325884 369776 325936 369782
rect 325884 369718 325936 369724
rect 322940 369708 322992 369714
rect 322940 369650 322992 369656
rect 276020 369028 276072 369034
rect 276020 368970 276072 368976
rect 266360 368484 266412 368490
rect 266360 368426 266412 368432
rect 342916 356726 342944 371282
rect 343100 371278 343128 371311
rect 343508 371311 343510 371320
rect 343456 371282 343508 371288
rect 343088 371272 343140 371278
rect 343088 371214 343140 371220
rect 343100 364342 343128 371214
rect 343088 364336 343140 364342
rect 343088 364278 343140 364284
rect 342904 356720 342956 356726
rect 342904 356662 342956 356668
rect 356624 355434 356652 456078
rect 340052 355428 340104 355434
rect 340052 355370 340104 355376
rect 356612 355428 356664 355434
rect 356612 355370 356664 355376
rect 340064 355065 340092 355370
rect 351736 355360 351788 355366
rect 351736 355302 351788 355308
rect 351748 355065 351776 355302
rect 340050 355056 340106 355065
rect 340050 354991 340106 355000
rect 351734 355056 351790 355065
rect 356624 355026 356652 355370
rect 351734 354991 351790 355000
rect 356612 355020 356664 355026
rect 356612 354962 356664 354968
rect 338120 354816 338172 354822
rect 338118 354784 338120 354793
rect 338172 354784 338174 354793
rect 338118 354719 338174 354728
rect 221004 353320 221056 353326
rect 221004 353262 221056 353268
rect 250718 269784 250774 269793
rect 250718 269719 250774 269728
rect 250732 269346 250760 269719
rect 283470 269648 283526 269657
rect 283470 269583 283526 269592
rect 288254 269648 288310 269657
rect 288254 269583 288310 269592
rect 291014 269648 291070 269657
rect 291014 269583 291070 269592
rect 293406 269648 293462 269657
rect 293406 269583 293462 269592
rect 305918 269648 305974 269657
rect 305918 269583 305974 269592
rect 318430 269648 318486 269657
rect 318430 269583 318486 269592
rect 250720 269340 250772 269346
rect 250720 269282 250772 269288
rect 283484 269278 283512 269583
rect 283472 269272 283524 269278
rect 283472 269214 283524 269220
rect 288268 269210 288296 269583
rect 288256 269204 288308 269210
rect 288256 269146 288308 269152
rect 291028 269142 291056 269583
rect 291016 269136 291068 269142
rect 291016 269078 291068 269084
rect 236000 268932 236052 268938
rect 236000 268874 236052 268880
rect 236012 267986 236040 268874
rect 243082 268832 243138 268841
rect 243082 268767 243138 268776
rect 258078 268832 258134 268841
rect 258078 268767 258134 268776
rect 261666 268832 261722 268841
rect 261666 268767 261722 268776
rect 236000 267980 236052 267986
rect 236000 267922 236052 267928
rect 220818 267880 220874 267889
rect 220818 267815 220874 267824
rect 220832 251190 220860 267815
rect 230388 265056 230440 265062
rect 230388 264998 230440 265004
rect 230400 264722 230428 264998
rect 233148 264988 233200 264994
rect 233148 264930 233200 264936
rect 230388 264716 230440 264722
rect 230388 264658 230440 264664
rect 233160 264654 233188 264930
rect 233148 264648 233200 264654
rect 233148 264590 233200 264596
rect 220820 251184 220872 251190
rect 220820 251126 220872 251132
rect 221372 251184 221424 251190
rect 221372 251126 221424 251132
rect 221384 249830 221412 251126
rect 236012 250578 236040 267922
rect 243096 267918 243124 268767
rect 247040 267980 247092 267986
rect 247040 267922 247092 267928
rect 243084 267912 243136 267918
rect 243084 267854 243136 267860
rect 247052 267714 247080 267922
rect 258092 267850 258120 268767
rect 258080 267844 258132 267850
rect 258080 267786 258132 267792
rect 261680 267782 261708 268767
rect 293420 268734 293448 269583
rect 298468 268864 298520 268870
rect 295890 268832 295946 268841
rect 295890 268767 295892 268776
rect 295944 268767 295946 268776
rect 298466 268832 298468 268841
rect 298520 268832 298522 268841
rect 298466 268767 298522 268776
rect 300858 268832 300914 268841
rect 300858 268767 300914 268776
rect 303434 268832 303490 268841
rect 303434 268767 303490 268776
rect 295892 268738 295944 268744
rect 293408 268728 293460 268734
rect 293408 268670 293460 268676
rect 300872 268666 300900 268767
rect 300860 268660 300912 268666
rect 300860 268602 300912 268608
rect 303448 268530 303476 268767
rect 305932 268598 305960 269583
rect 305920 268592 305972 268598
rect 305920 268534 305972 268540
rect 303436 268524 303488 268530
rect 303436 268466 303488 268472
rect 318444 268394 318472 269583
rect 323306 269104 323362 269113
rect 323306 269039 323362 269048
rect 323320 268462 323348 269039
rect 323308 268456 323360 268462
rect 323308 268398 323360 268404
rect 318432 268388 318484 268394
rect 318432 268330 318484 268336
rect 265162 268152 265218 268161
rect 265162 268087 265218 268096
rect 275926 268152 275982 268161
rect 275926 268087 275982 268096
rect 261668 267776 261720 267782
rect 255318 267744 255374 267753
rect 247040 267708 247092 267714
rect 255318 267679 255320 267688
rect 247040 267650 247092 267656
rect 255372 267679 255374 267688
rect 258262 267744 258318 267753
rect 258262 267679 258318 267688
rect 260838 267744 260894 267753
rect 261668 267718 261720 267724
rect 263598 267744 263654 267753
rect 260838 267679 260894 267688
rect 263598 267679 263654 267688
rect 264978 267744 265034 267753
rect 264978 267679 265034 267688
rect 255320 267650 255372 267656
rect 258276 267170 258304 267679
rect 258264 267164 258316 267170
rect 258264 267106 258316 267112
rect 260852 267102 260880 267679
rect 263612 267442 263640 267679
rect 264992 267510 265020 267679
rect 264980 267504 265032 267510
rect 264980 267446 265032 267452
rect 263600 267436 263652 267442
rect 263600 267378 263652 267384
rect 260840 267096 260892 267102
rect 255318 267064 255374 267073
rect 260840 267038 260892 267044
rect 255318 266999 255374 267008
rect 255332 266966 255360 266999
rect 255320 266960 255372 266966
rect 247038 266928 247094 266937
rect 247038 266863 247094 266872
rect 252558 266928 252614 266937
rect 255320 266902 255372 266908
rect 252558 266863 252560 266872
rect 247052 266830 247080 266863
rect 252612 266863 252614 266872
rect 252560 266834 252612 266840
rect 247040 266824 247092 266830
rect 247040 266766 247092 266772
rect 249798 266656 249854 266665
rect 249798 266591 249854 266600
rect 244370 266520 244426 266529
rect 244370 266455 244426 266464
rect 244278 266384 244334 266393
rect 244278 266319 244334 266328
rect 244292 265606 244320 266319
rect 244280 265600 244332 265606
rect 244280 265542 244332 265548
rect 244384 264586 244412 266455
rect 245658 266384 245714 266393
rect 245658 266319 245714 266328
rect 247038 266384 247094 266393
rect 247038 266319 247094 266328
rect 248510 266384 248566 266393
rect 248510 266319 248566 266328
rect 245672 266082 245700 266319
rect 247052 266286 247080 266319
rect 247040 266280 247092 266286
rect 247040 266222 247092 266228
rect 245660 266076 245712 266082
rect 245660 266018 245712 266024
rect 248524 265946 248552 266319
rect 249812 266014 249840 266591
rect 251270 266520 251326 266529
rect 251270 266455 251326 266464
rect 259550 266520 259606 266529
rect 259550 266455 259606 266464
rect 251178 266384 251234 266393
rect 251178 266319 251234 266328
rect 251192 266150 251220 266319
rect 251284 266218 251312 266455
rect 252558 266384 252614 266393
rect 252558 266319 252614 266328
rect 253938 266384 253994 266393
rect 253938 266319 253994 266328
rect 256698 266384 256754 266393
rect 256698 266319 256754 266328
rect 259458 266384 259514 266393
rect 259458 266319 259514 266328
rect 251272 266212 251324 266218
rect 251272 266154 251324 266160
rect 251180 266144 251232 266150
rect 251180 266086 251232 266092
rect 249800 266008 249852 266014
rect 249800 265950 249852 265956
rect 248512 265940 248564 265946
rect 248512 265882 248564 265888
rect 252572 265878 252600 266319
rect 252560 265872 252612 265878
rect 252560 265814 252612 265820
rect 253952 264790 253980 266319
rect 253940 264784 253992 264790
rect 253940 264726 253992 264732
rect 244372 264580 244424 264586
rect 244372 264522 244424 264528
rect 256712 264314 256740 266319
rect 259472 264654 259500 266319
rect 259564 264722 259592 266455
rect 262218 266384 262274 266393
rect 262218 266319 262220 266328
rect 262272 266319 262274 266328
rect 263598 266384 263654 266393
rect 263598 266319 263654 266328
rect 262220 266290 262272 266296
rect 263612 265810 263640 266319
rect 263600 265804 263652 265810
rect 263600 265746 263652 265752
rect 265176 265742 265204 268087
rect 267830 267744 267886 267753
rect 267830 267679 267886 267688
rect 270498 267744 270554 267753
rect 270498 267679 270554 267688
rect 273258 267744 273314 267753
rect 273258 267679 273314 267688
rect 267844 267578 267872 267679
rect 267832 267572 267884 267578
rect 267832 267514 267884 267520
rect 270512 267238 270540 267679
rect 273272 267374 273300 267679
rect 273260 267368 273312 267374
rect 273260 267310 273312 267316
rect 270500 267232 270552 267238
rect 270500 267174 270552 267180
rect 273258 267064 273314 267073
rect 275940 267034 275968 268087
rect 276018 267744 276074 267753
rect 276018 267679 276074 267688
rect 277030 267744 277086 267753
rect 277030 267679 277086 267688
rect 278134 267744 278190 267753
rect 278134 267679 278190 267688
rect 280158 267744 280214 267753
rect 280158 267679 280214 267688
rect 276032 267306 276060 267679
rect 276020 267300 276072 267306
rect 276020 267242 276072 267248
rect 277044 267102 277072 267679
rect 278148 267238 278176 267679
rect 280172 267646 280200 267679
rect 280160 267640 280212 267646
rect 280160 267582 280212 267588
rect 343454 267472 343510 267481
rect 343454 267407 343510 267416
rect 343468 267306 343496 267407
rect 343456 267300 343508 267306
rect 343456 267242 343508 267248
rect 278136 267232 278188 267238
rect 356612 267232 356664 267238
rect 278136 267174 278188 267180
rect 279146 267200 279202 267209
rect 356612 267174 356664 267180
rect 279146 267135 279148 267144
rect 279200 267135 279202 267144
rect 279148 267106 279200 267112
rect 356624 267102 356652 267174
rect 277032 267096 277084 267102
rect 356612 267096 356664 267102
rect 277032 267038 277084 267044
rect 343454 267064 343510 267073
rect 273258 266999 273260 267008
rect 273312 266999 273314 267008
rect 275928 267028 275980 267034
rect 273260 266970 273312 266976
rect 356612 267038 356664 267044
rect 343454 266999 343510 267008
rect 275928 266970 275980 266976
rect 285678 266928 285734 266937
rect 285678 266863 285734 266872
rect 285692 266762 285720 266863
rect 285680 266756 285732 266762
rect 285680 266698 285732 266704
rect 266358 266520 266414 266529
rect 266358 266455 266414 266464
rect 265164 265736 265216 265742
rect 265164 265678 265216 265684
rect 266372 265674 266400 266455
rect 343468 266422 343496 266999
rect 343456 266416 343508 266422
rect 266450 266384 266506 266393
rect 266450 266319 266506 266328
rect 267738 266384 267794 266393
rect 267738 266319 267794 266328
rect 269118 266384 269174 266393
rect 269118 266319 269174 266328
rect 270498 266384 270554 266393
rect 270498 266319 270554 266328
rect 273166 266384 273222 266393
rect 343456 266358 343508 266364
rect 273166 266319 273222 266328
rect 266360 265668 266412 265674
rect 266360 265610 266412 265616
rect 259552 264716 259604 264722
rect 259552 264658 259604 264664
rect 259460 264648 259512 264654
rect 259460 264590 259512 264596
rect 256700 264308 256752 264314
rect 256700 264250 256752 264256
rect 266464 251190 266492 266319
rect 266452 251184 266504 251190
rect 266452 251126 266504 251132
rect 236000 250572 236052 250578
rect 236000 250514 236052 250520
rect 267752 250510 267780 266319
rect 269132 264246 269160 266319
rect 270512 264858 270540 266319
rect 273180 264926 273208 266319
rect 273168 264920 273220 264926
rect 273168 264862 273220 264868
rect 270500 264852 270552 264858
rect 270500 264794 270552 264800
rect 269120 264240 269172 264246
rect 269120 264182 269172 264188
rect 340052 250640 340104 250646
rect 340052 250582 340104 250588
rect 338488 250572 338540 250578
rect 338488 250514 338540 250520
rect 267740 250504 267792 250510
rect 267740 250446 267792 250452
rect 338500 249937 338528 250514
rect 340064 249937 340092 250582
rect 351736 250504 351788 250510
rect 351736 250446 351788 250452
rect 351748 249937 351776 250446
rect 338486 249928 338542 249937
rect 338486 249863 338542 249872
rect 340050 249928 340106 249937
rect 340050 249863 340106 249872
rect 351734 249928 351790 249937
rect 351734 249863 351790 249872
rect 221372 249824 221424 249830
rect 221372 249766 221424 249772
rect 261022 164792 261078 164801
rect 261022 164727 261078 164736
rect 261036 164354 261064 164727
rect 288254 164656 288310 164665
rect 288254 164591 288310 164600
rect 305918 164656 305974 164665
rect 305918 164591 305974 164600
rect 265898 164520 265954 164529
rect 265898 164455 265954 164464
rect 261024 164348 261076 164354
rect 261024 164290 261076 164296
rect 265912 163946 265940 164455
rect 288268 164286 288296 164591
rect 288256 164280 288308 164286
rect 288256 164222 288308 164228
rect 298466 164248 298522 164257
rect 298466 164183 298522 164192
rect 300858 164248 300914 164257
rect 300858 164183 300914 164192
rect 303434 164248 303490 164257
rect 303434 164183 303490 164192
rect 265900 163940 265952 163946
rect 265900 163882 265952 163888
rect 285956 163872 286008 163878
rect 285954 163840 285956 163849
rect 286008 163840 286010 163849
rect 285954 163775 286010 163784
rect 298480 163742 298508 164183
rect 298468 163736 298520 163742
rect 298468 163678 298520 163684
rect 300872 163674 300900 164183
rect 303448 163810 303476 164183
rect 303436 163804 303488 163810
rect 303436 163746 303488 163752
rect 300860 163668 300912 163674
rect 300860 163610 300912 163616
rect 305932 163606 305960 164591
rect 313370 164248 313426 164257
rect 313370 164183 313426 164192
rect 305920 163600 305972 163606
rect 305920 163542 305972 163548
rect 313384 163538 313412 164183
rect 313372 163532 313424 163538
rect 313372 163474 313424 163480
rect 220452 163464 220504 163470
rect 220452 163406 220504 163412
rect 220464 162926 220492 163406
rect 235998 163160 236054 163169
rect 235998 163095 236054 163104
rect 264978 163160 265034 163169
rect 264978 163095 265034 163104
rect 276110 163160 276166 163169
rect 276110 163095 276166 163104
rect 220452 162920 220504 162926
rect 220452 162862 220504 162868
rect 236012 145382 236040 163095
rect 236644 162988 236696 162994
rect 236644 162930 236696 162936
rect 236090 162752 236146 162761
rect 236090 162687 236146 162696
rect 236104 145450 236132 162687
rect 236656 146198 236684 162930
rect 263690 162888 263746 162897
rect 263690 162823 263746 162832
rect 237378 162752 237434 162761
rect 237378 162687 237434 162696
rect 240138 162752 240194 162761
rect 240138 162687 240194 162696
rect 241518 162752 241574 162761
rect 241518 162687 241574 162696
rect 242898 162752 242954 162761
rect 242898 162687 242954 162696
rect 244370 162752 244426 162761
rect 244370 162687 244426 162696
rect 245658 162752 245714 162761
rect 245658 162687 245714 162696
rect 247038 162752 247094 162761
rect 247038 162687 247094 162696
rect 248234 162752 248290 162761
rect 248234 162687 248290 162696
rect 248418 162752 248474 162761
rect 248418 162687 248474 162696
rect 249798 162752 249854 162761
rect 249798 162687 249854 162696
rect 250626 162752 250682 162761
rect 250626 162687 250682 162696
rect 251178 162752 251234 162761
rect 251178 162687 251234 162696
rect 252558 162752 252614 162761
rect 252558 162687 252614 162696
rect 253570 162752 253626 162761
rect 253570 162687 253626 162696
rect 253938 162752 253994 162761
rect 253938 162687 253994 162696
rect 255318 162752 255374 162761
rect 255318 162687 255374 162696
rect 256146 162752 256202 162761
rect 256146 162687 256202 162696
rect 256698 162752 256754 162761
rect 256698 162687 256754 162696
rect 258354 162752 258410 162761
rect 258354 162687 258410 162696
rect 259458 162752 259514 162761
rect 259458 162687 259514 162696
rect 260838 162752 260894 162761
rect 260838 162687 260894 162696
rect 262218 162752 262274 162761
rect 262218 162687 262274 162696
rect 263598 162752 263654 162761
rect 263598 162687 263654 162696
rect 236644 146192 236696 146198
rect 236644 146134 236696 146140
rect 237392 145897 237420 162687
rect 238758 161528 238814 161537
rect 238758 161463 238814 161472
rect 238772 148850 238800 161463
rect 240152 148986 240180 162687
rect 240140 148980 240192 148986
rect 240140 148922 240192 148928
rect 241532 148918 241560 162687
rect 241520 148912 241572 148918
rect 241520 148854 241572 148860
rect 238760 148844 238812 148850
rect 238760 148786 238812 148792
rect 237378 145888 237434 145897
rect 237378 145823 237434 145832
rect 242912 145518 242940 162687
rect 244278 162072 244334 162081
rect 244278 162007 244334 162016
rect 244292 145722 244320 162007
rect 244384 145790 244412 162687
rect 244372 145784 244424 145790
rect 244372 145726 244424 145732
rect 244280 145716 244332 145722
rect 244280 145658 244332 145664
rect 245672 145586 245700 162687
rect 247052 145654 247080 162687
rect 248248 162042 248276 162687
rect 248236 162036 248288 162042
rect 248236 161978 248288 161984
rect 248432 145858 248460 162687
rect 249812 145926 249840 162687
rect 250640 162110 250668 162687
rect 250628 162104 250680 162110
rect 250628 162046 250680 162052
rect 251192 145994 251220 162687
rect 251270 162072 251326 162081
rect 251270 162007 251326 162016
rect 251180 145988 251232 145994
rect 251180 145930 251232 145936
rect 249800 145920 249852 145926
rect 249800 145862 249852 145868
rect 248420 145852 248472 145858
rect 248420 145794 248472 145800
rect 247040 145648 247092 145654
rect 247040 145590 247092 145596
rect 245660 145580 245712 145586
rect 245660 145522 245712 145528
rect 242900 145512 242952 145518
rect 242900 145454 242952 145460
rect 236092 145444 236144 145450
rect 236092 145386 236144 145392
rect 236000 145376 236052 145382
rect 236000 145318 236052 145324
rect 251284 145314 251312 162007
rect 252572 146062 252600 162687
rect 253584 162178 253612 162687
rect 253572 162172 253624 162178
rect 253572 162114 253624 162120
rect 253952 146130 253980 162687
rect 255332 146266 255360 162687
rect 256160 162314 256188 162687
rect 256148 162308 256200 162314
rect 256148 162250 256200 162256
rect 255320 146260 255372 146266
rect 255320 146202 255372 146208
rect 256712 146198 256740 162687
rect 258368 162246 258396 162687
rect 258356 162240 258408 162246
rect 258356 162182 258408 162188
rect 258078 161528 258134 161537
rect 258078 161463 258134 161472
rect 258092 161090 258120 161463
rect 258080 161084 258132 161090
rect 258080 161026 258132 161032
rect 259472 160002 259500 162687
rect 259550 162072 259606 162081
rect 259550 162007 259606 162016
rect 259564 160070 259592 162007
rect 260852 161294 260880 162687
rect 260840 161288 260892 161294
rect 260840 161230 260892 161236
rect 259552 160064 259604 160070
rect 259552 160006 259604 160012
rect 259460 159996 259512 160002
rect 259460 159938 259512 159944
rect 262232 146305 262260 162687
rect 263612 161158 263640 162687
rect 263704 162586 263732 162823
rect 263692 162580 263744 162586
rect 263692 162522 263744 162528
rect 264992 161226 265020 163095
rect 267556 162920 267608 162926
rect 267556 162862 267608 162868
rect 268290 162888 268346 162897
rect 267568 162761 267596 162862
rect 268290 162823 268346 162832
rect 273442 162888 273498 162897
rect 273442 162823 273498 162832
rect 266358 162752 266414 162761
rect 266358 162687 266414 162696
rect 267554 162752 267610 162761
rect 267554 162687 267610 162696
rect 267738 162752 267794 162761
rect 267738 162687 267794 162696
rect 266372 161362 266400 162687
rect 267752 161430 267780 162687
rect 268304 162450 268332 162823
rect 269118 162752 269174 162761
rect 269118 162687 269174 162696
rect 270498 162752 270554 162761
rect 270498 162687 270554 162696
rect 271878 162752 271934 162761
rect 271878 162687 271934 162696
rect 273258 162752 273314 162761
rect 273258 162687 273314 162696
rect 268292 162444 268344 162450
rect 268292 162386 268344 162392
rect 267740 161424 267792 161430
rect 267740 161366 267792 161372
rect 266360 161356 266412 161362
rect 266360 161298 266412 161304
rect 264980 161220 265032 161226
rect 264980 161162 265032 161168
rect 263600 161152 263652 161158
rect 263600 161094 263652 161100
rect 262218 146296 262274 146305
rect 262218 146231 262274 146240
rect 256700 146192 256752 146198
rect 256700 146134 256752 146140
rect 253940 146124 253992 146130
rect 253940 146066 253992 146072
rect 252560 146056 252612 146062
rect 252560 145998 252612 146004
rect 269132 145761 269160 162687
rect 269118 145752 269174 145761
rect 269118 145687 269174 145696
rect 270512 145625 270540 162687
rect 271892 148374 271920 162687
rect 273272 160750 273300 162687
rect 273456 162518 273484 162823
rect 274822 162752 274878 162761
rect 274822 162687 274878 162696
rect 276018 162752 276074 162761
rect 276018 162687 276074 162696
rect 273444 162512 273496 162518
rect 273444 162454 273496 162460
rect 274546 162072 274602 162081
rect 274546 162007 274602 162016
rect 274560 161474 274588 162007
rect 274560 161446 274772 161474
rect 273260 160744 273312 160750
rect 273260 160686 273312 160692
rect 274744 149054 274772 161446
rect 274732 149048 274784 149054
rect 274732 148990 274784 148996
rect 271880 148368 271932 148374
rect 271880 148310 271932 148316
rect 274836 146266 274864 162687
rect 276032 146441 276060 162687
rect 276124 162382 276152 163095
rect 320916 162852 320968 162858
rect 320916 162794 320968 162800
rect 293224 162784 293276 162790
rect 280066 162752 280122 162761
rect 280066 162687 280122 162696
rect 280802 162752 280858 162761
rect 280802 162687 280804 162696
rect 276112 162376 276164 162382
rect 276112 162318 276164 162324
rect 278042 161528 278098 161537
rect 278042 161463 278098 161472
rect 278056 151814 278084 161463
rect 278056 151786 278268 151814
rect 278240 149025 278268 151786
rect 278226 149016 278282 149025
rect 278226 148951 278282 148960
rect 278240 148345 278268 148951
rect 278226 148336 278282 148345
rect 278226 148271 278282 148280
rect 276018 146432 276074 146441
rect 276018 146367 276074 146376
rect 274824 146260 274876 146266
rect 274824 146202 274876 146208
rect 276032 146198 276060 146367
rect 276020 146192 276072 146198
rect 276020 146134 276072 146140
rect 280080 145654 280108 162687
rect 280856 162687 280858 162696
rect 283746 162752 283802 162761
rect 283746 162687 283802 162696
rect 293222 162752 293224 162761
rect 320928 162761 320956 162794
rect 293276 162752 293278 162761
rect 293222 162687 293278 162696
rect 320914 162752 320970 162761
rect 320914 162687 320970 162696
rect 343454 162752 343510 162761
rect 343454 162687 343510 162696
rect 280804 162658 280856 162664
rect 283760 162654 283788 162687
rect 283748 162648 283800 162654
rect 283748 162590 283800 162596
rect 343362 162616 343418 162625
rect 343362 162551 343418 162560
rect 343376 162178 343404 162551
rect 343468 162314 343496 162687
rect 343456 162308 343508 162314
rect 343456 162250 343508 162256
rect 343364 162172 343416 162178
rect 343364 162114 343416 162120
rect 356624 146198 356652 267038
rect 356716 164150 356744 478518
rect 357452 477873 357480 478790
rect 358360 478508 358412 478514
rect 358360 478450 358412 478456
rect 358268 478440 358320 478446
rect 358268 478382 358320 478388
rect 357438 477864 357494 477873
rect 357438 477799 357494 477808
rect 356796 477284 356848 477290
rect 356796 477226 356848 477232
rect 356808 268666 356836 477226
rect 356888 471912 356940 471918
rect 356888 471854 356940 471860
rect 356900 369714 356928 471854
rect 358176 469940 358228 469946
rect 358176 469882 358228 469888
rect 357072 466336 357124 466342
rect 357072 466278 357124 466284
rect 356980 461100 357032 461106
rect 356980 461042 357032 461048
rect 356992 456142 357020 461042
rect 356980 456136 357032 456142
rect 356980 456078 357032 456084
rect 356980 371884 357032 371890
rect 356980 371826 357032 371832
rect 356888 369708 356940 369714
rect 356888 369650 356940 369656
rect 356888 355020 356940 355026
rect 356888 354962 356940 354968
rect 356796 268660 356848 268666
rect 356796 268602 356848 268608
rect 356796 266416 356848 266422
rect 356796 266358 356848 266364
rect 356704 164144 356756 164150
rect 356704 164086 356756 164092
rect 356704 162852 356756 162858
rect 356704 162794 356756 162800
rect 356716 162314 356744 162794
rect 356704 162308 356756 162314
rect 356704 162250 356756 162256
rect 356612 146192 356664 146198
rect 356612 146134 356664 146140
rect 338488 146124 338540 146130
rect 338488 146066 338540 146072
rect 280068 145648 280120 145654
rect 270498 145616 270554 145625
rect 280068 145590 280120 145596
rect 270498 145551 270554 145560
rect 251272 145308 251324 145314
rect 251272 145250 251324 145256
rect 338500 144945 338528 146066
rect 340236 146056 340288 146062
rect 340236 145998 340288 146004
rect 340248 144945 340276 145998
rect 356612 145648 356664 145654
rect 356612 145590 356664 145596
rect 351644 145580 351696 145586
rect 351644 145522 351696 145528
rect 351656 144945 351684 145522
rect 338486 144936 338542 144945
rect 338486 144871 338542 144880
rect 340234 144936 340290 144945
rect 340234 144871 340290 144880
rect 351642 144936 351698 144945
rect 351642 144871 351698 144880
rect 237102 59800 237158 59809
rect 237102 59735 237158 59744
rect 255870 59800 255926 59809
rect 255870 59735 255926 59744
rect 256974 59800 257030 59809
rect 256974 59735 257030 59744
rect 261758 59800 261814 59809
rect 261758 59735 261814 59744
rect 263874 59800 263930 59809
rect 263874 59735 263930 59744
rect 237116 59702 237144 59735
rect 237104 59696 237156 59702
rect 237104 59638 237156 59644
rect 255884 59634 255912 59735
rect 255872 59628 255924 59634
rect 255872 59570 255924 59576
rect 256988 59566 257016 59735
rect 260654 59664 260710 59673
rect 260654 59599 260710 59608
rect 256976 59560 257028 59566
rect 256976 59502 257028 59508
rect 260668 59226 260696 59599
rect 261772 59430 261800 59735
rect 262770 59528 262826 59537
rect 263888 59498 263916 59735
rect 305918 59664 305974 59673
rect 305918 59599 305974 59608
rect 318430 59664 318486 59673
rect 318430 59599 318486 59608
rect 262770 59463 262826 59472
rect 263876 59492 263928 59498
rect 261760 59424 261812 59430
rect 261760 59366 261812 59372
rect 260656 59220 260708 59226
rect 260656 59162 260708 59168
rect 262784 59158 262812 59463
rect 263876 59434 263928 59440
rect 279238 59256 279294 59265
rect 279238 59191 279294 59200
rect 290922 59256 290978 59265
rect 290922 59191 290978 59200
rect 298466 59256 298522 59265
rect 298466 59191 298522 59200
rect 279252 59158 279280 59191
rect 262772 59152 262824 59158
rect 262772 59094 262824 59100
rect 279240 59152 279292 59158
rect 279240 59094 279292 59100
rect 290936 59090 290964 59191
rect 290924 59084 290976 59090
rect 290924 59026 290976 59032
rect 298480 59022 298508 59191
rect 298468 59016 298520 59022
rect 298468 58958 298520 58964
rect 305932 58886 305960 59599
rect 313370 59256 313426 59265
rect 313370 59191 313426 59200
rect 313384 58954 313412 59191
rect 313372 58948 313424 58954
rect 313372 58890 313424 58896
rect 305920 58880 305972 58886
rect 305920 58822 305972 58828
rect 318444 58818 318472 59599
rect 325882 59256 325938 59265
rect 325882 59191 325938 59200
rect 318432 58812 318484 58818
rect 318432 58754 318484 58760
rect 325896 58750 325924 59191
rect 356624 59158 356652 145590
rect 356612 59152 356664 59158
rect 356612 59094 356664 59100
rect 325884 58744 325936 58750
rect 259458 58712 259514 58721
rect 325884 58686 325936 58692
rect 259458 58647 259514 58656
rect 259472 58614 259500 58647
rect 259460 58608 259512 58614
rect 259460 58550 259512 58556
rect 323308 57928 323360 57934
rect 235998 57896 236054 57905
rect 235998 57831 236054 57840
rect 237378 57896 237434 57905
rect 237378 57831 237434 57840
rect 239218 57896 239274 57905
rect 239218 57831 239274 57840
rect 240138 57896 240194 57905
rect 240138 57831 240194 57840
rect 241610 57896 241666 57905
rect 241610 57831 241666 57840
rect 242898 57896 242954 57905
rect 242898 57831 242954 57840
rect 244370 57896 244426 57905
rect 244370 57831 244426 57840
rect 245290 57896 245346 57905
rect 245290 57831 245346 57840
rect 245658 57896 245714 57905
rect 245658 57831 245714 57840
rect 247038 57896 247094 57905
rect 247038 57831 247094 57840
rect 248602 57896 248658 57905
rect 248602 57831 248658 57840
rect 249798 57896 249854 57905
rect 249798 57831 249854 57840
rect 251178 57896 251234 57905
rect 251178 57831 251234 57840
rect 251362 57896 251418 57905
rect 251362 57831 251418 57840
rect 253386 57896 253442 57905
rect 253386 57831 253442 57840
rect 253938 57896 253994 57905
rect 253938 57831 253994 57840
rect 264978 57896 265034 57905
rect 264978 57831 265034 57840
rect 265898 57896 265954 57905
rect 265898 57831 265954 57840
rect 266358 57896 266414 57905
rect 266358 57831 266414 57840
rect 268474 57896 268530 57905
rect 268474 57831 268530 57840
rect 271234 57896 271290 57905
rect 271234 57831 271290 57840
rect 271878 57896 271934 57905
rect 271878 57831 271934 57840
rect 273258 57896 273314 57905
rect 273258 57831 273314 57840
rect 275466 57896 275522 57905
rect 275466 57831 275522 57840
rect 287610 57896 287666 57905
rect 287610 57831 287666 57840
rect 293314 57896 293370 57905
rect 293314 57831 293370 57840
rect 295890 57896 295946 57905
rect 295890 57831 295946 57840
rect 300858 57896 300914 57905
rect 300858 57831 300914 57840
rect 303434 57896 303490 57905
rect 303434 57831 303490 57840
rect 308494 57896 308550 57905
rect 308494 57831 308550 57840
rect 310978 57896 311034 57905
rect 310978 57831 311034 57840
rect 315762 57896 315818 57905
rect 315762 57831 315764 57840
rect 236012 56438 236040 57831
rect 236000 56432 236052 56438
rect 236000 56374 236052 56380
rect 219992 55820 220044 55826
rect 219992 55762 220044 55768
rect 219808 54868 219860 54874
rect 219808 54810 219860 54816
rect 217140 54800 217192 54806
rect 217140 54742 217192 54748
rect 217048 54732 217100 54738
rect 217048 54674 217100 54680
rect 216036 54664 216088 54670
rect 216036 54606 216088 54612
rect 215116 54528 215168 54534
rect 215116 54470 215168 54476
rect 237392 54330 237420 57831
rect 239232 56506 239260 57831
rect 239220 56500 239272 56506
rect 239220 56442 239272 56448
rect 240152 54398 240180 57831
rect 241624 56574 241652 57831
rect 241612 56568 241664 56574
rect 241612 56510 241664 56516
rect 242912 55214 242940 57831
rect 242900 55208 242952 55214
rect 242900 55150 242952 55156
rect 244384 54534 244412 57831
rect 245304 55962 245332 57831
rect 245292 55956 245344 55962
rect 245292 55898 245344 55904
rect 245672 54602 245700 57831
rect 247052 54670 247080 57831
rect 248616 56030 248644 57831
rect 248604 56024 248656 56030
rect 248604 55966 248656 55972
rect 249812 54738 249840 57831
rect 251192 56098 251220 57831
rect 251180 56092 251232 56098
rect 251180 56034 251232 56040
rect 251376 54806 251404 57831
rect 253400 56166 253428 57831
rect 253388 56160 253440 56166
rect 253388 56102 253440 56108
rect 253952 54874 253980 57831
rect 264992 54942 265020 57831
rect 265912 57254 265940 57831
rect 265900 57248 265952 57254
rect 265900 57190 265952 57196
rect 266372 56234 266400 57831
rect 266450 57624 266506 57633
rect 266450 57559 266506 57568
rect 266360 56228 266412 56234
rect 266360 56170 266412 56176
rect 266464 55010 266492 57559
rect 268488 56302 268516 57831
rect 269118 57624 269174 57633
rect 269118 57559 269174 57568
rect 268476 56296 268528 56302
rect 268476 56238 268528 56244
rect 269132 55078 269160 57559
rect 271248 56370 271276 57831
rect 271236 56364 271288 56370
rect 271236 56306 271288 56312
rect 271892 55146 271920 57831
rect 273272 55758 273300 57831
rect 273350 57624 273406 57633
rect 273350 57559 273406 57568
rect 273260 55752 273312 55758
rect 273260 55694 273312 55700
rect 271880 55140 271932 55146
rect 271880 55082 271932 55088
rect 269120 55072 269172 55078
rect 269120 55014 269172 55020
rect 266452 55004 266504 55010
rect 266452 54946 266504 54952
rect 264980 54936 265032 54942
rect 264980 54878 265032 54884
rect 253940 54868 253992 54874
rect 253940 54810 253992 54816
rect 251364 54800 251416 54806
rect 251364 54742 251416 54748
rect 249800 54732 249852 54738
rect 249800 54674 249852 54680
rect 247040 54664 247092 54670
rect 247040 54606 247092 54612
rect 245660 54596 245712 54602
rect 245660 54538 245712 54544
rect 244372 54528 244424 54534
rect 244372 54470 244424 54476
rect 273364 54466 273392 57559
rect 275480 55894 275508 57831
rect 276018 57624 276074 57633
rect 276018 57559 276074 57568
rect 275468 55888 275520 55894
rect 275468 55830 275520 55836
rect 276032 55185 276060 57559
rect 287624 57322 287652 57831
rect 293328 57390 293356 57831
rect 295904 57526 295932 57831
rect 295892 57520 295944 57526
rect 295892 57462 295944 57468
rect 300872 57458 300900 57831
rect 303448 57594 303476 57831
rect 308508 57730 308536 57831
rect 308496 57724 308548 57730
rect 308496 57666 308548 57672
rect 310992 57662 311020 57831
rect 315816 57831 315818 57840
rect 320914 57896 320970 57905
rect 320914 57831 320970 57840
rect 323306 57896 323308 57905
rect 343180 57928 343232 57934
rect 323360 57896 323362 57905
rect 323306 57831 323362 57840
rect 343178 57896 343180 57905
rect 343232 57896 343234 57905
rect 343178 57831 343234 57840
rect 343454 57896 343510 57905
rect 356716 57866 356744 162250
rect 356808 146266 356836 266358
rect 356900 250646 356928 354962
rect 356992 267034 357020 371826
rect 357084 368014 357112 466278
rect 357256 464976 357308 464982
rect 357256 464918 357308 464924
rect 357164 463616 357216 463622
rect 357164 463558 357216 463564
rect 357176 371074 357204 463558
rect 357268 372026 357296 464918
rect 357808 462936 357860 462942
rect 357808 462878 357860 462884
rect 357820 407794 357848 462878
rect 358084 462120 358136 462126
rect 358084 462062 358136 462068
rect 357992 461984 358044 461990
rect 357992 461926 358044 461932
rect 357900 459468 357952 459474
rect 357900 459410 357952 459416
rect 357808 407788 357860 407794
rect 357808 407730 357860 407736
rect 357256 372020 357308 372026
rect 357256 371962 357308 371968
rect 357256 371816 357308 371822
rect 357256 371758 357308 371764
rect 357164 371068 357216 371074
rect 357164 371010 357216 371016
rect 357072 368008 357124 368014
rect 357072 367950 357124 367956
rect 357268 267238 357296 371758
rect 357440 371680 357492 371686
rect 357440 371622 357492 371628
rect 357348 356040 357400 356046
rect 357348 355982 357400 355988
rect 357360 354822 357388 355982
rect 357348 354816 357400 354822
rect 357348 354758 357400 354764
rect 357256 267232 357308 267238
rect 357256 267174 357308 267180
rect 356980 267028 357032 267034
rect 356980 266970 357032 266976
rect 356992 266422 357020 266970
rect 357072 266484 357124 266490
rect 357072 266426 357124 266432
rect 356980 266416 357032 266422
rect 356980 266358 357032 266364
rect 356888 250640 356940 250646
rect 356888 250582 356940 250588
rect 356796 146260 356848 146266
rect 356796 146202 356848 146208
rect 356900 146062 356928 250582
rect 357084 162858 357112 266426
rect 357360 252362 357388 354758
rect 357452 267734 357480 371622
rect 357912 368082 357940 459410
rect 358004 371142 358032 461926
rect 358096 405006 358124 462062
rect 358084 405000 358136 405006
rect 358084 404942 358136 404948
rect 358084 382288 358136 382294
rect 358084 382230 358136 382236
rect 357992 371136 358044 371142
rect 357992 371078 358044 371084
rect 357900 368076 357952 368082
rect 357900 368018 357952 368024
rect 358096 355366 358124 382230
rect 358084 355360 358136 355366
rect 358084 355302 358136 355308
rect 358096 278050 358124 355302
rect 358084 278044 358136 278050
rect 358084 277986 358136 277992
rect 357452 267706 357756 267734
rect 357728 267306 357756 267706
rect 357716 267300 357768 267306
rect 357716 267242 357768 267248
rect 357360 252334 357664 252362
rect 357636 250578 357664 252334
rect 357624 250572 357676 250578
rect 357624 250514 357676 250520
rect 357532 164212 357584 164218
rect 357532 164154 357584 164160
rect 357072 162852 357124 162858
rect 357072 162794 357124 162800
rect 357544 162178 357572 164154
rect 357532 162172 357584 162178
rect 357532 162114 357584 162120
rect 356888 146056 356940 146062
rect 356888 145998 356940 146004
rect 357544 57934 357572 162114
rect 357636 146130 357664 250514
rect 357728 149025 357756 267242
rect 358096 250510 358124 277986
rect 358084 250504 358136 250510
rect 358084 250446 358136 250452
rect 358096 173194 358124 250446
rect 358084 173188 358136 173194
rect 358084 173130 358136 173136
rect 357714 149016 357770 149025
rect 357714 148951 357770 148960
rect 357624 146124 357676 146130
rect 357624 146066 357676 146072
rect 358096 145586 358124 173130
rect 358084 145580 358136 145586
rect 358084 145522 358136 145528
rect 358084 68468 358136 68474
rect 358084 68410 358136 68416
rect 358096 59362 358124 68410
rect 358084 59356 358136 59362
rect 358084 59298 358136 59304
rect 357532 57928 357584 57934
rect 357532 57870 357584 57876
rect 343454 57831 343456 57840
rect 315764 57802 315816 57808
rect 320928 57798 320956 57831
rect 343508 57831 343510 57840
rect 356704 57860 356756 57866
rect 343456 57802 343508 57808
rect 356704 57802 356756 57808
rect 358188 57798 358216 469882
rect 358280 164082 358308 478382
rect 358268 164076 358320 164082
rect 358268 164018 358320 164024
rect 358372 163946 358400 478450
rect 362224 478304 362276 478310
rect 362224 478246 362276 478252
rect 359832 477488 359884 477494
rect 359832 477430 359884 477436
rect 358452 474292 358504 474298
rect 358452 474234 358504 474240
rect 358464 266966 358492 474234
rect 359464 470416 359516 470422
rect 359464 470358 359516 470364
rect 358544 469124 358596 469130
rect 358544 469066 358596 469072
rect 358556 269113 358584 469066
rect 358728 467764 358780 467770
rect 358728 467706 358780 467712
rect 358634 407824 358690 407833
rect 358634 407759 358690 407768
rect 358542 269104 358598 269113
rect 358542 269039 358598 269048
rect 358452 266960 358504 266966
rect 358452 266902 358504 266908
rect 358360 163940 358412 163946
rect 358360 163882 358412 163888
rect 358648 58750 358676 407759
rect 358740 373522 358768 467706
rect 358820 458312 358872 458318
rect 358820 458254 358872 458260
rect 358832 454753 358860 458254
rect 358818 454744 358874 454753
rect 358874 454702 358952 454730
rect 358818 454679 358874 454688
rect 358728 373516 358780 373522
rect 358728 373458 358780 373464
rect 358818 373280 358874 373289
rect 358818 373215 358874 373224
rect 358832 267170 358860 373215
rect 358924 349625 358952 454702
rect 359094 389328 359150 389337
rect 359094 389263 359150 389272
rect 359004 367804 359056 367810
rect 359004 367746 359056 367752
rect 359016 366382 359044 367746
rect 359004 366376 359056 366382
rect 359004 366318 359056 366324
rect 358910 349616 358966 349625
rect 358910 349551 358966 349560
rect 358820 267164 358872 267170
rect 358820 267106 358872 267112
rect 358832 145654 358860 267106
rect 358924 243817 358952 349551
rect 359016 288425 359044 366318
rect 359108 362234 359136 389263
rect 359476 373386 359504 470358
rect 359648 467560 359700 467566
rect 359648 467502 359700 467508
rect 359556 463276 359608 463282
rect 359556 463218 359608 463224
rect 359464 373380 359516 373386
rect 359464 373322 359516 373328
rect 359568 370734 359596 463218
rect 359660 383586 359688 467502
rect 359740 459332 359792 459338
rect 359740 459274 359792 459280
rect 359752 385014 359780 459274
rect 359844 403646 359872 477430
rect 361028 477148 361080 477154
rect 361028 477090 361080 477096
rect 359924 475924 359976 475930
rect 359924 475866 359976 475872
rect 359936 406434 359964 475866
rect 360016 473204 360068 473210
rect 360016 473146 360068 473152
rect 360028 409154 360056 473146
rect 360936 472932 360988 472938
rect 360936 472874 360988 472880
rect 360844 468580 360896 468586
rect 360844 468522 360896 468528
rect 360752 463684 360804 463690
rect 360752 463626 360804 463632
rect 360200 460964 360252 460970
rect 360200 460906 360252 460912
rect 360016 409148 360068 409154
rect 360016 409090 360068 409096
rect 359924 406428 359976 406434
rect 359924 406370 359976 406376
rect 359832 403640 359884 403646
rect 359832 403582 359884 403588
rect 360014 393816 360070 393825
rect 360014 393751 360070 393760
rect 359922 392184 359978 392193
rect 359922 392119 359978 392128
rect 359830 390824 359886 390833
rect 359830 390759 359886 390768
rect 359740 385008 359792 385014
rect 359740 384950 359792 384956
rect 359648 383580 359700 383586
rect 359648 383522 359700 383528
rect 359556 370728 359608 370734
rect 359556 370670 359608 370676
rect 359464 369912 359516 369918
rect 359464 369854 359516 369860
rect 359476 364334 359504 369854
rect 359556 369164 359608 369170
rect 359556 369106 359608 369112
rect 359200 364306 359504 364334
rect 359096 362228 359148 362234
rect 359096 362170 359148 362176
rect 359200 360194 359228 364306
rect 359464 362228 359516 362234
rect 359464 362170 359516 362176
rect 359188 360188 359240 360194
rect 359188 360130 359240 360136
rect 359200 354674 359228 360130
rect 359280 359508 359332 359514
rect 359280 359450 359332 359456
rect 359292 358086 359320 359450
rect 359476 358154 359504 362170
rect 359464 358148 359516 358154
rect 359464 358090 359516 358096
rect 359280 358080 359332 358086
rect 359280 358022 359332 358028
rect 359108 354646 359228 354674
rect 359108 289377 359136 354646
rect 359188 353320 359240 353326
rect 359188 353262 359240 353268
rect 359094 289368 359150 289377
rect 359094 289303 359150 289312
rect 359002 288416 359058 288425
rect 359002 288351 359058 288360
rect 359002 283112 359058 283121
rect 359002 283047 359058 283056
rect 358910 243808 358966 243817
rect 358910 243743 358966 243752
rect 358910 183560 358966 183569
rect 358910 183495 358966 183504
rect 358924 182753 358952 183495
rect 358910 182744 358966 182753
rect 358910 182679 358966 182688
rect 358820 145648 358872 145654
rect 358820 145590 358872 145596
rect 358728 145580 358780 145586
rect 358728 145522 358780 145528
rect 358740 68474 358768 145522
rect 358924 78305 358952 182679
rect 359016 178673 359044 283047
rect 359108 184929 359136 289303
rect 359200 283121 359228 353262
rect 359292 286385 359320 358022
rect 359278 286376 359334 286385
rect 359278 286311 359334 286320
rect 359186 283112 359242 283121
rect 359186 283047 359242 283056
rect 359094 184920 359150 184929
rect 359094 184855 359150 184864
rect 359002 178664 359058 178673
rect 359002 178599 359058 178608
rect 358910 78296 358966 78305
rect 358910 78231 358966 78240
rect 359016 74089 359044 178599
rect 359108 79937 359136 184855
rect 359292 181393 359320 286311
rect 359476 284889 359504 358090
rect 359568 354006 359596 369106
rect 359844 359514 359872 390759
rect 359936 367810 359964 392119
rect 360028 370530 360056 393751
rect 360106 388104 360162 388113
rect 360106 388039 360162 388048
rect 360016 370524 360068 370530
rect 360016 370466 360068 370472
rect 360028 369918 360056 370466
rect 360016 369912 360068 369918
rect 360016 369854 360068 369860
rect 360120 369170 360148 388039
rect 360212 383654 360240 460906
rect 360200 383648 360252 383654
rect 360200 383590 360252 383596
rect 360212 382294 360240 383590
rect 360200 382288 360252 382294
rect 360200 382230 360252 382236
rect 360764 371958 360792 463626
rect 360752 371952 360804 371958
rect 360752 371894 360804 371900
rect 360200 371272 360252 371278
rect 360200 371214 360252 371220
rect 360108 369164 360160 369170
rect 360108 369106 360160 369112
rect 359924 367804 359976 367810
rect 359924 367746 359976 367752
rect 359832 359508 359884 359514
rect 359832 359450 359884 359456
rect 359556 354000 359608 354006
rect 359556 353942 359608 353948
rect 359568 353326 359596 353942
rect 359556 353320 359608 353326
rect 359556 353262 359608 353268
rect 359554 288416 359610 288425
rect 359554 288351 359610 288360
rect 359462 284880 359518 284889
rect 359462 284815 359518 284824
rect 359370 243808 359426 243817
rect 359370 243743 359426 243752
rect 359278 181384 359334 181393
rect 359278 181319 359334 181328
rect 359292 180794 359320 181319
rect 359200 180766 359320 180794
rect 359094 79928 359150 79937
rect 359094 79863 359150 79872
rect 359200 76945 359228 180766
rect 359278 179480 359334 179489
rect 359278 179415 359334 179424
rect 359186 76936 359242 76945
rect 359186 76871 359242 76880
rect 359292 75449 359320 179415
rect 359384 139369 359412 243743
rect 359476 179489 359504 284815
rect 359568 183569 359596 288351
rect 360212 267374 360240 371214
rect 360200 267368 360252 267374
rect 360200 267310 360252 267316
rect 359554 183560 359610 183569
rect 359554 183495 359610 183504
rect 359462 179480 359518 179489
rect 359462 179415 359518 179424
rect 360212 164218 360240 267310
rect 360200 164212 360252 164218
rect 360200 164154 360252 164160
rect 359370 139360 359426 139369
rect 359370 139295 359426 139304
rect 359278 75440 359334 75449
rect 359278 75375 359334 75384
rect 359002 74080 359058 74089
rect 359002 74015 359058 74024
rect 358728 68468 358780 68474
rect 358728 68410 358780 68416
rect 358636 58744 358688 58750
rect 358636 58686 358688 58692
rect 360856 57866 360884 468522
rect 360948 162586 360976 472874
rect 361040 268734 361068 477090
rect 361212 471572 361264 471578
rect 361212 471514 361264 471520
rect 361120 460828 361172 460834
rect 361120 460770 361172 460776
rect 361028 268728 361080 268734
rect 361028 268670 361080 268676
rect 361132 266937 361160 460770
rect 361224 278730 361252 471514
rect 361304 471232 361356 471238
rect 361304 471174 361356 471180
rect 361316 369034 361344 471174
rect 361396 467492 361448 467498
rect 361396 467434 361448 467440
rect 361408 373794 361436 467434
rect 362040 464704 362092 464710
rect 362040 464646 362092 464652
rect 361488 463548 361540 463554
rect 361488 463490 361540 463496
rect 361396 373788 361448 373794
rect 361396 373730 361448 373736
rect 361500 370870 361528 463490
rect 362052 410582 362080 464646
rect 362132 459264 362184 459270
rect 362132 459206 362184 459212
rect 362040 410576 362092 410582
rect 362040 410518 362092 410524
rect 361488 370864 361540 370870
rect 361488 370806 361540 370812
rect 362144 370326 362172 459206
rect 362132 370320 362184 370326
rect 362132 370262 362184 370268
rect 361304 369028 361356 369034
rect 361304 368970 361356 368976
rect 361212 278724 361264 278730
rect 361212 278666 361264 278672
rect 361118 266928 361174 266937
rect 361118 266863 361174 266872
rect 360936 162580 360988 162586
rect 360936 162522 360988 162528
rect 362236 59430 362264 478246
rect 363604 478236 363656 478242
rect 363604 478178 363656 478184
rect 362408 475448 362460 475454
rect 362408 475390 362460 475396
rect 362316 471300 362368 471306
rect 362316 471242 362368 471248
rect 362224 59424 362276 59430
rect 362224 59366 362276 59372
rect 360844 57860 360896 57866
rect 360844 57802 360896 57808
rect 320916 57792 320968 57798
rect 320916 57734 320968 57740
rect 358176 57792 358228 57798
rect 358176 57734 358228 57740
rect 310980 57656 311032 57662
rect 310980 57598 311032 57604
rect 362328 57594 362356 471242
rect 362420 162178 362448 475390
rect 362776 474632 362828 474638
rect 362776 474574 362828 474580
rect 362592 471776 362644 471782
rect 362592 471718 362644 471724
rect 362500 463004 362552 463010
rect 362500 462946 362552 462952
rect 362512 163878 362540 462946
rect 362604 267306 362632 471718
rect 362684 470212 362736 470218
rect 362684 470154 362736 470160
rect 362696 268394 362724 470154
rect 362788 367946 362816 474574
rect 362868 473068 362920 473074
rect 362868 473010 362920 473016
rect 362880 373590 362908 473010
rect 363512 464636 363564 464642
rect 363512 464578 363564 464584
rect 362960 461032 363012 461038
rect 362960 460974 363012 460980
rect 362868 373584 362920 373590
rect 362868 373526 362920 373532
rect 362776 367940 362828 367946
rect 362776 367882 362828 367888
rect 362972 356046 363000 460974
rect 363524 411942 363552 464578
rect 363512 411936 363564 411942
rect 363512 411878 363564 411884
rect 363052 371340 363104 371346
rect 363052 371282 363104 371288
rect 362960 356040 363012 356046
rect 362960 355982 363012 355988
rect 362684 268388 362736 268394
rect 362684 268330 362736 268336
rect 362592 267300 362644 267306
rect 362592 267242 362644 267248
rect 363064 266490 363092 371282
rect 363052 266484 363104 266490
rect 363052 266426 363104 266432
rect 362500 163872 362552 163878
rect 362500 163814 362552 163820
rect 362408 162172 362460 162178
rect 362408 162114 362460 162120
rect 363616 58886 363644 478178
rect 363788 476876 363840 476882
rect 363788 476818 363840 476824
rect 363696 467220 363748 467226
rect 363696 467162 363748 467168
rect 363604 58880 363656 58886
rect 363604 58822 363656 58828
rect 363708 57730 363736 467162
rect 363800 162450 363828 476818
rect 365168 475516 365220 475522
rect 365168 475458 365220 475464
rect 364984 472796 365036 472802
rect 364984 472738 365036 472744
rect 364156 470348 364208 470354
rect 364156 470290 364208 470296
rect 364064 469192 364116 469198
rect 364064 469134 364116 469140
rect 363972 461848 364024 461854
rect 363972 461790 364024 461796
rect 363880 460760 363932 460766
rect 363880 460702 363932 460708
rect 363892 267374 363920 460702
rect 363984 269482 364012 461790
rect 364076 373318 364104 469134
rect 364168 374066 364196 470290
rect 364892 463480 364944 463486
rect 364892 463422 364944 463428
rect 364248 459400 364300 459406
rect 364248 459342 364300 459348
rect 364156 374060 364208 374066
rect 364156 374002 364208 374008
rect 364064 373312 364116 373318
rect 364064 373254 364116 373260
rect 364260 367878 364288 459342
rect 364800 459128 364852 459134
rect 364800 459070 364852 459076
rect 364812 374134 364840 459070
rect 364800 374128 364852 374134
rect 364800 374070 364852 374076
rect 364904 370802 364932 463422
rect 364892 370796 364944 370802
rect 364892 370738 364944 370744
rect 364248 367872 364300 367878
rect 364248 367814 364300 367820
rect 363972 269476 364024 269482
rect 363972 269418 364024 269424
rect 363880 267368 363932 267374
rect 363880 267310 363932 267316
rect 363788 162444 363840 162450
rect 363788 162386 363840 162392
rect 364996 57934 365024 472738
rect 365076 470008 365128 470014
rect 365076 469950 365128 469956
rect 365088 70378 365116 469950
rect 365180 162858 365208 475458
rect 365352 471844 365404 471850
rect 365352 471786 365404 471792
rect 365260 463140 365312 463146
rect 365260 463082 365312 463088
rect 365272 164286 365300 463082
rect 365364 269142 365392 471786
rect 365444 467424 365496 467430
rect 365444 467366 365496 467372
rect 365352 269136 365404 269142
rect 365352 269078 365404 269084
rect 365456 267034 365484 467366
rect 365536 466132 365588 466138
rect 365536 466074 365588 466080
rect 365548 368150 365576 466074
rect 365628 464908 365680 464914
rect 365628 464850 365680 464856
rect 365640 369306 365668 464850
rect 366272 464840 366324 464846
rect 366272 464782 366324 464788
rect 366180 461916 366232 461922
rect 366180 461858 366232 461864
rect 366192 371006 366220 461858
rect 366180 371000 366232 371006
rect 366180 370942 366232 370948
rect 365628 369300 365680 369306
rect 365628 369242 365680 369248
rect 366284 369238 366312 464782
rect 366272 369232 366324 369238
rect 366272 369174 366324 369180
rect 365536 368144 365588 368150
rect 365536 368086 365588 368092
rect 365444 267028 365496 267034
rect 365444 266970 365496 266976
rect 365260 164280 365312 164286
rect 365260 164222 365312 164228
rect 365168 162852 365220 162858
rect 365168 162794 365220 162800
rect 365076 70372 365128 70378
rect 365076 70314 365128 70320
rect 364984 57928 365036 57934
rect 364984 57870 365036 57876
rect 363696 57724 363748 57730
rect 363696 57666 363748 57672
rect 303436 57588 303488 57594
rect 303436 57530 303488 57536
rect 362316 57588 362368 57594
rect 362316 57530 362368 57536
rect 300860 57452 300912 57458
rect 300860 57394 300912 57400
rect 293316 57384 293368 57390
rect 293316 57326 293368 57332
rect 287612 57316 287664 57322
rect 287612 57258 287664 57264
rect 276018 55176 276074 55185
rect 276018 55111 276074 55120
rect 273352 54460 273404 54466
rect 273352 54402 273404 54408
rect 240140 54392 240192 54398
rect 240140 54334 240192 54340
rect 214564 54324 214616 54330
rect 214564 54266 214616 54272
rect 237380 54324 237432 54330
rect 237380 54266 237432 54272
rect 136454 4040 136510 4049
rect 136454 3975 136510 3984
rect 132958 3904 133014 3913
rect 132958 3839 133014 3848
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 57244 3460 57296 3466
rect 57244 3402 57296 3408
rect 125876 3460 125928 3466
rect 125876 3402 125928 3408
rect 584 480 612 3402
rect 125888 480 125916 3402
rect 129370 3360 129426 3369
rect 129370 3295 129426 3304
rect 129384 480 129412 3295
rect 132972 480 133000 3839
rect 136468 480 136496 3975
rect 147126 3768 147182 3777
rect 147126 3703 147182 3712
rect 143538 3632 143594 3641
rect 143538 3567 143594 3576
rect 140042 3224 140098 3233
rect 140042 3159 140098 3168
rect 140056 480 140084 3159
rect 143552 480 143580 3567
rect 147140 480 147168 3703
rect 150622 3496 150678 3505
rect 366376 3466 366404 480791
rect 366456 478372 366508 478378
rect 366456 478314 366508 478320
rect 366468 58818 366496 478314
rect 373264 478168 373316 478174
rect 373264 478110 373316 478116
rect 371056 477216 371108 477222
rect 371056 477158 371108 477164
rect 369492 477012 369544 477018
rect 369492 476954 369544 476960
rect 368112 476944 368164 476950
rect 368112 476886 368164 476892
rect 367008 475788 367060 475794
rect 367008 475730 367060 475736
rect 366732 474020 366784 474026
rect 366732 473962 366784 473968
rect 366548 468716 366600 468722
rect 366548 468658 366600 468664
rect 366560 162654 366588 468658
rect 366640 465928 366692 465934
rect 366640 465870 366692 465876
rect 366652 163538 366680 465870
rect 366744 173874 366772 473962
rect 366824 470144 366876 470150
rect 366824 470086 366876 470092
rect 366836 267102 366864 470086
rect 366916 459060 366968 459066
rect 366916 459002 366968 459008
rect 366928 268598 366956 459002
rect 367020 374338 367048 475730
rect 367744 471436 367796 471442
rect 367744 471378 367796 471384
rect 367652 460896 367704 460902
rect 367652 460838 367704 460844
rect 367560 459196 367612 459202
rect 367560 459138 367612 459144
rect 367008 374332 367060 374338
rect 367008 374274 367060 374280
rect 367572 373454 367600 459138
rect 367560 373448 367612 373454
rect 367560 373390 367612 373396
rect 367664 373250 367692 460838
rect 367652 373244 367704 373250
rect 367652 373186 367704 373192
rect 366916 268592 366968 268598
rect 366916 268534 366968 268540
rect 366824 267096 366876 267102
rect 366824 267038 366876 267044
rect 366732 173868 366784 173874
rect 366732 173810 366784 173816
rect 366640 163532 366692 163538
rect 366640 163474 366692 163480
rect 366548 162648 366600 162654
rect 366548 162590 366600 162596
rect 367756 162110 367784 471378
rect 368020 468784 368072 468790
rect 368020 468726 368072 468732
rect 367836 468648 367888 468654
rect 367836 468590 367888 468596
rect 367848 164014 367876 468590
rect 367928 460624 367980 460630
rect 367928 460566 367980 460572
rect 367836 164008 367888 164014
rect 367836 163950 367888 163956
rect 367940 163674 367968 460566
rect 368032 175234 368060 468726
rect 368124 268802 368152 476886
rect 369124 475380 369176 475386
rect 369124 475322 369176 475328
rect 368204 474156 368256 474162
rect 368204 474098 368256 474104
rect 368112 268796 368164 268802
rect 368112 268738 368164 268744
rect 368216 267510 368244 474098
rect 368296 471980 368348 471986
rect 368296 471922 368348 471928
rect 368308 369102 368336 471922
rect 368388 466064 368440 466070
rect 368388 466006 368440 466012
rect 368400 372094 368428 466006
rect 369032 464772 369084 464778
rect 369032 464714 369084 464720
rect 368940 463344 368992 463350
rect 368940 463286 368992 463292
rect 368388 372088 368440 372094
rect 368388 372030 368440 372036
rect 368952 370938 368980 463286
rect 368940 370932 368992 370938
rect 368940 370874 368992 370880
rect 369044 370598 369072 464714
rect 369032 370592 369084 370598
rect 369032 370534 369084 370540
rect 368296 369096 368348 369102
rect 368296 369038 368348 369044
rect 368388 368076 368440 368082
rect 368388 368018 368440 368024
rect 368296 367872 368348 367878
rect 368296 367814 368348 367820
rect 368204 267504 368256 267510
rect 368204 267446 368256 267452
rect 368308 251054 368336 367814
rect 368400 251122 368428 368018
rect 368388 251116 368440 251122
rect 368388 251058 368440 251064
rect 368296 251048 368348 251054
rect 368296 250990 368348 250996
rect 368020 175228 368072 175234
rect 368020 175170 368072 175176
rect 367928 163668 367980 163674
rect 367928 163610 367980 163616
rect 369136 162246 369164 475322
rect 369216 474088 369268 474094
rect 369216 474030 369268 474036
rect 369228 162790 369256 474030
rect 369308 465860 369360 465866
rect 369308 465802 369360 465808
rect 369320 164121 369348 465802
rect 369400 460420 369452 460426
rect 369400 460362 369452 460368
rect 369412 164354 369440 460362
rect 369504 267646 369532 476954
rect 369676 474496 369728 474502
rect 369676 474438 369728 474444
rect 369584 474360 369636 474366
rect 369584 474302 369636 474308
rect 369596 268530 369624 474302
rect 369688 374270 369716 474438
rect 370688 472864 370740 472870
rect 370688 472806 370740 472812
rect 370504 467152 370556 467158
rect 370504 467094 370556 467100
rect 369860 466268 369912 466274
rect 369860 466210 369912 466216
rect 369676 374264 369728 374270
rect 369676 374206 369728 374212
rect 369872 373994 369900 466210
rect 370412 464568 370464 464574
rect 370412 464510 370464 464516
rect 370320 463412 370372 463418
rect 370320 463354 370372 463360
rect 369780 373966 369900 373994
rect 369676 372700 369728 372706
rect 369676 372642 369728 372648
rect 369584 268524 369636 268530
rect 369584 268466 369636 268472
rect 369492 267640 369544 267646
rect 369492 267582 369544 267588
rect 369688 262206 369716 372642
rect 369780 372450 369808 373966
rect 369860 372564 369912 372570
rect 369860 372506 369912 372512
rect 369872 372450 369900 372506
rect 369780 372422 369900 372450
rect 369676 262200 369728 262206
rect 369676 262142 369728 262148
rect 369780 251190 369808 372422
rect 370332 368966 370360 463354
rect 370424 369578 370452 464510
rect 370412 369572 370464 369578
rect 370412 369514 370464 369520
rect 370320 368960 370372 368966
rect 370320 368902 370372 368908
rect 370412 367940 370464 367946
rect 370412 367882 370464 367888
rect 370318 269376 370374 269385
rect 370318 269311 370374 269320
rect 370228 265940 370280 265946
rect 370228 265882 370280 265888
rect 369768 251184 369820 251190
rect 369768 251126 369820 251132
rect 369400 164348 369452 164354
rect 369400 164290 369452 164296
rect 369306 164112 369362 164121
rect 369306 164047 369362 164056
rect 369216 162784 369268 162790
rect 369216 162726 369268 162732
rect 369124 162240 369176 162246
rect 369124 162182 369176 162188
rect 367744 162104 367796 162110
rect 367744 162046 367796 162052
rect 370240 148510 370268 265882
rect 370228 148504 370280 148510
rect 370228 148446 370280 148452
rect 370332 148442 370360 269311
rect 370424 267578 370452 367882
rect 370412 267572 370464 267578
rect 370412 267514 370464 267520
rect 370412 251184 370464 251190
rect 370412 251126 370464 251132
rect 370424 250646 370452 251126
rect 370412 250640 370464 250646
rect 370412 250582 370464 250588
rect 370424 160750 370452 250582
rect 370412 160744 370464 160750
rect 370412 160686 370464 160692
rect 370320 148436 370372 148442
rect 370320 148378 370372 148384
rect 366456 58812 366508 58818
rect 366456 58754 366508 58760
rect 370516 57322 370544 467094
rect 370596 465724 370648 465730
rect 370596 465666 370648 465672
rect 370608 57458 370636 465666
rect 370700 162722 370728 472806
rect 370872 468920 370924 468926
rect 370872 468862 370924 468868
rect 370780 460556 370832 460562
rect 370780 460498 370832 460504
rect 370792 163742 370820 460498
rect 370884 267238 370912 468862
rect 370964 468852 371016 468858
rect 370964 468794 371016 468800
rect 370976 269278 371004 468794
rect 371068 374610 371096 477158
rect 371792 475720 371844 475726
rect 371792 475662 371844 475668
rect 371700 468444 371752 468450
rect 371700 468386 371752 468392
rect 371056 374604 371108 374610
rect 371056 374546 371108 374552
rect 371606 372736 371662 372745
rect 371606 372671 371662 372680
rect 371056 371748 371108 371754
rect 371056 371690 371108 371696
rect 371068 371550 371096 371690
rect 371148 371612 371200 371618
rect 371148 371554 371200 371560
rect 371056 371544 371108 371550
rect 371056 371486 371108 371492
rect 370964 269272 371016 269278
rect 370964 269214 371016 269220
rect 370872 267232 370924 267238
rect 370872 267174 370924 267180
rect 371068 265810 371096 371486
rect 371056 265804 371108 265810
rect 371056 265746 371108 265752
rect 371160 265674 371188 371554
rect 371148 265668 371200 265674
rect 371148 265610 371200 265616
rect 371620 265577 371648 372671
rect 371712 369374 371740 468386
rect 371804 373726 371832 475662
rect 372160 474224 372212 474230
rect 372160 474166 372212 474172
rect 371884 472660 371936 472666
rect 371884 472602 371936 472608
rect 371792 373720 371844 373726
rect 371792 373662 371844 373668
rect 371700 369368 371752 369374
rect 371700 369310 371752 369316
rect 371792 369232 371844 369238
rect 371792 369174 371844 369180
rect 371700 269340 371752 269346
rect 371700 269282 371752 269288
rect 371606 265568 371662 265577
rect 371606 265503 371662 265512
rect 370964 251116 371016 251122
rect 370964 251058 371016 251064
rect 370872 251048 370924 251054
rect 370872 250990 370924 250996
rect 370884 250510 370912 250990
rect 370976 250578 371004 251058
rect 370964 250572 371016 250578
rect 370964 250514 371016 250520
rect 370872 250504 370924 250510
rect 370872 250446 370924 250452
rect 370780 163736 370832 163742
rect 370780 163678 370832 163684
rect 370688 162716 370740 162722
rect 370688 162658 370740 162664
rect 370884 159390 370912 250446
rect 370872 159384 370924 159390
rect 370872 159326 370924 159332
rect 370976 148481 371004 250514
rect 371712 160818 371740 269282
rect 371804 265169 371832 369174
rect 371790 265160 371846 265169
rect 371790 265095 371846 265104
rect 371700 160812 371752 160818
rect 371700 160754 371752 160760
rect 370962 148472 371018 148481
rect 370962 148407 371018 148416
rect 371896 57526 371924 472602
rect 371976 470076 372028 470082
rect 371976 470018 372028 470024
rect 371988 162518 372016 470018
rect 372068 463072 372120 463078
rect 372068 463014 372120 463020
rect 372080 163606 372108 463014
rect 372172 268462 372200 474166
rect 372620 473136 372672 473142
rect 372620 473078 372672 473084
rect 372252 473000 372304 473006
rect 372252 472942 372304 472948
rect 372160 268456 372212 268462
rect 372160 268398 372212 268404
rect 372264 267714 372292 472942
rect 372436 469056 372488 469062
rect 372436 468998 372488 469004
rect 372344 458992 372396 458998
rect 372344 458934 372396 458940
rect 372252 267708 372304 267714
rect 372252 267650 372304 267656
rect 372356 267170 372384 458934
rect 372448 374202 372476 468998
rect 372436 374196 372488 374202
rect 372436 374138 372488 374144
rect 372632 373862 372660 473078
rect 373172 468988 373224 468994
rect 373172 468930 373224 468936
rect 373078 374096 373134 374105
rect 373078 374031 373134 374040
rect 372620 373856 372672 373862
rect 372620 373798 372672 373804
rect 372528 372632 372580 372638
rect 372528 372574 372580 372580
rect 372540 269346 372568 372574
rect 372988 371816 373040 371822
rect 372988 371758 373040 371764
rect 373000 371482 373028 371758
rect 372988 371476 373040 371482
rect 372988 371418 373040 371424
rect 372528 269340 372580 269346
rect 372528 269282 372580 269288
rect 372528 269204 372580 269210
rect 372528 269146 372580 269152
rect 372344 267164 372396 267170
rect 372344 267106 372396 267112
rect 372436 265804 372488 265810
rect 372436 265746 372488 265752
rect 372344 265668 372396 265674
rect 372344 265610 372396 265616
rect 372068 163600 372120 163606
rect 372068 163542 372120 163548
rect 371976 162512 372028 162518
rect 371976 162454 372028 162460
rect 372252 159384 372304 159390
rect 372252 159326 372304 159332
rect 371976 148504 372028 148510
rect 371976 148446 372028 148452
rect 371884 57520 371936 57526
rect 371884 57462 371936 57468
rect 370596 57452 370648 57458
rect 370596 57394 370648 57400
rect 370504 57316 370556 57322
rect 370504 57258 370556 57264
rect 371988 55894 372016 148446
rect 372264 56438 372292 159326
rect 372356 148578 372384 265610
rect 372344 148572 372396 148578
rect 372344 148514 372396 148520
rect 372448 144906 372476 265746
rect 372540 145625 372568 269146
rect 373000 265946 373028 371418
rect 373092 269074 373120 374031
rect 373184 369646 373212 468930
rect 373172 369640 373224 369646
rect 373172 369582 373224 369588
rect 373172 354000 373224 354006
rect 373172 353942 373224 353948
rect 373184 269822 373212 353942
rect 373172 269816 373224 269822
rect 373172 269758 373224 269764
rect 373080 269068 373132 269074
rect 373080 269010 373132 269016
rect 373172 268184 373224 268190
rect 373172 268126 373224 268132
rect 373184 267578 373212 268126
rect 373172 267572 373224 267578
rect 373172 267514 373224 267520
rect 372988 265940 373040 265946
rect 372988 265882 373040 265888
rect 373184 163198 373212 267514
rect 373172 163192 373224 163198
rect 373172 163134 373224 163140
rect 372526 145616 372582 145625
rect 372526 145551 372582 145560
rect 372436 144900 372488 144906
rect 372436 144842 372488 144848
rect 373276 58954 373304 478110
rect 375196 477420 375248 477426
rect 375196 477362 375248 477368
rect 374920 475584 374972 475590
rect 374920 475526 374972 475532
rect 374644 469872 374696 469878
rect 374644 469814 374696 469820
rect 373356 467288 373408 467294
rect 373356 467230 373408 467236
rect 373368 162382 373396 467230
rect 373816 466200 373868 466206
rect 373816 466142 373868 466148
rect 373448 465792 373500 465798
rect 373448 465734 373500 465740
rect 373460 164422 373488 465734
rect 373632 461712 373684 461718
rect 373632 461654 373684 461660
rect 373540 460488 373592 460494
rect 373540 460430 373592 460436
rect 373448 164416 373500 164422
rect 373448 164358 373500 164364
rect 373552 163810 373580 460430
rect 373644 266830 373672 461654
rect 373724 460692 373776 460698
rect 373724 460634 373776 460640
rect 373736 374542 373764 460634
rect 373724 374536 373776 374542
rect 373724 374478 373776 374484
rect 373724 373856 373776 373862
rect 373724 373798 373776 373804
rect 373736 372706 373764 373798
rect 373724 372700 373776 372706
rect 373724 372642 373776 372648
rect 373828 371793 373856 466142
rect 374460 463208 374512 463214
rect 374460 463150 374512 463156
rect 374000 462052 374052 462058
rect 374000 461994 374052 462000
rect 373908 407856 373960 407862
rect 373908 407798 373960 407804
rect 373814 371784 373870 371793
rect 373814 371719 373870 371728
rect 373816 370660 373868 370666
rect 373816 370602 373868 370608
rect 373724 269068 373776 269074
rect 373724 269010 373776 269016
rect 373736 268258 373764 269010
rect 373724 268252 373776 268258
rect 373724 268194 373776 268200
rect 373632 266824 373684 266830
rect 373632 266766 373684 266772
rect 373540 163804 373592 163810
rect 373540 163746 373592 163752
rect 373736 163062 373764 268194
rect 373828 267986 373856 370602
rect 373920 369850 373948 407798
rect 374012 372638 374040 461994
rect 374000 372632 374052 372638
rect 374000 372574 374052 372580
rect 374000 370592 374052 370598
rect 374000 370534 374052 370540
rect 373908 369844 373960 369850
rect 373908 369786 373960 369792
rect 374012 269210 374040 370534
rect 374472 369782 374500 463150
rect 374460 369776 374512 369782
rect 374460 369718 374512 369724
rect 374552 369436 374604 369442
rect 374552 369378 374604 369384
rect 374460 269816 374512 269822
rect 374460 269758 374512 269764
rect 374472 269414 374500 269758
rect 374460 269408 374512 269414
rect 374380 269356 374460 269362
rect 374380 269350 374512 269356
rect 374380 269334 374500 269350
rect 374000 269204 374052 269210
rect 374000 269146 374052 269152
rect 373816 267980 373868 267986
rect 373816 267922 373868 267928
rect 374276 267980 374328 267986
rect 374276 267922 374328 267928
rect 373908 266212 373960 266218
rect 373908 266154 373960 266160
rect 373814 265568 373870 265577
rect 373814 265503 373870 265512
rect 373724 163056 373776 163062
rect 373724 162998 373776 163004
rect 373356 162376 373408 162382
rect 373356 162318 373408 162324
rect 373828 160886 373856 265503
rect 373816 160880 373868 160886
rect 373816 160822 373868 160828
rect 373632 160812 373684 160818
rect 373632 160754 373684 160760
rect 373264 58948 373316 58954
rect 373264 58890 373316 58896
rect 372252 56432 372304 56438
rect 372252 56374 372304 56380
rect 371976 55888 372028 55894
rect 371976 55830 372028 55836
rect 373644 54466 373672 160754
rect 373724 148912 373776 148918
rect 373724 148854 373776 148860
rect 373736 54534 373764 148854
rect 373920 144906 373948 266154
rect 374092 265260 374144 265266
rect 374092 265202 374144 265208
rect 373908 144900 373960 144906
rect 373908 144842 373960 144848
rect 374104 144838 374132 265202
rect 374184 163192 374236 163198
rect 374184 163134 374236 163140
rect 374092 144832 374144 144838
rect 374092 144774 374144 144780
rect 374196 55078 374224 163134
rect 374288 145926 374316 267922
rect 374380 147694 374408 269334
rect 374460 269204 374512 269210
rect 374460 269146 374512 269152
rect 374472 268870 374500 269146
rect 374460 268864 374512 268870
rect 374460 268806 374512 268812
rect 374564 251190 374592 369378
rect 374552 251184 374604 251190
rect 374552 251126 374604 251132
rect 374564 238754 374592 251126
rect 374472 238726 374592 238754
rect 374368 147688 374420 147694
rect 374368 147630 374420 147636
rect 374472 146305 374500 238726
rect 374552 160744 374604 160750
rect 374552 160686 374604 160692
rect 374458 146296 374514 146305
rect 374458 146231 374514 146240
rect 374276 145920 374328 145926
rect 374276 145862 374328 145868
rect 374288 144702 374316 145862
rect 374276 144696 374328 144702
rect 374276 144638 374328 144644
rect 374564 56506 374592 160686
rect 374656 57662 374684 469814
rect 374736 460216 374788 460222
rect 374736 460158 374788 460164
rect 374748 162042 374776 460158
rect 374828 458924 374880 458930
rect 374828 458866 374880 458872
rect 374840 162314 374868 458866
rect 374932 267442 374960 475526
rect 375104 474564 375156 474570
rect 375104 474506 375156 474512
rect 375012 471504 375064 471510
rect 375012 471446 375064 471452
rect 375024 269210 375052 471446
rect 375116 371210 375144 474506
rect 375208 375018 375236 477362
rect 377312 477352 377364 477358
rect 377312 477294 377364 477300
rect 376484 475652 376536 475658
rect 376484 475594 376536 475600
rect 376024 468512 376076 468518
rect 376024 468454 376076 468460
rect 375380 464432 375432 464438
rect 375380 464374 375432 464380
rect 375196 375012 375248 375018
rect 375196 374954 375248 374960
rect 375392 374746 375420 464374
rect 375932 405680 375984 405686
rect 375932 405622 375984 405628
rect 375380 374740 375432 374746
rect 375380 374682 375432 374688
rect 375392 374626 375420 374682
rect 375300 374598 375420 374626
rect 375196 372632 375248 372638
rect 375196 372574 375248 372580
rect 375208 372502 375236 372574
rect 375196 372496 375248 372502
rect 375196 372438 375248 372444
rect 375196 371884 375248 371890
rect 375196 371826 375248 371832
rect 375208 371414 375236 371826
rect 375196 371408 375248 371414
rect 375196 371350 375248 371356
rect 375104 371204 375156 371210
rect 375104 371146 375156 371152
rect 375104 368008 375156 368014
rect 375104 367950 375156 367956
rect 375012 269204 375064 269210
rect 375012 269146 375064 269152
rect 374920 267436 374972 267442
rect 374920 267378 374972 267384
rect 375116 263566 375144 367950
rect 375208 266014 375236 371350
rect 375196 266008 375248 266014
rect 375196 265950 375248 265956
rect 375104 263560 375156 263566
rect 375104 263502 375156 263508
rect 375116 263106 375144 263502
rect 374932 263078 375144 263106
rect 374932 164218 374960 263078
rect 375208 258074 375236 265950
rect 375300 265470 375328 374598
rect 375944 370666 375972 405622
rect 375932 370660 375984 370666
rect 375932 370602 375984 370608
rect 375932 369368 375984 369374
rect 375932 369310 375984 369316
rect 375838 266384 375894 266393
rect 375838 266319 375894 266328
rect 375288 265464 375340 265470
rect 375288 265406 375340 265412
rect 375024 258046 375236 258074
rect 374920 164212 374972 164218
rect 374920 164154 374972 164160
rect 374920 163056 374972 163062
rect 374920 162998 374972 163004
rect 374828 162308 374880 162314
rect 374828 162250 374880 162256
rect 374736 162036 374788 162042
rect 374736 161978 374788 161984
rect 374736 160880 374788 160886
rect 374736 160822 374788 160828
rect 374644 57656 374696 57662
rect 374644 57598 374696 57604
rect 374552 56500 374604 56506
rect 374552 56442 374604 56448
rect 374184 55072 374236 55078
rect 374184 55014 374236 55020
rect 374748 55010 374776 160822
rect 374736 55004 374788 55010
rect 374736 54946 374788 54952
rect 374932 54942 374960 162998
rect 375024 148918 375052 258046
rect 375748 164212 375800 164218
rect 375748 164154 375800 164160
rect 375288 163192 375340 163198
rect 375288 163134 375340 163140
rect 375300 162994 375328 163134
rect 375288 162988 375340 162994
rect 375288 162930 375340 162936
rect 375760 162926 375788 164154
rect 375748 162920 375800 162926
rect 375748 162862 375800 162868
rect 375012 148912 375064 148918
rect 375012 148854 375064 148860
rect 375012 148572 375064 148578
rect 375012 148514 375064 148520
rect 375024 56574 375052 148514
rect 375196 145784 375248 145790
rect 375196 145726 375248 145732
rect 375104 144968 375156 144974
rect 375104 144910 375156 144916
rect 375012 56568 375064 56574
rect 375012 56510 375064 56516
rect 375116 55146 375144 144910
rect 375208 144786 375236 145726
rect 375288 145716 375340 145722
rect 375288 145658 375340 145664
rect 375300 144974 375328 145658
rect 375288 144968 375340 144974
rect 375288 144910 375340 144916
rect 375208 144758 375328 144786
rect 375196 144696 375248 144702
rect 375196 144638 375248 144644
rect 375208 59294 375236 144638
rect 375196 59288 375248 59294
rect 375196 59230 375248 59236
rect 375104 55140 375156 55146
rect 375104 55082 375156 55088
rect 374920 54936 374972 54942
rect 374920 54878 374972 54884
rect 375300 54670 375328 144758
rect 375760 55214 375788 162862
rect 375852 146198 375880 266319
rect 375944 265198 375972 369310
rect 375932 265192 375984 265198
rect 375932 265134 375984 265140
rect 375944 164218 375972 265134
rect 375932 164212 375984 164218
rect 375932 164154 375984 164160
rect 375930 146296 375986 146305
rect 375930 146231 375986 146240
rect 375840 146192 375892 146198
rect 375840 146134 375892 146140
rect 375944 145761 375972 146231
rect 375930 145752 375986 145761
rect 375930 145687 375986 145696
rect 375944 59566 375972 145687
rect 375932 59560 375984 59566
rect 375932 59502 375984 59508
rect 376036 57390 376064 468454
rect 376392 461780 376444 461786
rect 376392 461722 376444 461728
rect 376208 461644 376260 461650
rect 376208 461586 376260 461592
rect 376116 460352 376168 460358
rect 376116 460294 376168 460300
rect 376128 162489 376156 460294
rect 376220 266898 376248 461586
rect 376300 460284 376352 460290
rect 376300 460226 376352 460232
rect 376208 266892 376260 266898
rect 376208 266834 376260 266840
rect 376206 265160 376262 265169
rect 376206 265095 376262 265104
rect 376114 162480 376170 162489
rect 376114 162415 376170 162424
rect 376220 161474 376248 265095
rect 376312 161809 376340 460226
rect 376404 267578 376432 461722
rect 376496 373930 376524 475594
rect 376760 470280 376812 470286
rect 376760 470222 376812 470228
rect 376668 467696 376720 467702
rect 376668 467638 376720 467644
rect 376576 465996 376628 466002
rect 376576 465938 376628 465944
rect 376484 373924 376536 373930
rect 376484 373866 376536 373872
rect 376484 371952 376536 371958
rect 376484 371894 376536 371900
rect 376496 371482 376524 371894
rect 376588 371618 376616 465938
rect 376576 371612 376628 371618
rect 376576 371554 376628 371560
rect 376484 371476 376536 371482
rect 376484 371418 376536 371424
rect 376392 267572 376444 267578
rect 376392 267514 376444 267520
rect 376496 266218 376524 371418
rect 376576 371204 376628 371210
rect 376576 371146 376628 371152
rect 376588 370394 376616 371146
rect 376680 370462 376708 467638
rect 376772 405686 376800 470222
rect 376852 464500 376904 464506
rect 376852 464442 376904 464448
rect 376864 407862 376892 464442
rect 377036 411936 377088 411942
rect 377034 411904 377036 411913
rect 377088 411904 377090 411913
rect 377034 411839 377090 411848
rect 376852 407856 376904 407862
rect 376852 407798 376904 407804
rect 376760 405680 376812 405686
rect 376760 405622 376812 405628
rect 376944 385008 376996 385014
rect 376942 384976 376944 384985
rect 376996 384976 376998 384985
rect 376942 384911 376998 384920
rect 376944 383648 376996 383654
rect 376944 383590 376996 383596
rect 376852 383580 376904 383586
rect 376852 383522 376904 383528
rect 376864 383081 376892 383522
rect 376956 383353 376984 383590
rect 376942 383344 376998 383353
rect 376942 383279 376998 383288
rect 376850 383072 376906 383081
rect 376850 383007 376906 383016
rect 376760 373244 376812 373250
rect 376760 373186 376812 373192
rect 376772 372706 376800 373186
rect 376760 372700 376812 372706
rect 376760 372642 376812 372648
rect 376760 372088 376812 372094
rect 376760 372030 376812 372036
rect 376772 371414 376800 372030
rect 376760 371408 376812 371414
rect 376760 371350 376812 371356
rect 376760 371204 376812 371210
rect 376760 371146 376812 371152
rect 376772 370666 376800 371146
rect 376760 370660 376812 370666
rect 376760 370602 376812 370608
rect 376668 370456 376720 370462
rect 376668 370398 376720 370404
rect 376576 370388 376628 370394
rect 376576 370330 376628 370336
rect 376588 267209 376616 370330
rect 376944 369844 376996 369850
rect 376944 369786 376996 369792
rect 376668 369096 376720 369102
rect 376668 369038 376720 369044
rect 376574 267200 376630 267209
rect 376574 267135 376630 267144
rect 376588 266393 376616 267135
rect 376574 266384 376630 266393
rect 376574 266319 376630 266328
rect 376484 266212 376536 266218
rect 376484 266154 376536 266160
rect 376680 265826 376708 369038
rect 376956 368529 376984 369786
rect 376942 368520 376998 368529
rect 376942 368455 376998 368464
rect 377048 306921 377076 411839
rect 377218 410952 377274 410961
rect 377218 410887 377274 410896
rect 377232 410582 377260 410887
rect 377220 410576 377272 410582
rect 377220 410518 377272 410524
rect 377220 409148 377272 409154
rect 377220 409090 377272 409096
rect 377232 408785 377260 409090
rect 377218 408776 377274 408785
rect 377218 408711 377274 408720
rect 377126 407824 377182 407833
rect 377126 407759 377128 407768
rect 377180 407759 377182 407768
rect 377128 407730 377180 407736
rect 377220 406428 377272 406434
rect 377220 406370 377272 406376
rect 377232 406065 377260 406370
rect 377218 406056 377274 406065
rect 377218 405991 377274 406000
rect 377128 369300 377180 369306
rect 377128 369242 377180 369248
rect 377034 306912 377090 306921
rect 377034 306847 377090 306856
rect 377048 306374 377076 306847
rect 376956 306346 377076 306374
rect 376760 278724 376812 278730
rect 376760 278666 376812 278672
rect 376772 278089 376800 278666
rect 376850 278352 376906 278361
rect 376850 278287 376906 278296
rect 376758 278080 376814 278089
rect 376864 278050 376892 278287
rect 376758 278015 376814 278024
rect 376852 278044 376904 278050
rect 376852 277986 376904 277992
rect 376404 265798 376708 265826
rect 376404 265334 376432 265798
rect 376576 265736 376628 265742
rect 376576 265678 376628 265684
rect 376588 265470 376616 265678
rect 376576 265464 376628 265470
rect 376576 265406 376628 265412
rect 376392 265328 376444 265334
rect 376392 265270 376444 265276
rect 376298 161800 376354 161809
rect 376298 161735 376354 161744
rect 376220 161446 376340 161474
rect 376312 160070 376340 161446
rect 376300 160064 376352 160070
rect 376300 160006 376352 160012
rect 376208 146260 376260 146266
rect 376208 146202 376260 146208
rect 376116 145444 376168 145450
rect 376116 145386 376168 145392
rect 376128 58614 376156 145386
rect 376116 58608 376168 58614
rect 376116 58550 376168 58556
rect 376024 57384 376076 57390
rect 376024 57326 376076 57332
rect 376220 56030 376248 146202
rect 376312 59090 376340 160006
rect 376404 159458 376432 265270
rect 376484 263628 376536 263634
rect 376484 263570 376536 263576
rect 376392 159452 376444 159458
rect 376392 159394 376444 159400
rect 376392 148368 376444 148374
rect 376392 148310 376444 148316
rect 376404 147694 376432 148310
rect 376392 147688 376444 147694
rect 376392 147630 376444 147636
rect 376300 59084 376352 59090
rect 376300 59026 376352 59032
rect 376404 56370 376432 147630
rect 376496 145994 376524 263570
rect 376484 145988 376536 145994
rect 376484 145930 376536 145936
rect 376392 56364 376444 56370
rect 376392 56306 376444 56312
rect 376208 56024 376260 56030
rect 376208 55966 376260 55972
rect 375748 55208 375800 55214
rect 375748 55150 375800 55156
rect 376496 54738 376524 145930
rect 376588 145858 376616 265406
rect 376852 264988 376904 264994
rect 376852 264930 376904 264936
rect 376864 180794 376892 264930
rect 376956 202881 376984 306346
rect 377034 303648 377090 303657
rect 377034 303583 377090 303592
rect 376942 202872 376998 202881
rect 376942 202807 376998 202816
rect 377048 200114 377076 303583
rect 377140 265033 377168 369242
rect 377232 301073 377260 405991
rect 377324 373658 377352 477294
rect 377956 477080 378008 477086
rect 377956 477022 378008 477028
rect 377680 471640 377732 471646
rect 377680 471582 377732 471588
rect 377494 407824 377550 407833
rect 377494 407759 377550 407768
rect 377404 388748 377456 388754
rect 377404 388690 377456 388696
rect 377416 374678 377444 388690
rect 377404 374672 377456 374678
rect 377404 374614 377456 374620
rect 377312 373652 377364 373658
rect 377312 373594 377364 373600
rect 377310 305008 377366 305017
rect 377310 304943 377366 304952
rect 377218 301064 377274 301073
rect 377218 300999 377274 301008
rect 377126 265024 377182 265033
rect 377126 264959 377182 264968
rect 376956 200086 377076 200114
rect 376956 198801 376984 200086
rect 376942 198792 376998 198801
rect 376942 198727 376998 198736
rect 376772 180766 376892 180794
rect 376772 171134 376800 180766
rect 376852 175228 376904 175234
rect 376852 175170 376904 175176
rect 376864 175001 376892 175170
rect 376850 174992 376906 175001
rect 376850 174927 376906 174936
rect 376850 173360 376906 173369
rect 376850 173295 376906 173304
rect 376864 173194 376892 173295
rect 376852 173188 376904 173194
rect 376852 173130 376904 173136
rect 376772 171106 376892 171134
rect 376668 158772 376720 158778
rect 376668 158714 376720 158720
rect 376576 145852 376628 145858
rect 376576 145794 376628 145800
rect 376588 145450 376616 145794
rect 376576 145444 376628 145450
rect 376576 145386 376628 145392
rect 376680 59158 376708 158714
rect 376864 146266 376892 171106
rect 376852 146260 376904 146266
rect 376852 146202 376904 146208
rect 376864 146062 376892 146202
rect 376852 146056 376904 146062
rect 376852 145998 376904 146004
rect 376956 93809 376984 198727
rect 377232 196081 377260 300999
rect 377324 200977 377352 304943
rect 377508 302841 377536 407759
rect 377692 405686 377720 471582
rect 377770 410952 377826 410961
rect 377770 410887 377826 410896
rect 377680 405680 377732 405686
rect 377680 405622 377732 405628
rect 377588 405000 377640 405006
rect 377586 404968 377588 404977
rect 377640 404968 377642 404977
rect 377586 404903 377642 404912
rect 377494 302832 377550 302841
rect 377494 302767 377550 302776
rect 377310 200968 377366 200977
rect 377310 200903 377366 200912
rect 377034 196072 377090 196081
rect 377034 196007 377090 196016
rect 377218 196072 377274 196081
rect 377218 196007 377274 196016
rect 376942 93800 376998 93809
rect 376942 93735 376998 93744
rect 377048 91089 377076 196007
rect 377218 193216 377274 193225
rect 377218 193151 377274 193160
rect 377128 173868 377180 173874
rect 377128 173810 377180 173816
rect 377140 173097 377168 173810
rect 377126 173088 377182 173097
rect 377126 173023 377182 173032
rect 377034 91080 377090 91089
rect 377034 91015 377090 91024
rect 377232 88233 377260 193151
rect 377324 95985 377352 200903
rect 377508 197849 377536 302767
rect 377600 299985 377628 404903
rect 377680 403640 377732 403646
rect 377680 403582 377732 403588
rect 377692 403209 377720 403582
rect 377678 403200 377734 403209
rect 377678 403135 377734 403144
rect 377692 300370 377720 403135
rect 377784 388754 377812 410887
rect 377862 408776 377918 408785
rect 377862 408711 377918 408720
rect 377772 388748 377824 388754
rect 377772 388690 377824 388696
rect 377876 388634 377904 408711
rect 377784 388606 377904 388634
rect 377784 379514 377812 388606
rect 377968 388498 377996 477022
rect 378152 476814 378180 520118
rect 383672 518430 383700 520118
rect 387904 518498 387932 520118
rect 387892 518492 387944 518498
rect 387892 518434 387944 518440
rect 383660 518424 383712 518430
rect 383660 518366 383712 518372
rect 391952 485081 391980 520118
rect 396920 519110 396948 520118
rect 396908 519104 396960 519110
rect 396908 519046 396960 519052
rect 401612 518634 401640 520118
rect 401600 518628 401652 518634
rect 401600 518570 401652 518576
rect 406028 518566 406056 520118
rect 406016 518560 406068 518566
rect 406016 518502 406068 518508
rect 410536 518022 410564 520118
rect 414952 519042 414980 520118
rect 414940 519036 414992 519042
rect 414940 518978 414992 518984
rect 419552 518090 419580 520118
rect 423968 518702 423996 520118
rect 423956 518696 424008 518702
rect 423956 518638 424008 518644
rect 419540 518084 419592 518090
rect 419540 518026 419592 518032
rect 410524 518016 410576 518022
rect 410524 517958 410576 517964
rect 427832 514690 427860 520231
rect 428384 514758 428412 558175
rect 429212 518974 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 429384 636880 429436 636886
rect 429384 636822 429436 636828
rect 429290 583332 429346 583341
rect 429290 583267 429346 583276
rect 429200 518968 429252 518974
rect 429200 518910 429252 518916
rect 428372 514752 428424 514758
rect 428372 514694 428424 514700
rect 427820 514684 427872 514690
rect 427820 514626 427872 514632
rect 391938 485072 391994 485081
rect 391938 485007 391994 485016
rect 378140 476808 378192 476814
rect 378140 476750 378192 476756
rect 379152 475856 379204 475862
rect 379152 475798 379204 475804
rect 378784 472728 378836 472734
rect 378784 472670 378836 472676
rect 378048 471708 378100 471714
rect 378048 471650 378100 471656
rect 377876 388470 377996 388498
rect 377876 383654 377904 388470
rect 377876 383626 377996 383654
rect 377784 379486 377904 379514
rect 377772 374672 377824 374678
rect 377772 374614 377824 374620
rect 377784 305969 377812 374614
rect 377770 305960 377826 305969
rect 377770 305895 377826 305904
rect 377784 305017 377812 305895
rect 377770 305008 377826 305017
rect 377770 304943 377826 304952
rect 377876 303657 377904 379486
rect 377968 373998 377996 383626
rect 378060 374406 378088 471650
rect 378600 405680 378652 405686
rect 378600 405622 378652 405628
rect 378048 374400 378100 374406
rect 378048 374342 378100 374348
rect 377956 373992 378008 373998
rect 377956 373934 378008 373940
rect 378048 372700 378100 372706
rect 378048 372642 378100 372648
rect 377956 371408 378008 371414
rect 377956 371350 378008 371356
rect 377862 303648 377918 303657
rect 377862 303583 377918 303592
rect 377692 300342 377904 300370
rect 377586 299976 377642 299985
rect 377586 299911 377642 299920
rect 377770 299976 377826 299985
rect 377770 299911 377826 299920
rect 377678 265024 377734 265033
rect 377678 264959 377734 264968
rect 377586 202872 377642 202881
rect 377586 202807 377642 202816
rect 377600 201929 377628 202807
rect 377586 201920 377642 201929
rect 377586 201855 377642 201864
rect 377494 197840 377550 197849
rect 377494 197775 377550 197784
rect 377310 95976 377366 95985
rect 377310 95911 377366 95920
rect 377508 92857 377536 197775
rect 377600 96937 377628 201855
rect 377692 160002 377720 264959
rect 377784 194993 377812 299911
rect 377876 298217 377904 300342
rect 377862 298208 377918 298217
rect 377862 298143 377918 298152
rect 377770 194984 377826 194993
rect 377770 194919 377826 194928
rect 377680 159996 377732 160002
rect 377680 159938 377732 159944
rect 377692 158778 377720 159938
rect 377680 158772 377732 158778
rect 377680 158714 377732 158720
rect 377680 148300 377732 148306
rect 377680 148242 377732 148248
rect 377586 96928 377642 96937
rect 377586 96863 377642 96872
rect 377494 92848 377550 92857
rect 377494 92783 377550 92792
rect 377218 88224 377274 88233
rect 377218 88159 377274 88168
rect 376944 70372 376996 70378
rect 376944 70314 376996 70320
rect 376956 70009 376984 70314
rect 376942 70000 376998 70009
rect 376942 69935 376998 69944
rect 376942 68368 376998 68377
rect 376942 68303 376944 68312
rect 376996 68303 376998 68312
rect 376944 68274 376996 68280
rect 377692 59498 377720 148242
rect 377784 90001 377812 194919
rect 377876 193225 377904 298143
rect 377968 265606 377996 371350
rect 378060 370002 378088 372642
rect 378060 369974 378180 370002
rect 378048 369844 378100 369850
rect 378048 369786 378100 369792
rect 378060 369510 378088 369786
rect 378048 369504 378100 369510
rect 378048 369446 378100 369452
rect 378152 369322 378180 369974
rect 378612 369578 378640 405622
rect 378600 369572 378652 369578
rect 378600 369514 378652 369520
rect 378060 369294 378180 369322
rect 378060 266150 378088 369294
rect 378692 369028 378744 369034
rect 378692 368970 378744 368976
rect 378600 353388 378652 353394
rect 378600 353330 378652 353336
rect 378612 270502 378640 353330
rect 378600 270496 378652 270502
rect 378600 270438 378652 270444
rect 378048 266144 378100 266150
rect 378048 266086 378100 266092
rect 377956 265600 378008 265606
rect 377956 265542 378008 265548
rect 377862 193216 377918 193225
rect 377862 193151 377918 193160
rect 377968 146266 377996 265542
rect 378060 264994 378088 266086
rect 378508 265056 378560 265062
rect 378508 264998 378560 265004
rect 378048 264988 378100 264994
rect 378048 264930 378100 264936
rect 377956 146260 378008 146266
rect 377956 146202 378008 146208
rect 377770 89992 377826 90001
rect 377770 89927 377826 89936
rect 377680 59492 377732 59498
rect 377680 59434 377732 59440
rect 376668 59152 376720 59158
rect 376668 59094 376720 59100
rect 377968 54874 377996 146202
rect 378520 145790 378548 264998
rect 378600 264988 378652 264994
rect 378600 264930 378652 264936
rect 378612 146130 378640 264930
rect 378704 264790 378732 368970
rect 378692 264784 378744 264790
rect 378692 264726 378744 264732
rect 378704 263634 378732 264726
rect 378692 263628 378744 263634
rect 378692 263570 378744 263576
rect 378796 161974 378824 472670
rect 378876 471368 378928 471374
rect 378876 471310 378928 471316
rect 378888 162353 378916 471310
rect 378968 467356 379020 467362
rect 378968 467298 379020 467304
rect 378980 267617 379008 467298
rect 379060 458856 379112 458862
rect 379060 458798 379112 458804
rect 378966 267608 379022 267617
rect 378966 267543 379022 267552
rect 378968 262880 379020 262886
rect 378968 262822 379020 262828
rect 378980 262206 379008 262822
rect 378968 262200 379020 262206
rect 378968 262142 379020 262148
rect 378874 162344 378930 162353
rect 378874 162279 378930 162288
rect 378784 161968 378836 161974
rect 378784 161910 378836 161916
rect 378980 147422 379008 262142
rect 379072 162625 379100 458798
rect 379164 372638 379192 475798
rect 429304 475425 429332 583267
rect 429396 530913 429424 636822
rect 430948 635520 431000 635526
rect 430948 635462 431000 635468
rect 430580 634908 430632 634914
rect 430580 634850 430632 634856
rect 429844 631100 429896 631106
rect 429844 631042 429896 631048
rect 429856 620974 429884 631042
rect 429844 620968 429896 620974
rect 429844 620910 429896 620916
rect 430592 607209 430620 634850
rect 430856 634840 430908 634846
rect 430856 634782 430908 634788
rect 430762 633448 430818 633457
rect 430762 633383 430818 633392
rect 430670 632224 430726 632233
rect 430670 632159 430726 632168
rect 430684 612513 430712 632159
rect 430776 616865 430804 633383
rect 430868 622033 430896 634782
rect 430960 626521 430988 635462
rect 494072 634098 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 543476 700330 543504 703520
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 494060 634092 494112 634098
rect 494060 634034 494112 634040
rect 435364 633684 435416 633690
rect 435364 633626 435416 633632
rect 432604 633616 432656 633622
rect 432604 633558 432656 633564
rect 430946 626512 431002 626521
rect 430946 626447 431002 626456
rect 430854 622024 430910 622033
rect 430854 621959 430910 621968
rect 432616 621790 432644 633558
rect 432696 631236 432748 631242
rect 432696 631178 432748 631184
rect 432604 621784 432656 621790
rect 432604 621726 432656 621732
rect 432708 621722 432736 631178
rect 432696 621716 432748 621722
rect 432696 621658 432748 621664
rect 430762 616856 430818 616865
rect 430762 616791 430818 616800
rect 430670 612504 430726 612513
rect 430670 612439 430726 612448
rect 435376 608598 435404 633626
rect 494336 633548 494388 633554
rect 494336 633490 494388 633496
rect 457444 632120 457496 632126
rect 457444 632062 457496 632068
rect 456800 620968 456852 620974
rect 456800 620910 456852 620916
rect 456812 619721 456840 620910
rect 456798 619712 456854 619721
rect 456798 619647 456854 619656
rect 435364 608592 435416 608598
rect 435364 608534 435416 608540
rect 456800 608592 456852 608598
rect 456800 608534 456852 608540
rect 456812 607481 456840 608534
rect 456798 607472 456854 607481
rect 456798 607407 456854 607416
rect 430578 607200 430634 607209
rect 430578 607135 430634 607144
rect 430578 588024 430634 588033
rect 430578 587959 430634 587968
rect 429474 553480 429530 553489
rect 429474 553415 429530 553424
rect 429382 530904 429438 530913
rect 429382 530839 429438 530848
rect 429488 515710 429516 553415
rect 430592 517206 430620 587959
rect 457456 582321 457484 632062
rect 457536 631168 457588 631174
rect 457536 631110 457588 631116
rect 457548 613601 457576 631110
rect 471152 631032 471204 631038
rect 471152 630974 471204 630980
rect 465172 621036 465224 621042
rect 465172 620978 465224 620984
rect 465184 619956 465212 620978
rect 471164 619970 471192 630974
rect 483204 621784 483256 621790
rect 483204 621726 483256 621732
rect 477130 619984 477186 619993
rect 471164 619942 471638 619970
rect 477186 619942 477434 619970
rect 483216 619956 483244 621726
rect 488722 619984 488778 619993
rect 477130 619919 477186 619928
rect 494348 619970 494376 633490
rect 510712 633480 510764 633486
rect 510712 633422 510764 633428
rect 510620 630964 510672 630970
rect 510620 630906 510672 630912
rect 501236 621716 501288 621722
rect 501236 621658 501288 621664
rect 488778 619942 489026 619970
rect 494348 619942 494822 619970
rect 501248 619956 501276 621658
rect 506754 619984 506810 619993
rect 488722 619919 488778 619928
rect 506810 619942 507058 619970
rect 506754 619919 506810 619928
rect 457534 613592 457590 613601
rect 457534 613527 457590 613536
rect 510632 604081 510660 630906
rect 510724 617001 510752 633422
rect 512000 630896 512052 630902
rect 512000 630838 512052 630844
rect 580170 630864 580226 630873
rect 510710 616992 510766 617001
rect 510710 616927 510766 616936
rect 512012 610881 512040 630838
rect 580170 630799 580172 630808
rect 580224 630799 580226 630808
rect 580172 630770 580224 630776
rect 515404 621036 515456 621042
rect 515404 620978 515456 620984
rect 511998 610872 512054 610881
rect 511998 610807 512054 610816
rect 510618 604072 510674 604081
rect 510618 604007 510674 604016
rect 457626 601352 457682 601361
rect 457626 601287 457682 601296
rect 457534 588432 457590 588441
rect 457534 588367 457590 588376
rect 457442 582312 457498 582321
rect 457442 582247 457498 582256
rect 430670 578368 430726 578377
rect 430670 578303 430726 578312
rect 430684 525026 430712 578303
rect 457442 576192 457498 576201
rect 457442 576127 457498 576136
rect 430762 572792 430818 572801
rect 430762 572727 430818 572736
rect 430672 525020 430724 525026
rect 430672 524962 430724 524968
rect 430670 524920 430726 524929
rect 430670 524855 430726 524864
rect 430684 519994 430712 524855
rect 430672 519988 430724 519994
rect 430672 519930 430724 519936
rect 430580 517200 430632 517206
rect 430580 517142 430632 517148
rect 430776 517070 430804 572727
rect 430854 567760 430910 567769
rect 430854 567695 430910 567704
rect 430868 520130 430896 567695
rect 430946 563136 431002 563145
rect 430946 563071 431002 563080
rect 430960 525162 430988 563071
rect 431038 549400 431094 549409
rect 431038 549335 431094 549344
rect 430948 525156 431000 525162
rect 430948 525098 431000 525104
rect 430948 525020 431000 525026
rect 430948 524962 431000 524968
rect 430856 520124 430908 520130
rect 430856 520066 430908 520072
rect 430960 519858 430988 524962
rect 430948 519852 431000 519858
rect 430948 519794 431000 519800
rect 431052 517138 431080 549335
rect 431130 543960 431186 543969
rect 431130 543895 431186 543904
rect 431144 518158 431172 543895
rect 431222 539608 431278 539617
rect 431222 539543 431278 539552
rect 431236 525298 431264 539543
rect 431314 534440 431370 534449
rect 431314 534375 431370 534384
rect 431224 525292 431276 525298
rect 431224 525234 431276 525240
rect 431224 525156 431276 525162
rect 431224 525098 431276 525104
rect 431236 519926 431264 525098
rect 431328 520062 431356 534375
rect 431408 525292 431460 525298
rect 431408 525234 431460 525240
rect 431316 520056 431368 520062
rect 431316 519998 431368 520004
rect 431224 519920 431276 519926
rect 431224 519862 431276 519868
rect 431420 519790 431448 525234
rect 457456 520198 457484 576127
rect 457444 520192 457496 520198
rect 457444 520134 457496 520140
rect 431408 519784 431460 519790
rect 431408 519726 431460 519732
rect 431132 518152 431184 518158
rect 431132 518094 431184 518100
rect 431040 517132 431092 517138
rect 431040 517074 431092 517080
rect 430764 517064 430816 517070
rect 430764 517006 430816 517012
rect 429476 515704 429528 515710
rect 429476 515646 429528 515652
rect 457548 479641 457576 588367
rect 457640 515778 457668 601287
rect 511998 597952 512054 597961
rect 511998 597887 512054 597896
rect 457718 594552 457774 594561
rect 457718 594487 457774 594496
rect 457732 517274 457760 594487
rect 459572 570030 460046 570058
rect 465092 570030 465842 570058
rect 470612 570030 471638 570058
rect 476132 570030 477434 570058
rect 483032 570030 483230 570058
rect 488552 570030 489670 570058
rect 459572 517342 459600 570030
rect 459560 517336 459612 517342
rect 459560 517278 459612 517284
rect 457720 517268 457772 517274
rect 457720 517210 457772 517216
rect 465092 515846 465120 570030
rect 470612 515914 470640 570030
rect 476132 520266 476160 570030
rect 476120 520260 476172 520266
rect 476120 520202 476172 520208
rect 470600 515908 470652 515914
rect 470600 515850 470652 515856
rect 465080 515840 465132 515846
rect 465080 515782 465132 515788
rect 457628 515772 457680 515778
rect 457628 515714 457680 515720
rect 483032 482225 483060 570030
rect 488552 515982 488580 570030
rect 495452 517410 495480 570044
rect 500972 570030 501262 570058
rect 506492 570030 507058 570058
rect 495440 517404 495492 517410
rect 495440 517346 495492 517352
rect 500972 516050 501000 570030
rect 500960 516044 501012 516050
rect 500960 515986 501012 515992
rect 488540 515976 488592 515982
rect 488540 515918 488592 515924
rect 483018 482216 483074 482225
rect 483018 482151 483074 482160
rect 506492 479777 506520 570030
rect 506478 479768 506534 479777
rect 506478 479703 506534 479712
rect 457534 479632 457590 479641
rect 457534 479567 457590 479576
rect 512012 478417 512040 597887
rect 512182 591832 512238 591841
rect 512182 591767 512238 591776
rect 512090 585712 512146 585721
rect 512090 585647 512146 585656
rect 511998 478408 512054 478417
rect 511998 478343 512054 478352
rect 429290 475416 429346 475425
rect 429290 475351 429346 475360
rect 379980 474428 380032 474434
rect 379980 474370 380032 474376
rect 379244 467628 379296 467634
rect 379244 467570 379296 467576
rect 379152 372632 379204 372638
rect 379152 372574 379204 372580
rect 379256 370666 379284 467570
rect 379336 464364 379388 464370
rect 379336 464306 379388 464312
rect 379348 383654 379376 464306
rect 379348 383626 379468 383654
rect 379336 372632 379388 372638
rect 379336 372574 379388 372580
rect 379244 370660 379296 370666
rect 379244 370602 379296 370608
rect 379256 354674 379284 370602
rect 379348 369854 379376 372574
rect 379440 371958 379468 383626
rect 379992 372026 380020 474370
rect 512104 474065 512132 585647
rect 512196 516118 512224 591767
rect 515416 585818 515444 620978
rect 515404 585812 515456 585818
rect 515404 585754 515456 585760
rect 580172 585812 580224 585818
rect 580172 585754 580224 585760
rect 512274 579592 512330 579601
rect 512274 579527 512330 579536
rect 512288 517478 512316 579527
rect 580184 577697 580212 585754
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 513286 572792 513342 572801
rect 513286 572727 513288 572736
rect 513340 572727 513342 572736
rect 560944 572756 560996 572762
rect 513288 572698 513340 572704
rect 560944 572698 560996 572704
rect 512276 517472 512328 517478
rect 512276 517414 512328 517420
rect 519544 516180 519596 516186
rect 519544 516122 519596 516128
rect 512184 516112 512236 516118
rect 512184 516054 512236 516060
rect 512090 474056 512146 474065
rect 512090 473991 512146 474000
rect 498200 461168 498252 461174
rect 498200 461110 498252 461116
rect 517704 461168 517756 461174
rect 517704 461110 517756 461116
rect 498212 461009 498240 461110
rect 499856 461032 499908 461038
rect 498198 461000 498254 461009
rect 498198 460935 498200 460944
rect 498252 460935 498254 460944
rect 499854 461000 499856 461009
rect 517612 461032 517664 461038
rect 499908 461000 499910 461009
rect 499854 460935 499910 460944
rect 510894 461000 510950 461009
rect 517612 460974 517664 460980
rect 510894 460935 510896 460944
rect 498200 460906 498252 460912
rect 510948 460935 510950 460944
rect 517520 460964 517572 460970
rect 510896 460906 510948 460912
rect 517520 460906 517572 460912
rect 516600 458312 516652 458318
rect 516600 458254 516652 458260
rect 516612 454753 516640 458254
rect 516598 454744 516654 454753
rect 516598 454679 516654 454688
rect 407762 375048 407818 375057
rect 380900 375012 380952 375018
rect 407762 374983 407818 374992
rect 425058 375048 425114 375057
rect 425058 374983 425114 374992
rect 440330 375048 440386 375057
rect 440330 374983 440386 374992
rect 443090 375048 443146 375057
rect 443090 374983 443146 374992
rect 380900 374954 380952 374960
rect 380912 374474 380940 374954
rect 404174 374776 404230 374785
rect 404174 374711 404230 374720
rect 404188 374678 404216 374711
rect 404176 374672 404228 374678
rect 404176 374614 404228 374620
rect 407776 374610 407804 374983
rect 410706 374640 410762 374649
rect 407764 374604 407816 374610
rect 410706 374575 410762 374584
rect 407764 374546 407816 374552
rect 410720 374542 410748 374575
rect 410708 374536 410760 374542
rect 410708 374478 410760 374484
rect 425072 374474 425100 374983
rect 433614 374504 433670 374513
rect 380900 374468 380952 374474
rect 380900 374410 380952 374416
rect 425060 374468 425112 374474
rect 433614 374439 433670 374448
rect 436006 374504 436062 374513
rect 436006 374439 436062 374448
rect 438490 374504 438546 374513
rect 438490 374439 438546 374448
rect 425060 374410 425112 374416
rect 379520 372020 379572 372026
rect 379520 371962 379572 371968
rect 379980 372020 380032 372026
rect 379980 371962 380032 371968
rect 379428 371952 379480 371958
rect 379428 371894 379480 371900
rect 379440 371362 379468 371894
rect 379532 371686 379560 371962
rect 379520 371680 379572 371686
rect 379520 371622 379572 371628
rect 379888 371680 379940 371686
rect 379888 371622 379940 371628
rect 379440 371334 379560 371362
rect 379348 369826 379468 369854
rect 379336 368144 379388 368150
rect 379336 368086 379388 368092
rect 379164 354646 379284 354674
rect 379164 251122 379192 354646
rect 379244 353320 379296 353326
rect 379244 353262 379296 353268
rect 379256 266286 379284 353262
rect 379244 266280 379296 266286
rect 379244 266222 379296 266228
rect 379152 251116 379204 251122
rect 379152 251058 379204 251064
rect 379058 162616 379114 162625
rect 379058 162551 379114 162560
rect 378968 147416 379020 147422
rect 378968 147358 379020 147364
rect 379150 146296 379206 146305
rect 379150 146231 379206 146240
rect 379060 146192 379112 146198
rect 379060 146134 379112 146140
rect 378600 146124 378652 146130
rect 378600 146066 378652 146072
rect 378508 145784 378560 145790
rect 378508 145726 378560 145732
rect 378612 145654 378640 146066
rect 378048 145648 378100 145654
rect 378048 145590 378100 145596
rect 378600 145648 378652 145654
rect 378600 145590 378652 145596
rect 378784 145648 378836 145654
rect 378784 145590 378836 145596
rect 377956 54868 378008 54874
rect 377956 54810 378008 54816
rect 378060 54806 378088 145590
rect 378796 144906 378824 145590
rect 378876 145512 378928 145518
rect 378876 145454 378928 145460
rect 378784 144900 378836 144906
rect 378784 144842 378836 144848
rect 378048 54800 378100 54806
rect 378048 54742 378100 54748
rect 376484 54732 376536 54738
rect 376484 54674 376536 54680
rect 375288 54664 375340 54670
rect 375288 54606 375340 54612
rect 378796 54602 378824 144842
rect 378888 144838 378916 145454
rect 379072 145450 379100 146134
rect 379164 145897 379192 146231
rect 379256 146198 379284 266222
rect 379348 264246 379376 368086
rect 379440 265713 379468 369826
rect 379532 364334 379560 371334
rect 379796 370456 379848 370462
rect 379796 370398 379848 370404
rect 379532 364306 379744 364334
rect 379612 270496 379664 270502
rect 379612 270438 379664 270444
rect 379624 269550 379652 270438
rect 379612 269544 379664 269550
rect 379612 269486 379664 269492
rect 379520 269068 379572 269074
rect 379520 269010 379572 269016
rect 379532 267918 379560 269010
rect 379520 267912 379572 267918
rect 379520 267854 379572 267860
rect 379426 265704 379482 265713
rect 379426 265639 379482 265648
rect 379440 265033 379468 265639
rect 379426 265024 379482 265033
rect 379426 264959 379482 264968
rect 379336 264240 379388 264246
rect 379336 264182 379388 264188
rect 379348 263634 379376 264182
rect 379336 263628 379388 263634
rect 379336 263570 379388 263576
rect 379428 251116 379480 251122
rect 379428 251058 379480 251064
rect 379440 251025 379468 251058
rect 379426 251016 379482 251025
rect 379426 250951 379482 250960
rect 379428 147688 379480 147694
rect 379428 147630 379480 147636
rect 379336 147620 379388 147626
rect 379336 147562 379388 147568
rect 379348 147422 379376 147562
rect 379336 147416 379388 147422
rect 379336 147358 379388 147364
rect 379244 146192 379296 146198
rect 379244 146134 379296 146140
rect 379150 145888 379206 145897
rect 379150 145823 379206 145832
rect 379060 145444 379112 145450
rect 379060 145386 379112 145392
rect 378968 145376 379020 145382
rect 378968 145318 379020 145324
rect 378876 144832 378928 144838
rect 378876 144774 378928 144780
rect 378888 59702 378916 144774
rect 378876 59696 378928 59702
rect 378876 59638 378928 59644
rect 378980 59634 379008 145318
rect 379072 59770 379100 145386
rect 379060 59764 379112 59770
rect 379060 59706 379112 59712
rect 378968 59628 379020 59634
rect 378968 59570 379020 59576
rect 379164 57254 379192 145823
rect 379152 57248 379204 57254
rect 379152 57190 379204 57196
rect 379256 55962 379284 146134
rect 379348 56302 379376 147358
rect 379336 56296 379388 56302
rect 379336 56238 379388 56244
rect 379440 56098 379468 147630
rect 379532 146305 379560 267854
rect 379624 171134 379652 269486
rect 379716 265878 379744 364306
rect 379808 269074 379836 370398
rect 379796 269068 379848 269074
rect 379796 269010 379848 269016
rect 379900 266082 379928 371622
rect 379992 266354 380020 371962
rect 380912 353394 380940 374410
rect 433628 374134 433656 374439
rect 436020 374338 436048 374439
rect 436008 374332 436060 374338
rect 436008 374274 436060 374280
rect 438504 374270 438532 374439
rect 438492 374264 438544 374270
rect 438492 374206 438544 374212
rect 440344 374202 440372 374983
rect 443104 374406 443132 374983
rect 451002 374640 451058 374649
rect 451002 374575 451058 374584
rect 443092 374400 443144 374406
rect 443092 374342 443144 374348
rect 440332 374196 440384 374202
rect 440332 374138 440384 374144
rect 433616 374128 433668 374134
rect 433616 374070 433668 374076
rect 451016 374066 451044 374575
rect 451004 374060 451056 374066
rect 451004 374002 451056 374008
rect 421012 373992 421064 373998
rect 421012 373934 421064 373940
rect 421024 373833 421052 373934
rect 423036 373924 423088 373930
rect 423036 373866 423088 373872
rect 423048 373833 423076 373866
rect 426900 373856 426952 373862
rect 416042 373824 416098 373833
rect 416042 373759 416044 373768
rect 416096 373759 416098 373768
rect 421010 373824 421066 373833
rect 421010 373759 421066 373768
rect 423034 373824 423090 373833
rect 423034 373759 423090 373768
rect 426898 373824 426900 373833
rect 426952 373824 426954 373833
rect 426898 373759 426954 373768
rect 430578 373824 430634 373833
rect 430578 373759 430634 373768
rect 416044 373730 416096 373736
rect 430592 373726 430620 373759
rect 430580 373720 430632 373726
rect 430580 373662 430632 373668
rect 445850 373688 445906 373697
rect 445850 373623 445906 373632
rect 455418 373688 455474 373697
rect 455418 373623 455420 373632
rect 445864 373590 445892 373623
rect 455472 373623 455474 373632
rect 455420 373594 455472 373600
rect 445852 373584 445904 373590
rect 445852 373526 445904 373532
rect 447690 373552 447746 373561
rect 447690 373487 447692 373496
rect 447744 373487 447746 373496
rect 458178 373552 458234 373561
rect 458178 373487 458234 373496
rect 447692 373458 447744 373464
rect 458192 373454 458220 373487
rect 458180 373448 458232 373454
rect 452842 373416 452898 373425
rect 458180 373390 458232 373396
rect 485778 373416 485834 373425
rect 452842 373351 452844 373360
rect 452896 373351 452898 373360
rect 485778 373351 485834 373360
rect 452844 373322 452896 373328
rect 485792 373318 485820 373351
rect 485780 373312 485832 373318
rect 485780 373254 485832 373260
rect 408500 372700 408552 372706
rect 408500 372642 408552 372648
rect 408512 372609 408540 372642
rect 426440 372632 426492 372638
rect 408498 372600 408554 372609
rect 408498 372535 408554 372544
rect 426438 372600 426440 372609
rect 426492 372600 426494 372609
rect 426438 372535 426494 372544
rect 433338 372600 433394 372609
rect 433338 372535 433394 372544
rect 437478 372600 437534 372609
rect 437478 372535 437480 372544
rect 433352 372502 433380 372535
rect 437532 372535 437534 372544
rect 437480 372506 437532 372512
rect 433340 372496 433392 372502
rect 433340 372438 433392 372444
rect 470598 372328 470654 372337
rect 470598 372263 470654 372272
rect 404358 372192 404414 372201
rect 404358 372127 404414 372136
rect 396078 372056 396134 372065
rect 396078 371991 396080 372000
rect 396132 371991 396134 372000
rect 397458 372056 397514 372065
rect 397458 371991 397514 372000
rect 398838 372056 398894 372065
rect 398838 371991 398894 372000
rect 400218 372056 400274 372065
rect 400218 371991 400274 372000
rect 396080 371962 396132 371968
rect 381082 371920 381138 371929
rect 381082 371855 381138 371864
rect 380992 371612 381044 371618
rect 380992 371554 381044 371560
rect 380900 353388 380952 353394
rect 380900 353330 380952 353336
rect 381004 353326 381032 371554
rect 381096 354006 381124 371855
rect 397472 371754 397500 371991
rect 398852 371822 398880 371991
rect 400232 371890 400260 371991
rect 404372 371958 404400 372127
rect 409878 372056 409934 372065
rect 409878 371991 409934 372000
rect 404360 371952 404412 371958
rect 404360 371894 404412 371900
rect 400220 371884 400272 371890
rect 400220 371826 400272 371832
rect 398840 371816 398892 371822
rect 398840 371758 398892 371764
rect 397460 371748 397512 371754
rect 397460 371690 397512 371696
rect 409892 371686 409920 371991
rect 439870 371784 439926 371793
rect 439870 371719 439926 371728
rect 409880 371680 409932 371686
rect 401598 371648 401654 371657
rect 409880 371622 409932 371628
rect 411258 371648 411314 371657
rect 401598 371583 401654 371592
rect 411258 371583 411260 371592
rect 401612 371550 401640 371583
rect 411312 371583 411314 371592
rect 418342 371648 418398 371657
rect 418342 371583 418398 371592
rect 423678 371648 423734 371657
rect 423678 371583 423734 371592
rect 427818 371648 427874 371657
rect 427818 371583 427874 371592
rect 411260 371554 411312 371560
rect 401600 371544 401652 371550
rect 401600 371486 401652 371492
rect 407118 371512 407174 371521
rect 407118 371447 407120 371456
rect 407172 371447 407174 371456
rect 411258 371512 411314 371521
rect 411258 371447 411314 371456
rect 418250 371512 418306 371521
rect 418250 371447 418306 371456
rect 407120 371418 407172 371424
rect 411272 371414 411300 371447
rect 411260 371408 411312 371414
rect 396078 371376 396134 371385
rect 396078 371311 396134 371320
rect 402978 371376 403034 371385
rect 402978 371311 403034 371320
rect 405738 371376 405794 371385
rect 411260 371350 411312 371356
rect 412638 371376 412694 371385
rect 405738 371311 405794 371320
rect 412638 371311 412694 371320
rect 413190 371376 413246 371385
rect 413190 371311 413246 371320
rect 414018 371376 414074 371385
rect 414018 371311 414074 371320
rect 415398 371376 415454 371385
rect 415398 371311 415454 371320
rect 416778 371376 416834 371385
rect 416778 371311 416834 371320
rect 418158 371376 418214 371385
rect 418158 371311 418214 371320
rect 396092 370394 396120 371311
rect 402992 371210 403020 371311
rect 402980 371204 403032 371210
rect 402980 371146 403032 371152
rect 396080 370388 396132 370394
rect 396080 370330 396132 370336
rect 405752 369034 405780 371311
rect 405740 369028 405792 369034
rect 405740 368970 405792 368976
rect 412652 368150 412680 371311
rect 413204 370734 413232 371311
rect 413192 370728 413244 370734
rect 413192 370670 413244 370676
rect 414032 370462 414060 371311
rect 415412 370666 415440 371311
rect 415400 370660 415452 370666
rect 415400 370602 415452 370608
rect 414020 370456 414072 370462
rect 414020 370398 414072 370404
rect 416792 369442 416820 371311
rect 418172 369714 418200 371311
rect 418160 369708 418212 369714
rect 418160 369650 418212 369656
rect 416780 369436 416832 369442
rect 416780 369378 416832 369384
rect 418264 369374 418292 371447
rect 418252 369368 418304 369374
rect 418252 369310 418304 369316
rect 418356 369102 418384 371583
rect 420918 371512 420974 371521
rect 420918 371447 420974 371456
rect 419538 371376 419594 371385
rect 419538 371311 419594 371320
rect 419552 369306 419580 371311
rect 419540 369300 419592 369306
rect 419540 369242 419592 369248
rect 420932 369238 420960 371447
rect 422298 371376 422354 371385
rect 422298 371311 422354 371320
rect 422312 370598 422340 371311
rect 422300 370592 422352 370598
rect 422300 370534 422352 370540
rect 423692 369510 423720 371583
rect 425058 371376 425114 371385
rect 425058 371311 425114 371320
rect 425072 369578 425100 371311
rect 427832 369646 427860 371583
rect 439884 371414 439912 371719
rect 462318 371648 462374 371657
rect 462318 371583 462374 371592
rect 465078 371648 465134 371657
rect 465078 371583 465134 371592
rect 439872 371408 439924 371414
rect 427910 371376 427966 371385
rect 427910 371311 427966 371320
rect 431958 371376 432014 371385
rect 431958 371311 432014 371320
rect 434718 371376 434774 371385
rect 434718 371311 434774 371320
rect 436098 371376 436154 371385
rect 439872 371350 439924 371356
rect 460938 371376 460994 371385
rect 436098 371311 436154 371320
rect 460938 371311 460994 371320
rect 427820 369640 427872 369646
rect 427820 369582 427872 369588
rect 425060 369572 425112 369578
rect 425060 369514 425112 369520
rect 423680 369504 423732 369510
rect 423680 369446 423732 369452
rect 420920 369232 420972 369238
rect 420920 369174 420972 369180
rect 418344 369096 418396 369102
rect 418344 369038 418396 369044
rect 412640 368144 412692 368150
rect 412640 368086 412692 368092
rect 427924 368082 427952 371311
rect 427912 368076 427964 368082
rect 427912 368018 427964 368024
rect 431972 367946 432000 371311
rect 431960 367940 432012 367946
rect 431960 367882 432012 367888
rect 434732 367878 434760 371311
rect 436112 368014 436140 371311
rect 460952 370802 460980 371311
rect 462332 370870 462360 371583
rect 465092 371074 465120 371583
rect 467838 371376 467894 371385
rect 467838 371311 467894 371320
rect 465080 371068 465132 371074
rect 465080 371010 465132 371016
rect 467852 371006 467880 371311
rect 467840 371000 467892 371006
rect 467840 370942 467892 370948
rect 470612 370938 470640 372263
rect 503166 372192 503222 372201
rect 503166 372127 503222 372136
rect 503534 372192 503590 372201
rect 503534 372127 503590 372136
rect 477498 371648 477554 371657
rect 477498 371583 477554 371592
rect 473358 371376 473414 371385
rect 473358 371311 473414 371320
rect 473372 371142 473400 371311
rect 473360 371136 473412 371142
rect 473360 371078 473412 371084
rect 470600 370932 470652 370938
rect 470600 370874 470652 370880
rect 462320 370864 462372 370870
rect 462320 370806 462372 370812
rect 460940 370796 460992 370802
rect 460940 370738 460992 370744
rect 477512 369782 477540 371583
rect 480258 371512 480314 371521
rect 480258 371447 480314 371456
rect 477500 369776 477552 369782
rect 477500 369718 477552 369724
rect 480272 368966 480300 371447
rect 483018 371376 483074 371385
rect 483018 371311 483074 371320
rect 483032 370326 483060 371311
rect 503180 371278 503208 372127
rect 503548 371346 503576 372127
rect 516600 371408 516652 371414
rect 516600 371350 516652 371356
rect 503536 371340 503588 371346
rect 503536 371282 503588 371288
rect 503168 371272 503220 371278
rect 503168 371214 503220 371220
rect 483020 370320 483072 370326
rect 483020 370262 483072 370268
rect 480260 368960 480312 368966
rect 480260 368902 480312 368908
rect 436100 368008 436152 368014
rect 436100 367950 436152 367956
rect 434720 367872 434772 367878
rect 434720 367814 434772 367820
rect 500868 355496 500920 355502
rect 500868 355438 500920 355444
rect 498844 355428 498896 355434
rect 498844 355370 498896 355376
rect 498856 355065 498884 355370
rect 498842 355056 498898 355065
rect 498842 354991 498898 355000
rect 500880 354929 500908 355438
rect 500866 354920 500922 354929
rect 500866 354855 500922 354864
rect 510896 354816 510948 354822
rect 510894 354784 510896 354793
rect 510948 354784 510950 354793
rect 510894 354719 510950 354728
rect 381084 354000 381136 354006
rect 381084 353942 381136 353948
rect 380992 353320 381044 353326
rect 380992 353262 381044 353268
rect 416042 269784 416098 269793
rect 416042 269719 416098 269728
rect 425242 269784 425298 269793
rect 425242 269719 425298 269728
rect 433338 269784 433394 269793
rect 433338 269719 433394 269728
rect 434350 269784 434406 269793
rect 434350 269719 434406 269728
rect 416056 269482 416084 269719
rect 425256 269550 425284 269719
rect 429750 269648 429806 269657
rect 429750 269583 429806 269592
rect 425244 269544 425296 269550
rect 425244 269486 425296 269492
rect 416044 269476 416096 269482
rect 416044 269418 416096 269424
rect 422850 268968 422906 268977
rect 422850 268903 422906 268912
rect 425978 268968 426034 268977
rect 425978 268903 426034 268912
rect 422864 268870 422892 268903
rect 422852 268864 422904 268870
rect 416962 268832 417018 268841
rect 416962 268767 417018 268776
rect 421010 268832 421066 268841
rect 422852 268806 422904 268812
rect 421010 268767 421066 268776
rect 398194 268152 398250 268161
rect 396724 268116 396776 268122
rect 398194 268087 398250 268096
rect 401690 268152 401746 268161
rect 401690 268087 401746 268096
rect 415400 268116 415452 268122
rect 396724 268058 396776 268064
rect 395344 268048 395396 268054
rect 395344 267990 395396 267996
rect 379980 266348 380032 266354
rect 379980 266290 380032 266296
rect 379888 266076 379940 266082
rect 379888 266018 379940 266024
rect 379704 265872 379756 265878
rect 379704 265814 379756 265820
rect 379716 265062 379744 265814
rect 379704 265056 379756 265062
rect 379704 264998 379756 265004
rect 379900 264994 379928 266018
rect 379992 265266 380020 266290
rect 379980 265260 380032 265266
rect 379980 265202 380032 265208
rect 388442 265160 388498 265169
rect 388442 265095 388498 265104
rect 379978 265024 380034 265033
rect 379888 264988 379940 264994
rect 379978 264959 380034 264968
rect 379888 264930 379940 264936
rect 379888 263628 379940 263634
rect 379888 263570 379940 263576
rect 379624 171106 379744 171134
rect 379716 161362 379744 171106
rect 379704 161356 379756 161362
rect 379704 161298 379756 161304
rect 379612 159452 379664 159458
rect 379612 159394 379664 159400
rect 379518 146296 379574 146305
rect 379518 146231 379574 146240
rect 379624 59226 379652 159394
rect 379612 59220 379664 59226
rect 379612 59162 379664 59168
rect 379716 59022 379744 161298
rect 379796 160132 379848 160138
rect 379796 160074 379848 160080
rect 379704 59016 379756 59022
rect 379704 58958 379756 58964
rect 379808 56234 379836 160074
rect 379900 148986 379928 263570
rect 379992 161430 380020 264959
rect 388456 264926 388484 265095
rect 390560 265056 390612 265062
rect 389178 265024 389234 265033
rect 390560 264998 390612 265004
rect 389178 264959 389234 264968
rect 388444 264920 388496 264926
rect 388444 264862 388496 264868
rect 389192 264858 389220 264959
rect 389180 264852 389232 264858
rect 389180 264794 389232 264800
rect 390572 264722 390600 264998
rect 391940 264988 391992 264994
rect 391940 264930 391992 264936
rect 390560 264716 390612 264722
rect 390560 264658 390612 264664
rect 391952 264654 391980 264930
rect 391940 264648 391992 264654
rect 391940 264590 391992 264596
rect 395356 251190 395384 267990
rect 396078 266384 396134 266393
rect 396078 266319 396080 266328
rect 396132 266319 396134 266328
rect 396080 266290 396132 266296
rect 395344 251184 395396 251190
rect 395344 251126 395396 251132
rect 396736 251122 396764 268058
rect 398208 265810 398236 268087
rect 398838 266384 398894 266393
rect 398838 266319 398894 266328
rect 400218 266384 400274 266393
rect 400218 266319 400274 266328
rect 398852 265946 398880 266319
rect 400232 266014 400260 266319
rect 400220 266008 400272 266014
rect 400220 265950 400272 265956
rect 398840 265940 398892 265946
rect 398840 265882 398892 265888
rect 398196 265804 398248 265810
rect 398196 265746 398248 265752
rect 401704 265674 401732 268087
rect 415400 268058 415452 268064
rect 402980 267980 403032 267986
rect 402980 267922 403032 267928
rect 402992 267753 403020 267922
rect 414388 267912 414440 267918
rect 414388 267854 414440 267860
rect 414400 267753 414428 267854
rect 415412 267753 415440 268058
rect 416976 268054 417004 268767
rect 421024 268666 421052 268767
rect 425992 268734 426020 268903
rect 425980 268728 426032 268734
rect 425980 268670 426032 268676
rect 421012 268660 421064 268666
rect 421012 268602 421064 268608
rect 429764 268258 429792 269583
rect 433352 269414 433380 269719
rect 433340 269408 433392 269414
rect 433340 269350 433392 269356
rect 434364 269346 434392 269719
rect 436006 269648 436062 269657
rect 436006 269583 436062 269592
rect 468482 269648 468538 269657
rect 468482 269583 468538 269592
rect 470966 269648 471022 269657
rect 470966 269583 471022 269592
rect 480902 269648 480958 269657
rect 480902 269583 480958 269592
rect 434352 269340 434404 269346
rect 434352 269282 434404 269288
rect 436020 269278 436048 269583
rect 436008 269272 436060 269278
rect 436008 269214 436060 269220
rect 468496 269210 468524 269583
rect 468484 269204 468536 269210
rect 468484 269146 468536 269152
rect 470980 269142 471008 269583
rect 470968 269136 471020 269142
rect 470968 269078 471020 269084
rect 430946 268968 431002 268977
rect 430946 268903 431002 268912
rect 432234 268968 432290 268977
rect 432234 268903 432290 268912
rect 475842 268968 475898 268977
rect 475842 268903 475898 268912
rect 478418 268968 478474 268977
rect 478418 268903 478474 268912
rect 430960 268802 430988 268903
rect 430948 268796 431000 268802
rect 430948 268738 431000 268744
rect 429752 268252 429804 268258
rect 429752 268194 429804 268200
rect 432248 268190 432276 268903
rect 475856 268598 475884 268903
rect 475844 268592 475896 268598
rect 475844 268534 475896 268540
rect 478432 268530 478460 268903
rect 478420 268524 478472 268530
rect 478420 268466 478472 268472
rect 480916 268462 480944 269583
rect 483386 268968 483442 268977
rect 483386 268903 483442 268912
rect 480904 268456 480956 268462
rect 480904 268398 480956 268404
rect 483400 268394 483428 268903
rect 483388 268388 483440 268394
rect 483388 268330 483440 268336
rect 432236 268184 432288 268190
rect 432236 268126 432288 268132
rect 455786 268152 455842 268161
rect 455786 268087 455842 268096
rect 416964 268048 417016 268054
rect 416964 267990 417016 267996
rect 427084 267844 427136 267850
rect 427084 267786 427136 267792
rect 434720 267844 434772 267850
rect 434720 267786 434772 267792
rect 425704 267776 425756 267782
rect 402978 267744 403034 267753
rect 402978 267679 403034 267688
rect 414386 267744 414442 267753
rect 414386 267679 414442 267688
rect 415398 267744 415454 267753
rect 425704 267718 425756 267724
rect 415398 267679 415454 267688
rect 418158 267200 418214 267209
rect 418158 267135 418214 267144
rect 409878 267064 409934 267073
rect 409878 266999 409934 267008
rect 412914 267064 412970 267073
rect 412914 266999 412970 267008
rect 409892 266830 409920 266999
rect 412928 266898 412956 266999
rect 418172 266966 418200 267135
rect 418160 266960 418212 266966
rect 418160 266902 418212 266908
rect 412916 266892 412968 266898
rect 412916 266834 412968 266840
rect 409880 266824 409932 266830
rect 409880 266766 409932 266772
rect 408498 266656 408554 266665
rect 408498 266591 408554 266600
rect 403162 266384 403218 266393
rect 403162 266319 403218 266328
rect 404358 266384 404414 266393
rect 404358 266319 404414 266328
rect 405738 266384 405794 266393
rect 405738 266319 405794 266328
rect 407118 266384 407174 266393
rect 407118 266319 407174 266328
rect 403176 265742 403204 266319
rect 404372 265878 404400 266319
rect 404360 265872 404412 265878
rect 404360 265814 404412 265820
rect 403164 265736 403216 265742
rect 403164 265678 403216 265684
rect 401692 265668 401744 265674
rect 401692 265610 401744 265616
rect 405752 264790 405780 266319
rect 407132 266218 407160 266319
rect 407120 266212 407172 266218
rect 407120 266154 407172 266160
rect 408512 266150 408540 266591
rect 411350 266520 411406 266529
rect 411350 266455 411406 266464
rect 418250 266520 418306 266529
rect 418250 266455 418306 266464
rect 409878 266384 409934 266393
rect 409878 266319 409934 266328
rect 411258 266384 411314 266393
rect 411258 266319 411314 266328
rect 408500 266144 408552 266150
rect 408500 266086 408552 266092
rect 409892 266082 409920 266319
rect 411272 266286 411300 266319
rect 411260 266280 411312 266286
rect 411260 266222 411312 266228
rect 409880 266076 409932 266082
rect 409880 266018 409932 266024
rect 411364 265606 411392 266455
rect 413006 266384 413062 266393
rect 413006 266319 413062 266328
rect 418158 266384 418214 266393
rect 418158 266319 418214 266328
rect 411352 265600 411404 265606
rect 411352 265542 411404 265548
rect 405740 264784 405792 264790
rect 405740 264726 405792 264732
rect 413020 264246 413048 266319
rect 418172 264654 418200 266319
rect 418264 264722 418292 266455
rect 421564 266416 421616 266422
rect 419538 266384 419594 266393
rect 419538 266319 419594 266328
rect 420918 266384 420974 266393
rect 421564 266358 421616 266364
rect 420918 266319 420974 266328
rect 419552 264858 419580 266319
rect 420932 264926 420960 266319
rect 420920 264920 420972 264926
rect 420920 264862 420972 264868
rect 419540 264852 419592 264858
rect 419540 264794 419592 264800
rect 418252 264716 418304 264722
rect 418252 264658 418304 264664
rect 418160 264648 418212 264654
rect 418160 264590 418212 264596
rect 413008 264240 413060 264246
rect 413008 264182 413060 264188
rect 396724 251116 396776 251122
rect 396724 251058 396776 251064
rect 421576 250646 421604 266358
rect 421564 250640 421616 250646
rect 421564 250582 421616 250588
rect 425716 250578 425744 267718
rect 426438 266384 426494 266393
rect 426438 266319 426494 266328
rect 426452 262886 426480 266319
rect 426440 262880 426492 262886
rect 426440 262822 426492 262828
rect 425704 250572 425756 250578
rect 425704 250514 425756 250520
rect 427096 250510 427124 267786
rect 428556 267776 428608 267782
rect 434732 267753 434760 267786
rect 428646 267744 428702 267753
rect 428608 267724 428646 267734
rect 428556 267718 428646 267724
rect 428568 267706 428646 267718
rect 428646 267679 428702 267688
rect 434718 267744 434774 267753
rect 434718 267679 434774 267688
rect 449898 267744 449954 267753
rect 449898 267679 449954 267688
rect 452658 267744 452714 267753
rect 452658 267679 452714 267688
rect 449912 267510 449940 267679
rect 452672 267646 452700 267679
rect 452660 267640 452712 267646
rect 452660 267582 452712 267588
rect 449900 267504 449952 267510
rect 442998 267472 443054 267481
rect 449900 267446 449952 267452
rect 455800 267442 455828 268087
rect 458178 267744 458234 267753
rect 458178 267679 458234 267688
rect 460938 267744 460994 267753
rect 460938 267679 460940 267688
rect 458192 267578 458220 267679
rect 460992 267679 460994 267688
rect 460940 267650 460992 267656
rect 458180 267572 458232 267578
rect 458180 267514 458232 267520
rect 503166 267472 503222 267481
rect 442998 267407 443054 267416
rect 455788 267436 455840 267442
rect 443012 267374 443040 267407
rect 503166 267407 503222 267416
rect 503534 267472 503590 267481
rect 503534 267407 503590 267416
rect 455788 267378 455840 267384
rect 443000 267368 443052 267374
rect 440054 267336 440110 267345
rect 440054 267271 440110 267280
rect 440238 267336 440294 267345
rect 443000 267310 443052 267316
rect 447138 267336 447194 267345
rect 440238 267271 440240 267280
rect 437478 267200 437534 267209
rect 437478 267135 437534 267144
rect 437492 267102 437520 267135
rect 437480 267096 437532 267102
rect 433338 267064 433394 267073
rect 437480 267038 437532 267044
rect 440068 267034 440096 267271
rect 440292 267271 440294 267280
rect 447138 267271 447194 267280
rect 440240 267242 440292 267248
rect 447152 267238 447180 267271
rect 503180 267238 503208 267407
rect 447140 267232 447192 267238
rect 445758 267200 445814 267209
rect 447140 267174 447192 267180
rect 503168 267232 503220 267238
rect 503168 267174 503220 267180
rect 445758 267135 445760 267144
rect 445812 267135 445814 267144
rect 445760 267106 445812 267112
rect 503548 267102 503576 267407
rect 503536 267096 503588 267102
rect 503536 267038 503588 267044
rect 516612 267034 516640 371350
rect 517532 354822 517560 460906
rect 517624 355502 517652 460974
rect 517612 355496 517664 355502
rect 517612 355438 517664 355444
rect 517520 354816 517572 354822
rect 517520 354758 517572 354764
rect 433338 266999 433340 267008
rect 433392 266999 433394 267008
rect 440056 267028 440108 267034
rect 433340 266970 433392 266976
rect 440056 266970 440108 266976
rect 516600 267028 516652 267034
rect 516600 266970 516652 266976
rect 437478 266656 437534 266665
rect 437478 266591 437534 266600
rect 437492 266422 437520 266591
rect 437480 266416 437532 266422
rect 436098 266384 436154 266393
rect 437480 266358 437532 266364
rect 436098 266319 436154 266328
rect 436112 263566 436140 266319
rect 436100 263560 436152 263566
rect 436100 263502 436152 263508
rect 500040 250708 500092 250714
rect 500040 250650 500092 250656
rect 499028 250572 499080 250578
rect 499028 250514 499080 250520
rect 427084 250504 427136 250510
rect 427084 250446 427136 250452
rect 499040 249937 499068 250514
rect 500052 249937 500080 250650
rect 510896 249960 510948 249966
rect 499026 249928 499082 249937
rect 499026 249863 499082 249872
rect 500038 249928 500094 249937
rect 500038 249863 500094 249872
rect 510894 249928 510896 249937
rect 510948 249928 510950 249937
rect 510894 249863 510950 249872
rect 412546 164928 412602 164937
rect 412546 164863 412602 164872
rect 393964 164212 394016 164218
rect 393964 164154 394016 164160
rect 393976 162081 394004 164154
rect 401598 163160 401654 163169
rect 401598 163095 401654 163104
rect 396078 162752 396134 162761
rect 396078 162687 396134 162696
rect 397458 162752 397514 162761
rect 397458 162687 397514 162696
rect 398838 162752 398894 162761
rect 398838 162687 398894 162696
rect 400218 162752 400274 162761
rect 400218 162687 400274 162696
rect 393962 162072 394018 162081
rect 393962 162007 394018 162016
rect 379980 161424 380032 161430
rect 379980 161366 380032 161372
rect 379992 160138 380020 161366
rect 379980 160132 380032 160138
rect 379980 160074 380032 160080
rect 380808 149048 380860 149054
rect 380808 148990 380860 148996
rect 379888 148980 379940 148986
rect 379888 148922 379940 148928
rect 379900 147694 379928 148922
rect 380820 148481 380848 148990
rect 380806 148472 380862 148481
rect 380256 148436 380308 148442
rect 380806 148407 380862 148416
rect 380256 148378 380308 148384
rect 380268 148306 380296 148378
rect 380256 148300 380308 148306
rect 380256 148242 380308 148248
rect 379888 147688 379940 147694
rect 379888 147630 379940 147636
rect 379978 146296 380034 146305
rect 379978 146231 380034 146240
rect 379796 56228 379848 56234
rect 379796 56170 379848 56176
rect 379992 56166 380020 146231
rect 393976 145382 394004 162007
rect 396092 145518 396120 162687
rect 396170 162208 396226 162217
rect 396170 162143 396226 162152
rect 396080 145512 396132 145518
rect 396080 145454 396132 145460
rect 396184 145450 396212 162143
rect 397472 145722 397500 162687
rect 398852 148510 398880 162687
rect 400232 148918 400260 162687
rect 400220 148912 400272 148918
rect 400220 148854 400272 148860
rect 401612 148578 401640 163095
rect 403070 162752 403126 162761
rect 403070 162687 403126 162696
rect 404358 162752 404414 162761
rect 404358 162687 404414 162696
rect 405738 162752 405794 162761
rect 405738 162687 405794 162696
rect 407210 162752 407266 162761
rect 407210 162687 407266 162696
rect 408314 162752 408370 162761
rect 408314 162687 408370 162696
rect 408498 162752 408554 162761
rect 408498 162687 408554 162696
rect 409878 162752 409934 162761
rect 409878 162687 409934 162696
rect 410614 162752 410670 162761
rect 410614 162687 410670 162696
rect 411350 162752 411406 162761
rect 411350 162687 411406 162696
rect 402978 162208 403034 162217
rect 402978 162143 403034 162152
rect 401600 148572 401652 148578
rect 401600 148514 401652 148520
rect 398840 148504 398892 148510
rect 398840 148446 398892 148452
rect 402992 145858 403020 162143
rect 403084 145926 403112 162687
rect 403072 145920 403124 145926
rect 403072 145862 403124 145868
rect 402980 145852 403032 145858
rect 402980 145794 403032 145800
rect 404372 145790 404400 162687
rect 405752 145994 405780 162687
rect 405740 145988 405792 145994
rect 405740 145930 405792 145936
rect 404360 145784 404412 145790
rect 404360 145726 404412 145732
rect 397460 145716 397512 145722
rect 397460 145658 397512 145664
rect 407224 145654 407252 162687
rect 408328 162110 408356 162687
rect 408316 162104 408368 162110
rect 408316 162046 408368 162052
rect 408512 146062 408540 162687
rect 409892 146130 409920 162687
rect 410628 162178 410656 162687
rect 411258 162208 411314 162217
rect 410616 162172 410668 162178
rect 411258 162143 411314 162152
rect 410616 162114 410668 162120
rect 411272 146266 411300 162143
rect 411260 146260 411312 146266
rect 411260 146202 411312 146208
rect 411364 146198 411392 162687
rect 412560 161537 412588 164863
rect 425978 164792 426034 164801
rect 425978 164727 426034 164736
rect 451002 164792 451058 164801
rect 451002 164727 451058 164736
rect 423494 164656 423550 164665
rect 423494 164591 423550 164600
rect 418434 164248 418490 164257
rect 418434 164183 418490 164192
rect 421010 164248 421066 164257
rect 421010 164183 421066 164192
rect 418448 164150 418476 164183
rect 418436 164144 418488 164150
rect 418436 164086 418488 164092
rect 421024 164082 421052 164183
rect 421012 164076 421064 164082
rect 421012 164018 421064 164024
rect 423508 163946 423536 164591
rect 425992 164422 426020 164727
rect 429750 164656 429806 164665
rect 429750 164591 429806 164600
rect 436926 164656 436982 164665
rect 436926 164591 436982 164600
rect 425980 164416 426032 164422
rect 425980 164358 426032 164364
rect 428186 164248 428242 164257
rect 428186 164183 428242 164192
rect 423496 163940 423548 163946
rect 423496 163882 423548 163888
rect 428200 163878 428228 164183
rect 428188 163872 428240 163878
rect 428188 163814 428240 163820
rect 416042 163160 416098 163169
rect 416042 163095 416098 163104
rect 413558 162752 413614 162761
rect 413558 162687 413614 162696
rect 414018 162752 414074 162761
rect 414018 162687 414074 162696
rect 415490 162752 415546 162761
rect 415490 162687 415546 162696
rect 413572 162042 413600 162687
rect 413560 162036 413612 162042
rect 413560 161978 413612 161984
rect 412546 161528 412602 161537
rect 412546 161463 412602 161472
rect 412730 161528 412786 161537
rect 412730 161463 412786 161472
rect 412744 148986 412772 161463
rect 412732 148980 412784 148986
rect 412732 148922 412784 148928
rect 414032 146305 414060 162687
rect 415308 162172 415360 162178
rect 415308 162114 415360 162120
rect 415320 162081 415348 162114
rect 415306 162072 415362 162081
rect 415306 162007 415362 162016
rect 414018 146296 414074 146305
rect 414018 146231 414074 146240
rect 411352 146192 411404 146198
rect 411352 146134 411404 146140
rect 409880 146124 409932 146130
rect 409880 146066 409932 146072
rect 408500 146056 408552 146062
rect 408500 145998 408552 146004
rect 415504 145897 415532 162687
rect 416056 161974 416084 163095
rect 429764 163062 429792 164591
rect 430946 164248 431002 164257
rect 430946 164183 431002 164192
rect 430960 164014 430988 164183
rect 430948 164008 431000 164014
rect 430948 163950 431000 163956
rect 429752 163056 429804 163062
rect 429752 162998 429804 163004
rect 431960 162988 432012 162994
rect 431960 162930 432012 162936
rect 431972 162761 432000 162930
rect 436940 162926 436968 164591
rect 451016 164354 451044 164727
rect 470966 164656 471022 164665
rect 470966 164591 471022 164600
rect 480902 164656 480958 164665
rect 480902 164591 480958 164600
rect 451004 164348 451056 164354
rect 451004 164290 451056 164296
rect 438860 163872 438912 163878
rect 438860 163814 438912 163820
rect 436928 162920 436980 162926
rect 436928 162862 436980 162868
rect 438872 162761 438900 163814
rect 470980 163674 471008 164591
rect 480916 164286 480944 164591
rect 480904 164280 480956 164286
rect 473450 164248 473506 164257
rect 473450 164183 473506 164192
rect 475842 164248 475898 164257
rect 475842 164183 475898 164192
rect 478418 164248 478474 164257
rect 480904 164222 480956 164228
rect 483386 164248 483442 164257
rect 478418 164183 478474 164192
rect 483386 164183 483442 164192
rect 473464 163742 473492 164183
rect 475856 163810 475884 164183
rect 475844 163804 475896 163810
rect 475844 163746 475896 163752
rect 473452 163736 473504 163742
rect 473452 163678 473504 163684
rect 470968 163668 471020 163674
rect 470968 163610 471020 163616
rect 478432 163606 478460 164183
rect 478420 163600 478472 163606
rect 478420 163542 478472 163548
rect 483400 163538 483428 164183
rect 516612 163878 516640 266970
rect 517532 249966 517560 354758
rect 517624 250714 517652 355438
rect 517716 355434 517744 461110
rect 519556 454714 519584 516122
rect 560956 511970 560984 572698
rect 580264 515432 580316 515438
rect 580264 515374 580316 515380
rect 560944 511964 560996 511970
rect 560944 511906 560996 511912
rect 580172 511964 580224 511970
rect 580172 511906 580224 511912
rect 580184 511329 580212 511906
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 520924 487212 520976 487218
rect 520924 487154 520976 487160
rect 519544 454708 519596 454714
rect 519544 454650 519596 454656
rect 518898 454200 518954 454209
rect 518898 454135 518954 454144
rect 517888 371884 517940 371890
rect 517888 371826 517940 371832
rect 517900 371346 517928 371826
rect 517888 371340 517940 371346
rect 517888 371282 517940 371288
rect 517796 371272 517848 371278
rect 517796 371214 517848 371220
rect 517704 355428 517756 355434
rect 517704 355370 517756 355376
rect 517612 250708 517664 250714
rect 517612 250650 517664 250656
rect 517624 250306 517652 250650
rect 517716 250578 517744 355370
rect 517808 267238 517836 371214
rect 517796 267232 517848 267238
rect 517796 267174 517848 267180
rect 517808 266422 517836 267174
rect 517900 267102 517928 371282
rect 518912 349217 518940 454135
rect 518990 393816 519046 393825
rect 518990 393751 519046 393760
rect 519004 370530 519032 393751
rect 519174 392184 519230 392193
rect 519174 392119 519230 392128
rect 519082 388104 519138 388113
rect 519082 388039 519138 388048
rect 518992 370524 519044 370530
rect 518992 370466 519044 370472
rect 518898 349208 518954 349217
rect 518898 349143 518954 349152
rect 517888 267096 517940 267102
rect 517888 267038 517940 267044
rect 517796 266416 517848 266422
rect 517796 266358 517848 266364
rect 517704 250572 517756 250578
rect 517704 250514 517756 250520
rect 517612 250300 517664 250306
rect 517612 250242 517664 250248
rect 517520 249960 517572 249966
rect 517520 249902 517572 249908
rect 516600 163872 516652 163878
rect 516600 163814 516652 163820
rect 517532 163674 517560 249902
rect 517716 248414 517744 250514
rect 517716 248386 517836 248414
rect 510528 163668 510580 163674
rect 510528 163610 510580 163616
rect 517520 163668 517572 163674
rect 517520 163610 517572 163616
rect 483388 163532 483440 163538
rect 483388 163474 483440 163480
rect 455786 163160 455842 163169
rect 455786 163095 455842 163104
rect 455800 162790 455828 163095
rect 458364 162852 458416 162858
rect 458364 162794 458416 162800
rect 455788 162784 455840 162790
rect 416778 162752 416834 162761
rect 416778 162687 416834 162696
rect 418158 162752 418214 162761
rect 418158 162687 418214 162696
rect 419538 162752 419594 162761
rect 419538 162687 419594 162696
rect 420918 162752 420974 162761
rect 420918 162687 420974 162696
rect 422298 162752 422354 162761
rect 422298 162687 422354 162696
rect 423678 162752 423734 162761
rect 423678 162687 423734 162696
rect 425058 162752 425114 162761
rect 425058 162687 425114 162696
rect 426438 162752 426494 162761
rect 426438 162687 426494 162696
rect 429106 162752 429162 162761
rect 429106 162687 429162 162696
rect 430578 162752 430634 162761
rect 430578 162687 430634 162696
rect 431958 162752 432014 162761
rect 431958 162687 432014 162696
rect 433338 162752 433394 162761
rect 433338 162687 433394 162696
rect 435730 162752 435786 162761
rect 435730 162687 435786 162696
rect 435914 162752 435970 162761
rect 435914 162687 435970 162696
rect 437478 162752 437534 162761
rect 437478 162687 437534 162696
rect 438490 162752 438546 162761
rect 438490 162687 438546 162696
rect 438858 162752 438914 162761
rect 438858 162687 438914 162696
rect 440882 162752 440938 162761
rect 440882 162687 440938 162696
rect 443458 162752 443514 162761
rect 443458 162687 443514 162696
rect 445850 162752 445906 162761
rect 445850 162687 445906 162696
rect 448242 162752 448298 162761
rect 448242 162687 448298 162696
rect 453394 162752 453450 162761
rect 458376 162761 458404 162794
rect 455788 162726 455840 162732
rect 458362 162752 458418 162761
rect 453394 162687 453396 162696
rect 416044 161968 416096 161974
rect 416044 161910 416096 161916
rect 415490 145888 415546 145897
rect 415490 145823 415546 145832
rect 416792 145761 416820 162687
rect 418172 159458 418200 162687
rect 418250 162208 418306 162217
rect 418250 162143 418252 162152
rect 418304 162143 418306 162152
rect 418252 162114 418304 162120
rect 419552 160002 419580 162687
rect 420932 160070 420960 162687
rect 420920 160064 420972 160070
rect 420920 160006 420972 160012
rect 419540 159996 419592 160002
rect 419540 159938 419592 159944
rect 418160 159452 418212 159458
rect 418160 159394 418212 159400
rect 416778 145752 416834 145761
rect 416778 145687 416834 145696
rect 407212 145648 407264 145654
rect 422312 145625 422340 162687
rect 423692 148442 423720 162687
rect 425072 161362 425100 162687
rect 426452 161430 426480 162687
rect 426530 162208 426586 162217
rect 426530 162143 426586 162152
rect 426440 161424 426492 161430
rect 426440 161366 426492 161372
rect 425060 161356 425112 161362
rect 425060 161298 425112 161304
rect 423680 148436 423732 148442
rect 423680 148378 423732 148384
rect 426544 147626 426572 162143
rect 428740 161560 428792 161566
rect 428740 161502 428792 161508
rect 428752 159390 428780 161502
rect 429120 161474 429148 162687
rect 429120 161446 429240 161474
rect 428740 159384 428792 159390
rect 428740 159326 428792 159332
rect 429212 149054 429240 161446
rect 430592 160886 430620 162687
rect 430580 160880 430632 160886
rect 430580 160822 430632 160828
rect 433352 160818 433380 162687
rect 433524 162240 433576 162246
rect 433524 162182 433576 162188
rect 434626 162208 434682 162217
rect 433536 162081 433564 162182
rect 434626 162143 434682 162152
rect 433522 162072 433578 162081
rect 433522 162007 433578 162016
rect 434640 161474 434668 162143
rect 435744 161566 435772 162687
rect 435928 162586 435956 162687
rect 435916 162580 435968 162586
rect 435916 162522 435968 162528
rect 435732 161560 435784 161566
rect 435732 161502 435784 161508
rect 437492 161474 437520 162687
rect 438504 162450 438532 162687
rect 438492 162444 438544 162450
rect 438492 162386 438544 162392
rect 434640 161446 434760 161474
rect 433340 160812 433392 160818
rect 433340 160754 433392 160760
rect 429200 149048 429252 149054
rect 429200 148990 429252 148996
rect 434732 148374 434760 161446
rect 437400 161446 437520 161474
rect 437400 160750 437428 161446
rect 437388 160744 437440 160750
rect 437388 160686 437440 160692
rect 434720 148368 434772 148374
rect 438872 148345 438900 162687
rect 440896 162314 440924 162687
rect 443472 162382 443500 162687
rect 445864 162518 445892 162687
rect 448256 162654 448284 162687
rect 453448 162687 453450 162696
rect 458362 162687 458418 162696
rect 503258 162752 503314 162761
rect 503258 162687 503314 162696
rect 453396 162658 453448 162664
rect 448244 162648 448296 162654
rect 448244 162590 448296 162596
rect 445852 162512 445904 162518
rect 445852 162454 445904 162460
rect 443460 162376 443512 162382
rect 443460 162318 443512 162324
rect 503272 162314 503300 162687
rect 503626 162616 503682 162625
rect 503626 162551 503682 162560
rect 440884 162308 440936 162314
rect 440884 162250 440936 162256
rect 503260 162308 503312 162314
rect 503260 162250 503312 162256
rect 503640 162178 503668 162551
rect 503628 162172 503680 162178
rect 503628 162114 503680 162120
rect 434720 148310 434772 148316
rect 438858 148336 438914 148345
rect 438858 148271 438914 148280
rect 426532 147620 426584 147626
rect 426532 147562 426584 147568
rect 500224 146192 500276 146198
rect 500224 146134 500276 146140
rect 498660 146124 498712 146130
rect 498660 146066 498712 146072
rect 407212 145590 407264 145596
rect 422298 145616 422354 145625
rect 422298 145551 422354 145560
rect 396172 145444 396224 145450
rect 396172 145386 396224 145392
rect 393964 145376 394016 145382
rect 393964 145318 394016 145324
rect 498672 144945 498700 146066
rect 500236 144945 500264 146134
rect 510540 145586 510568 163610
rect 517612 162852 517664 162858
rect 517612 162794 517664 162800
rect 517520 162784 517572 162790
rect 517520 162726 517572 162732
rect 517532 162314 517560 162726
rect 517520 162308 517572 162314
rect 517520 162250 517572 162256
rect 510528 145580 510580 145586
rect 510528 145522 510580 145528
rect 510540 145466 510568 145522
rect 510618 145480 510674 145489
rect 510540 145438 510618 145466
rect 510618 145415 510674 145424
rect 498658 144936 498714 144945
rect 498658 144871 498714 144880
rect 500222 144936 500278 144945
rect 500222 144871 500278 144880
rect 396078 59800 396134 59809
rect 396078 59735 396134 59744
rect 397090 59800 397146 59809
rect 397090 59735 397092 59744
rect 396092 59702 396120 59735
rect 397144 59735 397146 59744
rect 416962 59800 417018 59809
rect 416962 59735 417018 59744
rect 418434 59800 418490 59809
rect 418434 59735 418490 59744
rect 423954 59800 424010 59809
rect 423954 59735 424010 59744
rect 397092 59706 397144 59712
rect 396080 59696 396132 59702
rect 396080 59638 396132 59644
rect 403070 59664 403126 59673
rect 403070 59599 403126 59608
rect 404174 59664 404230 59673
rect 404174 59599 404230 59608
rect 412546 59664 412602 59673
rect 412546 59599 412602 59608
rect 403084 59294 403112 59599
rect 403072 59288 403124 59294
rect 403072 59230 403124 59236
rect 404188 58614 404216 59599
rect 404176 58608 404228 58614
rect 404176 58550 404228 58556
rect 397458 57896 397514 57905
rect 397458 57831 397514 57840
rect 399482 57896 399538 57905
rect 399482 57831 399538 57840
rect 400218 57896 400274 57905
rect 400218 57831 400274 57840
rect 401690 57896 401746 57905
rect 401690 57831 401746 57840
rect 404358 57896 404414 57905
rect 404358 57831 404414 57840
rect 405830 57896 405886 57905
rect 405830 57831 405886 57840
rect 407210 57896 407266 57905
rect 407210 57831 407266 57840
rect 408314 57896 408370 57905
rect 408314 57831 408370 57840
rect 408682 57896 408738 57905
rect 408682 57831 408738 57840
rect 409878 57896 409934 57905
rect 409878 57831 409934 57840
rect 411350 57896 411406 57905
rect 411350 57831 411406 57840
rect 379980 56160 380032 56166
rect 379980 56102 380032 56108
rect 379428 56092 379480 56098
rect 379428 56034 379480 56040
rect 379244 55956 379296 55962
rect 379244 55898 379296 55904
rect 397472 55146 397500 57831
rect 399496 55894 399524 57831
rect 399484 55888 399536 55894
rect 399484 55830 399536 55836
rect 397460 55140 397512 55146
rect 397460 55082 397512 55088
rect 378784 54596 378836 54602
rect 378784 54538 378836 54544
rect 400232 54534 400260 57831
rect 401704 56574 401732 57831
rect 401692 56568 401744 56574
rect 401692 56510 401744 56516
rect 404372 54670 404400 57831
rect 405844 54738 405872 57831
rect 405832 54732 405884 54738
rect 405832 54674 405884 54680
rect 404360 54664 404412 54670
rect 404360 54606 404412 54612
rect 407224 54602 407252 57831
rect 408328 55826 408356 57831
rect 408696 56030 408724 57831
rect 408684 56024 408736 56030
rect 408684 55966 408736 55972
rect 408316 55820 408368 55826
rect 408316 55762 408368 55768
rect 409892 54806 409920 57831
rect 411258 56944 411314 56953
rect 411258 56879 411314 56888
rect 411272 55962 411300 56879
rect 411260 55956 411312 55962
rect 411260 55898 411312 55904
rect 411364 54874 411392 57831
rect 412560 56953 412588 59599
rect 416976 59566 417004 59735
rect 418160 59628 418212 59634
rect 418160 59570 418212 59576
rect 416964 59560 417016 59566
rect 418172 59537 418200 59570
rect 416964 59502 417016 59508
rect 418158 59528 418214 59537
rect 418158 59463 418214 59472
rect 418448 59430 418476 59735
rect 419446 59664 419502 59673
rect 419446 59599 419502 59608
rect 421746 59664 421802 59673
rect 421746 59599 421802 59608
rect 423494 59664 423550 59673
rect 423494 59599 423550 59608
rect 418436 59424 418488 59430
rect 418436 59366 418488 59372
rect 419460 59226 419488 59599
rect 420642 59528 420698 59537
rect 420642 59463 420698 59472
rect 419448 59220 419500 59226
rect 419448 59162 419500 59168
rect 420656 59158 420684 59463
rect 420644 59152 420696 59158
rect 420644 59094 420696 59100
rect 421760 59090 421788 59599
rect 421748 59084 421800 59090
rect 421748 59026 421800 59032
rect 423508 58954 423536 59599
rect 423968 59498 423996 59735
rect 503258 59664 503314 59673
rect 503258 59599 503314 59608
rect 423956 59492 424008 59498
rect 423956 59434 424008 59440
rect 425242 59392 425298 59401
rect 425242 59327 425298 59336
rect 425978 59392 426034 59401
rect 425978 59327 426034 59336
rect 428186 59392 428242 59401
rect 428186 59327 428242 59336
rect 465906 59392 465962 59401
rect 465906 59327 465962 59336
rect 425256 59022 425284 59327
rect 425244 59016 425296 59022
rect 425244 58958 425296 58964
rect 423496 58948 423548 58954
rect 423496 58890 423548 58896
rect 425992 58886 426020 59327
rect 425980 58880 426032 58886
rect 425980 58822 426032 58828
rect 428200 58682 428228 59327
rect 465920 58818 465948 59327
rect 485962 59256 486018 59265
rect 485962 59191 486018 59200
rect 465908 58812 465960 58818
rect 465908 58754 465960 58760
rect 485976 58750 486004 59191
rect 485964 58744 486016 58750
rect 485964 58686 486016 58692
rect 428188 58676 428240 58682
rect 428188 58618 428240 58624
rect 478420 57928 478472 57934
rect 414570 57896 414626 57905
rect 414570 57831 414626 57840
rect 415490 57896 415546 57905
rect 415490 57831 415546 57840
rect 416042 57896 416098 57905
rect 416042 57831 416098 57840
rect 426438 57896 426494 57905
rect 426438 57831 426494 57840
rect 427634 57896 427690 57905
rect 427634 57831 427690 57840
rect 427818 57896 427874 57905
rect 427818 57831 427874 57840
rect 429198 57896 429254 57905
rect 429198 57831 429254 57840
rect 430578 57896 430634 57905
rect 430578 57831 430634 57840
rect 431958 57896 432014 57905
rect 431958 57831 432014 57840
rect 433430 57896 433486 57905
rect 433430 57831 433486 57840
rect 435914 57896 435970 57905
rect 435914 57831 435970 57840
rect 436098 57896 436154 57905
rect 436098 57831 436154 57840
rect 438306 57896 438362 57905
rect 438306 57831 438362 57840
rect 438490 57896 438546 57905
rect 438490 57831 438546 57840
rect 438858 57896 438914 57905
rect 438858 57831 438914 57840
rect 440882 57896 440938 57905
rect 440882 57831 440938 57840
rect 443458 57896 443514 57905
rect 443458 57831 443460 57840
rect 412546 56944 412602 56953
rect 412546 56879 412602 56888
rect 412638 56808 412694 56817
rect 412638 56743 412694 56752
rect 412652 56098 412680 56743
rect 414584 56166 414612 57831
rect 415504 57254 415532 57831
rect 416056 57322 416084 57831
rect 416044 57316 416096 57322
rect 416044 57258 416096 57264
rect 415492 57248 415544 57254
rect 415492 57190 415544 57196
rect 426452 56234 426480 57831
rect 427648 56302 427676 57831
rect 427636 56296 427688 56302
rect 427636 56238 427688 56244
rect 426440 56228 426492 56234
rect 426440 56170 426492 56176
rect 414572 56160 414624 56166
rect 414572 56102 414624 56108
rect 412640 56092 412692 56098
rect 412640 56034 412692 56040
rect 427832 55049 427860 57831
rect 427818 55040 427874 55049
rect 427818 54975 427874 54984
rect 429212 54942 429240 57831
rect 430592 55010 430620 57831
rect 430948 57384 431000 57390
rect 430948 57326 431000 57332
rect 430960 57225 430988 57326
rect 430946 57216 431002 57225
rect 430946 57151 431002 57160
rect 431972 55078 432000 57831
rect 433338 57216 433394 57225
rect 433338 57151 433394 57160
rect 433352 56370 433380 57151
rect 433340 56364 433392 56370
rect 433340 56306 433392 56312
rect 431960 55072 432012 55078
rect 431960 55014 432012 55020
rect 430580 55004 430632 55010
rect 430580 54946 430632 54952
rect 429200 54936 429252 54942
rect 429200 54878 429252 54884
rect 411352 54868 411404 54874
rect 411352 54810 411404 54816
rect 409880 54800 409932 54806
rect 409880 54742 409932 54748
rect 407212 54596 407264 54602
rect 407212 54538 407264 54544
rect 373724 54528 373776 54534
rect 373724 54470 373776 54476
rect 400220 54528 400272 54534
rect 400220 54470 400272 54476
rect 433444 54466 433472 57831
rect 435928 57526 435956 57831
rect 435916 57520 435968 57526
rect 435916 57462 435968 57468
rect 433524 57452 433576 57458
rect 433524 57394 433576 57400
rect 433536 57225 433564 57394
rect 433522 57216 433578 57225
rect 433522 57151 433578 57160
rect 435730 57216 435786 57225
rect 435730 57151 435786 57160
rect 435744 56438 435772 57151
rect 435732 56432 435784 56438
rect 435732 56374 435784 56380
rect 436112 55214 436140 57831
rect 438320 56506 438348 57831
rect 438504 57594 438532 57831
rect 438492 57588 438544 57594
rect 438492 57530 438544 57536
rect 438308 56500 438360 56506
rect 438308 56442 438360 56448
rect 436100 55208 436152 55214
rect 438872 55185 438900 57831
rect 440896 57798 440924 57831
rect 443512 57831 443514 57840
rect 445850 57896 445906 57905
rect 445850 57831 445906 57840
rect 451002 57896 451058 57905
rect 451002 57831 451058 57840
rect 478418 57896 478420 57905
rect 478472 57896 478474 57905
rect 503272 57866 503300 59599
rect 503352 57928 503404 57934
rect 503350 57896 503352 57905
rect 503404 57896 503406 57905
rect 478418 57831 478474 57840
rect 503260 57860 503312 57866
rect 443460 57802 443512 57808
rect 440884 57792 440936 57798
rect 440884 57734 440936 57740
rect 445864 57730 445892 57831
rect 445852 57724 445904 57730
rect 445852 57666 445904 57672
rect 451016 57662 451044 57831
rect 517532 57866 517560 162250
rect 517624 162178 517652 162794
rect 517612 162172 517664 162178
rect 517612 162114 517664 162120
rect 517624 57934 517652 162114
rect 517808 151814 517836 248386
rect 517900 162858 517928 267038
rect 517980 266416 518032 266422
rect 517980 266358 518032 266364
rect 517888 162852 517940 162858
rect 517888 162794 517940 162800
rect 517992 162790 518020 266358
rect 518072 250300 518124 250306
rect 518072 250242 518124 250248
rect 517980 162784 518032 162790
rect 517980 162726 518032 162732
rect 517716 151786 517836 151814
rect 517716 146130 517744 151786
rect 518084 146198 518112 250242
rect 518912 244225 518940 349143
rect 519004 289377 519032 370466
rect 519096 369170 519124 388039
rect 519084 369164 519136 369170
rect 519084 369106 519136 369112
rect 518990 289368 519046 289377
rect 518990 289303 519046 289312
rect 518990 288416 519046 288425
rect 518990 288351 519046 288360
rect 519004 287201 519032 288351
rect 518990 287192 519046 287201
rect 518990 287127 519046 287136
rect 518898 244216 518954 244225
rect 518898 244151 518954 244160
rect 519004 182753 519032 287127
rect 519096 284209 519124 369106
rect 519188 367810 519216 392119
rect 519266 390824 519322 390833
rect 519266 390759 519322 390768
rect 519176 367804 519228 367810
rect 519176 367746 519228 367752
rect 519188 288425 519216 367746
rect 519280 359514 519308 390759
rect 519358 389328 519414 389337
rect 519358 389263 519414 389272
rect 519268 359508 519320 359514
rect 519268 359450 519320 359456
rect 519174 288416 519230 288425
rect 519174 288351 519230 288360
rect 519280 285841 519308 359450
rect 519372 358154 519400 389263
rect 520936 388482 520964 487154
rect 580276 458153 580304 515374
rect 580262 458144 580318 458153
rect 580262 458079 580318 458088
rect 580264 454708 580316 454714
rect 580264 454650 580316 454656
rect 580276 404977 580304 454650
rect 580262 404968 580318 404977
rect 580262 404903 580318 404912
rect 520924 388476 520976 388482
rect 520924 388418 520976 388424
rect 580356 388476 580408 388482
rect 580356 388418 580408 388424
rect 580264 371272 580316 371278
rect 580264 371214 580316 371220
rect 519360 358148 519412 358154
rect 519360 358090 519412 358096
rect 519266 285832 519322 285841
rect 519266 285767 519322 285776
rect 519372 284889 519400 358090
rect 580276 325281 580304 371214
rect 580368 351937 580396 388418
rect 580446 378448 580502 378457
rect 580446 378383 580502 378392
rect 580460 371890 580488 378383
rect 580448 371884 580500 371890
rect 580448 371826 580500 371832
rect 580354 351928 580410 351937
rect 580354 351863 580410 351872
rect 580262 325272 580318 325281
rect 580262 325207 580318 325216
rect 519542 289368 519598 289377
rect 519542 289303 519598 289312
rect 519358 284880 519414 284889
rect 519358 284815 519414 284824
rect 519082 284200 519138 284209
rect 519082 284135 519138 284144
rect 519096 282946 519124 284135
rect 519084 282940 519136 282946
rect 519084 282882 519136 282888
rect 518990 182744 519046 182753
rect 518990 182679 519046 182688
rect 519096 180794 519124 282882
rect 519372 277394 519400 284815
rect 519372 277366 519492 277394
rect 519358 244216 519414 244225
rect 519358 244151 519414 244160
rect 519266 184920 519322 184929
rect 519266 184855 519322 184864
rect 519174 182744 519230 182753
rect 519174 182679 519230 182688
rect 518912 180766 519124 180794
rect 518912 178809 518940 180766
rect 518990 179480 519046 179489
rect 518990 179415 519046 179424
rect 518898 178800 518954 178809
rect 518898 178735 518954 178744
rect 518072 146192 518124 146198
rect 518072 146134 518124 146140
rect 518256 146192 518308 146198
rect 518256 146134 518308 146140
rect 517704 146124 517756 146130
rect 517704 146066 517756 146072
rect 517716 145654 517744 146066
rect 517704 145648 517756 145654
rect 517704 145590 517756 145596
rect 518268 145586 518296 146134
rect 518256 145580 518308 145586
rect 518256 145522 518308 145528
rect 518912 74225 518940 178735
rect 519004 75449 519032 179415
rect 519188 78305 519216 182679
rect 519280 79937 519308 184855
rect 519372 139369 519400 244151
rect 519464 179489 519492 277366
rect 519556 184929 519584 289303
rect 519634 285832 519690 285841
rect 519634 285767 519690 285776
rect 519542 184920 519598 184929
rect 519542 184855 519598 184864
rect 519648 183682 519676 285767
rect 520186 284880 520242 284889
rect 520186 284815 520242 284824
rect 520200 284374 520228 284815
rect 520188 284368 520240 284374
rect 520188 284310 520240 284316
rect 580264 284368 580316 284374
rect 580264 284310 580316 284316
rect 580276 232393 580304 284310
rect 580356 282940 580408 282946
rect 580356 282882 580408 282888
rect 580368 272241 580396 282882
rect 580354 272232 580410 272241
rect 580354 272167 580410 272176
rect 580262 232384 580318 232393
rect 580262 232319 580318 232328
rect 580354 192536 580410 192545
rect 580354 192471 580410 192480
rect 519556 183654 519676 183682
rect 519556 182170 519584 183654
rect 520186 182744 520242 182753
rect 520186 182679 520242 182688
rect 520200 182238 520228 182679
rect 520188 182232 520240 182238
rect 520188 182174 520240 182180
rect 580264 182232 580316 182238
rect 580264 182174 580316 182180
rect 519544 182164 519596 182170
rect 519544 182106 519596 182112
rect 519556 181393 519584 182106
rect 519542 181384 519598 181393
rect 519542 181319 519598 181328
rect 519450 179480 519506 179489
rect 519450 179415 519506 179424
rect 519358 139360 519414 139369
rect 519358 139295 519414 139304
rect 519266 79928 519322 79937
rect 519266 79863 519322 79872
rect 519174 78296 519230 78305
rect 519174 78231 519230 78240
rect 519556 76809 519584 181319
rect 580276 152697 580304 182174
rect 580368 182170 580396 192471
rect 580356 182164 580408 182170
rect 580356 182106 580408 182112
rect 580262 152688 580318 152697
rect 580262 152623 580318 152632
rect 580356 145648 580408 145654
rect 580356 145590 580408 145596
rect 580264 145580 580316 145586
rect 580264 145522 580316 145528
rect 520188 80028 520240 80034
rect 520188 79970 520240 79976
rect 520200 79937 520228 79970
rect 520186 79928 520242 79937
rect 520186 79863 520242 79872
rect 519542 76800 519598 76809
rect 519542 76735 519598 76744
rect 518990 75440 519046 75449
rect 518990 75375 519046 75384
rect 518898 74216 518954 74225
rect 518898 74151 518954 74160
rect 517612 57928 517664 57934
rect 517612 57870 517664 57876
rect 503350 57831 503406 57840
rect 517520 57860 517572 57866
rect 503260 57802 503312 57808
rect 517520 57802 517572 57808
rect 451004 57656 451056 57662
rect 451004 57598 451056 57604
rect 436100 55150 436152 55156
rect 438858 55176 438914 55185
rect 438858 55111 438914 55120
rect 373632 54460 373684 54466
rect 373632 54402 373684 54408
rect 433432 54460 433484 54466
rect 433432 54402 433484 54408
rect 580276 33153 580304 145522
rect 580368 73001 580396 145590
rect 580446 112840 580502 112849
rect 580446 112775 580502 112784
rect 580460 80034 580488 112775
rect 580448 80028 580500 80034
rect 580448 79970 580500 79976
rect 580354 72992 580410 73001
rect 580354 72927 580410 72936
rect 580262 33144 580318 33153
rect 580262 33079 580318 33088
rect 150622 3431 150678 3440
rect 366364 3460 366416 3466
rect 150636 480 150664 3431
rect 366364 3402 366416 3408
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 632032 3570 632088
rect 3422 579944 3478 580000
rect 2962 410488 3018 410544
rect 3330 358400 3386 358456
rect 3054 201864 3110 201920
rect 3606 514800 3662 514856
rect 3606 475360 3662 475416
rect 3606 462576 3662 462632
rect 3514 97552 3570 97608
rect 3422 58520 3478 58576
rect 42062 632032 42118 632088
rect 57702 620608 57758 620664
rect 57518 614352 57574 614408
rect 57426 589872 57482 589928
rect 57334 586336 57390 586392
rect 57058 577632 57114 577688
rect 57150 574912 57206 574968
rect 57334 571512 57390 571568
rect 57242 565392 57298 565448
rect 57610 593408 57666 593464
rect 57518 583616 57574 583672
rect 59266 617752 59322 617808
rect 59082 611632 59138 611688
rect 58898 608232 58954 608288
rect 57886 599528 57942 599584
rect 57886 595992 57942 596048
rect 58530 568792 58586 568848
rect 58806 581032 58862 581088
rect 58990 602112 59046 602168
rect 59174 605512 59230 605568
rect 59542 562732 59598 562788
rect 120814 598304 120870 598360
rect 120998 576816 121054 576872
rect 121458 570968 121514 571024
rect 121090 564848 121146 564904
rect 121182 562128 121238 562184
rect 121734 613808 121790 613864
rect 121918 611088 121974 611144
rect 121826 601568 121882 601624
rect 122194 586608 122250 586664
rect 122102 583208 122158 583264
rect 122010 580488 122066 580544
rect 122930 619928 122986 619984
rect 123114 617208 123170 617264
rect 123022 607688 123078 607744
rect 123206 604968 123262 605024
rect 123390 595448 123446 595504
rect 123298 592728 123354 592784
rect 124126 589364 124128 589384
rect 124128 589364 124180 589384
rect 124180 589364 124182 589384
rect 124126 589328 124182 589364
rect 123482 574368 123538 574424
rect 123574 568248 123630 568304
rect 137374 620608 137430 620664
rect 136730 608232 136786 608288
rect 137282 594768 137338 594824
rect 136730 589872 136786 589928
rect 136730 577632 136786 577688
rect 137650 611632 137706 611688
rect 137466 574912 137522 574968
rect 137558 571512 137614 571568
rect 281078 632168 281134 632224
rect 137834 599528 137890 599584
rect 139030 617752 139086 617808
rect 138846 605512 138902 605568
rect 137926 596128 137982 596184
rect 137926 594768 137982 594824
rect 137926 593408 137982 593464
rect 137834 583752 137890 583808
rect 138754 587152 138810 587208
rect 138662 581032 138718 581088
rect 138570 568792 138626 568848
rect 138478 565392 138534 565448
rect 138938 602112 138994 602168
rect 139214 614352 139270 614408
rect 139398 562740 139454 562796
rect 200762 598304 200818 598360
rect 201590 619928 201646 619984
rect 201498 570968 201554 571024
rect 201130 568248 201186 568304
rect 201222 562128 201278 562184
rect 201774 613808 201830 613864
rect 201866 604968 201922 605024
rect 201958 592728 202014 592784
rect 202142 586608 202198 586664
rect 202050 583208 202106 583264
rect 202878 617208 202934 617264
rect 202326 580488 202382 580544
rect 203062 611088 203118 611144
rect 202970 607688 203026 607744
rect 203154 601568 203210 601624
rect 203062 595448 203118 595504
rect 203246 589348 203302 589384
rect 203246 589328 203248 589348
rect 203248 589328 203300 589348
rect 203300 589328 203302 589348
rect 203338 577088 203394 577144
rect 203246 574368 203302 574424
rect 203430 564848 203486 564904
rect 216678 620608 216734 620664
rect 216678 617752 216734 617808
rect 215942 611632 215998 611688
rect 216678 608232 216734 608288
rect 217230 602112 217286 602168
rect 216678 593428 216734 593464
rect 216678 593408 216680 593428
rect 216680 593408 216732 593428
rect 216732 593408 216734 593428
rect 216678 589872 216734 589928
rect 216678 587152 216734 587208
rect 216034 577632 216090 577688
rect 216678 574912 216734 574968
rect 216678 571512 216734 571568
rect 217138 562672 217194 562728
rect 217690 614352 217746 614408
rect 217414 583752 217470 583808
rect 217782 599528 217838 599584
rect 217690 581032 217746 581088
rect 217598 565392 217654 565448
rect 218702 596128 218758 596184
rect 219254 605512 219310 605568
rect 219162 568792 219218 568848
rect 239402 542952 239458 543008
rect 241518 542544 241574 542600
rect 248694 542680 248750 542736
rect 255134 543224 255190 543280
rect 256514 543088 256570 543144
rect 264426 541048 264482 541104
rect 280894 616936 280950 616992
rect 280986 594904 281042 594960
rect 281906 619928 281962 619984
rect 281630 611088 281686 611144
rect 281170 592728 281226 592784
rect 281538 568248 281594 568304
rect 281262 564848 281318 564904
rect 281722 586608 281778 586664
rect 281814 580488 281870 580544
rect 282918 613808 282974 613864
rect 281998 562128 282054 562184
rect 283010 607688 283066 607744
rect 283194 604968 283250 605024
rect 283102 601568 283158 601624
rect 283286 598848 283342 598904
rect 283654 589348 283710 589384
rect 283654 589328 283656 589348
rect 283656 589328 283708 589348
rect 283708 589328 283710 589348
rect 283378 583208 283434 583264
rect 283562 577088 283618 577144
rect 283470 574368 283526 574424
rect 283654 570968 283710 571024
rect 285034 543088 285090 543144
rect 284298 541592 284354 541648
rect 285954 542816 286010 542872
rect 286690 542408 286746 542464
rect 291658 541320 291714 541376
rect 294510 541184 294566 541240
rect 300214 542680 300270 542736
rect 300214 518744 300270 518800
rect 301502 542408 301558 542464
rect 57702 509924 57758 509960
rect 57702 509904 57704 509924
rect 57704 509904 57756 509924
rect 57756 509904 57758 509924
rect 57886 509904 57942 509960
rect 42154 373904 42210 373960
rect 42614 466248 42670 466304
rect 302330 532344 302386 532400
rect 302606 517384 302662 517440
rect 317786 629584 317842 629640
rect 317602 625232 317658 625288
rect 317970 620064 318026 620120
rect 317970 615576 318026 615632
rect 317878 610544 317934 610600
rect 317970 606056 318026 606112
rect 317602 601024 317658 601080
rect 317602 596400 317658 596456
rect 317418 586508 317420 586528
rect 317420 586508 317472 586528
rect 317472 586508 317474 586528
rect 317418 586472 317474 586508
rect 317970 582528 318026 582584
rect 317878 577224 317934 577280
rect 317970 571784 318026 571840
rect 317050 568248 317106 568304
rect 317418 557640 317474 557696
rect 317970 553444 318026 553480
rect 317970 553424 317972 553444
rect 317972 553424 318024 553444
rect 318024 553424 318026 553444
rect 317970 549072 318026 549128
rect 312542 518472 312598 518528
rect 314198 541320 314254 541376
rect 317970 543804 317972 543824
rect 317972 543804 318024 543824
rect 318024 543804 318026 543824
rect 317970 543768 318026 543804
rect 318798 592728 318854 592784
rect 318338 562264 318394 562320
rect 319534 632304 319590 632360
rect 346398 632032 346454 632088
rect 392122 632304 392178 632360
rect 328090 630808 328146 630864
rect 405370 630672 405426 630728
rect 428370 558184 428426 558240
rect 318246 543224 318302 543280
rect 317050 542816 317106 542872
rect 316774 541592 316830 541648
rect 316958 541184 317014 541240
rect 318062 539280 318118 539336
rect 317602 534928 317658 534984
rect 317602 529760 317658 529816
rect 317694 525408 317750 525464
rect 318246 520104 318302 520160
rect 319718 518336 319774 518392
rect 337658 518336 337714 518392
rect 427818 520240 427874 520296
rect 356242 518472 356298 518528
rect 374458 518608 374514 518664
rect 302238 502424 302294 502480
rect 302882 487464 302938 487520
rect 366362 480800 366418 480856
rect 43258 373768 43314 373824
rect 46846 475904 46902 475960
rect 43994 472912 44050 472968
rect 46478 475496 46534 475552
rect 46294 267416 46350 267472
rect 46294 266328 46350 266384
rect 46478 266328 46534 266384
rect 47490 374992 47546 375048
rect 47950 266872 48006 266928
rect 47858 249056 47914 249112
rect 48870 267280 48926 267336
rect 48870 266328 48926 266384
rect 49146 266328 49202 266384
rect 50894 477536 50950 477592
rect 50342 475632 50398 475688
rect 50802 465976 50858 466032
rect 50710 459584 50766 459640
rect 50986 462984 51042 463040
rect 50986 268368 51042 268424
rect 50710 162560 50766 162616
rect 51538 144744 51594 144800
rect 52366 375264 52422 375320
rect 52458 374856 52514 374912
rect 53470 477536 53526 477592
rect 53470 466112 53526 466168
rect 52918 267008 52974 267064
rect 53562 375264 53618 375320
rect 53746 459584 53802 459640
rect 54390 269048 54446 269104
rect 53746 268504 53802 268560
rect 55862 472504 55918 472560
rect 53746 146240 53802 146296
rect 55678 415248 55734 415304
rect 55494 375264 55550 375320
rect 55586 372952 55642 373008
rect 55678 372680 55734 372736
rect 56966 412256 57022 412312
rect 57058 410352 57114 410408
rect 57058 408584 57114 408640
rect 56966 407360 57022 407416
rect 57058 405748 57114 405784
rect 57058 405728 57060 405748
rect 57060 405728 57112 405748
rect 57112 405728 57114 405748
rect 57058 404388 57114 404424
rect 57058 404368 57060 404388
rect 57060 404368 57112 404388
rect 57112 404368 57114 404388
rect 56966 403028 57022 403064
rect 56966 403008 56968 403028
rect 56968 403008 57020 403028
rect 57020 403008 57022 403028
rect 56966 384956 56968 384976
rect 56968 384956 57020 384976
rect 57020 384956 57022 384976
rect 56966 384920 57022 384956
rect 56874 383288 56930 383344
rect 57150 383016 57206 383072
rect 56506 372816 56562 372872
rect 56690 303592 56746 303648
rect 56782 302232 56838 302288
rect 56690 198736 56746 198792
rect 57150 304952 57206 305008
rect 57058 300464 57114 300520
rect 56966 268912 57022 268968
rect 56782 197376 56838 197432
rect 56046 145560 56102 145616
rect 56874 160112 56930 160168
rect 56322 146240 56378 146296
rect 57426 306856 57482 306912
rect 57242 278704 57298 278760
rect 57242 262248 57298 262304
rect 57610 302232 57666 302288
rect 57334 201864 57390 201920
rect 57150 200912 57206 200968
rect 57058 195200 57114 195256
rect 57058 147500 57060 147520
rect 57060 147500 57112 147520
rect 57112 147500 57114 147520
rect 57058 147464 57114 147500
rect 56414 145832 56470 145888
rect 56322 145560 56378 145616
rect 56874 68040 56930 68096
rect 57334 197376 57390 197432
rect 57242 97416 57298 97472
rect 57150 96464 57206 96520
rect 57518 301280 57574 301336
rect 58622 372680 58678 372736
rect 57886 305904 57942 305960
rect 57886 304952 57942 305008
rect 57794 303592 57850 303648
rect 57702 300464 57758 300520
rect 57518 298152 57574 298208
rect 57426 196016 57482 196072
rect 57426 195200 57482 195256
rect 57334 93336 57390 93392
rect 57886 278704 57942 278760
rect 57610 198736 57666 198792
rect 57518 193160 57574 193216
rect 57426 90480 57482 90536
rect 57702 196016 57758 196072
rect 57610 93744 57666 93800
rect 58714 279928 58770 279984
rect 58990 472776 59046 472832
rect 58806 278024 58862 278080
rect 57886 173304 57942 173360
rect 57794 173032 57850 173088
rect 57702 91024 57758 91080
rect 57518 88168 57574 88224
rect 58622 249736 58678 249792
rect 59082 463256 59138 463312
rect 58990 175208 59046 175264
rect 58622 145968 58678 146024
rect 57886 68856 57942 68912
rect 2778 19352 2834 19408
rect 59358 407768 59414 407824
rect 59450 372952 59506 373008
rect 60002 463120 60058 463176
rect 66258 478216 66314 478272
rect 66258 477808 66314 477864
rect 66350 475904 66406 475960
rect 67914 461624 67970 461680
rect 67822 460672 67878 460728
rect 67638 459040 67694 459096
rect 69202 460808 69258 460864
rect 72054 478760 72110 478816
rect 70582 466248 70638 466304
rect 70490 463392 70546 463448
rect 72514 477944 72570 478000
rect 73158 478780 73214 478816
rect 73158 478760 73160 478780
rect 73160 478760 73212 478780
rect 73212 478760 73214 478780
rect 73158 478624 73214 478680
rect 73434 478896 73490 478952
rect 73250 461488 73306 461544
rect 74630 478352 74686 478408
rect 76010 478216 76066 478272
rect 76470 477808 76526 477864
rect 77758 478624 77814 478680
rect 74630 460400 74686 460456
rect 77390 460536 77446 460592
rect 75918 460264 75974 460320
rect 79506 478760 79562 478816
rect 80794 478080 80850 478136
rect 81254 472912 81310 472968
rect 81530 465840 81586 465896
rect 84290 465976 84346 466032
rect 85762 466112 85818 466168
rect 78678 460128 78734 460184
rect 74538 459992 74594 460048
rect 91190 463256 91246 463312
rect 92662 463120 92718 463176
rect 95790 472776 95846 472832
rect 93950 462984 94006 463040
rect 94042 462848 94098 462904
rect 69110 458904 69166 458960
rect 102230 465704 102286 465760
rect 107750 478896 107806 478952
rect 116306 474000 116362 474056
rect 121366 475768 121422 475824
rect 120906 475632 120962 475688
rect 120446 475496 120502 475552
rect 121826 472504 121882 472560
rect 122654 472640 122710 472696
rect 124310 469920 124366 469976
rect 124218 465704 124274 465760
rect 69018 458768 69074 458824
rect 128542 469784 128598 469840
rect 145562 478216 145618 478272
rect 145102 478080 145158 478136
rect 146022 471280 146078 471336
rect 143630 468424 143686 468480
rect 147310 478488 147366 478544
rect 148230 478352 148286 478408
rect 150438 474136 150494 474192
rect 153106 476720 153162 476776
rect 152646 472504 152702 472560
rect 151726 471144 151782 471200
rect 150438 468560 150494 468616
rect 147678 467064 147734 467120
rect 146482 462984 146538 463040
rect 146298 462848 146354 462904
rect 143722 460264 143778 460320
rect 155682 475496 155738 475552
rect 153290 469784 153346 469840
rect 155958 469920 156014 469976
rect 154578 467200 154634 467256
rect 157430 468696 157486 468752
rect 160098 465976 160154 466032
rect 163594 478624 163650 478680
rect 161662 465840 161718 465896
rect 157338 460400 157394 460456
rect 153198 460128 153254 460184
rect 164330 460536 164386 460592
rect 167182 460808 167238 460864
rect 166998 460672 167054 460728
rect 170218 478760 170274 478816
rect 169850 466112 169906 466168
rect 168562 459312 168618 459368
rect 171598 474272 171654 474328
rect 171230 463120 171286 463176
rect 172702 470056 172758 470112
rect 172610 464344 172666 464400
rect 172518 459448 172574 459504
rect 171138 459176 171194 459232
rect 178314 461352 178370 461408
rect 179970 472640 180026 472696
rect 179510 461624 179566 461680
rect 185674 477944 185730 478000
rect 186318 463256 186374 463312
rect 187882 466248 187938 466304
rect 190918 460964 190974 461000
rect 190918 460944 190920 460964
rect 190920 460944 190972 460964
rect 190972 460944 190974 460964
rect 168378 459040 168434 459096
rect 164238 458904 164294 458960
rect 125690 458768 125746 458824
rect 158534 374584 158590 374640
rect 165986 374604 166042 374640
rect 165986 374584 165988 374604
rect 165988 374584 166040 374604
rect 166040 374584 166042 374604
rect 195886 374584 195942 374640
rect 105450 374448 105506 374504
rect 116030 374448 116086 374504
rect 140962 374448 141018 374504
rect 143538 374448 143594 374504
rect 156510 374468 156566 374504
rect 156510 374448 156512 374468
rect 156512 374448 156564 374468
rect 156564 374448 156566 374468
rect 139214 374040 139270 374096
rect 160926 374448 160982 374504
rect 163410 374448 163466 374504
rect 146206 374312 146262 374368
rect 148966 374312 149022 374368
rect 95054 373632 95110 373688
rect 96066 373632 96122 373688
rect 103518 373668 103520 373688
rect 103520 373668 103572 373688
rect 103572 373668 103574 373688
rect 103518 373632 103574 373668
rect 107842 373632 107898 373688
rect 113546 373652 113602 373688
rect 113546 373632 113548 373652
rect 113548 373632 113600 373652
rect 113600 373632 113602 373652
rect 93674 373360 93730 373416
rect 118330 373632 118386 373688
rect 121366 373632 121422 373688
rect 110418 373496 110474 373552
rect 124126 373532 124128 373552
rect 124128 373532 124180 373552
rect 124180 373532 124182 373552
rect 124126 373496 124182 373532
rect 125690 373516 125746 373552
rect 125690 373496 125692 373516
rect 125692 373496 125744 373516
rect 125744 373496 125746 373516
rect 128910 373516 128966 373552
rect 128910 373496 128912 373516
rect 128912 373496 128964 373516
rect 128964 373496 128966 373516
rect 131026 373496 131082 373552
rect 133694 373496 133750 373552
rect 136454 373496 136510 373552
rect 151726 373496 151782 373552
rect 154118 373496 154174 373552
rect 98274 373380 98330 373416
rect 98274 373360 98276 373380
rect 98276 373360 98328 373380
rect 98328 373360 98330 373380
rect 88338 373224 88394 373280
rect 95974 373224 96030 373280
rect 90178 373108 90234 373144
rect 90178 373088 90180 373108
rect 90180 373088 90232 373108
rect 90232 373088 90234 373108
rect 92386 373088 92442 373144
rect 62118 372680 62174 372736
rect 77206 372544 77262 372600
rect 85486 372544 85542 372600
rect 86590 372544 86646 372600
rect 88062 372544 88118 372600
rect 89350 372564 89406 372600
rect 89350 372544 89352 372564
rect 89352 372544 89404 372564
rect 89404 372544 89406 372564
rect 78494 372408 78550 372464
rect 79966 372408 80022 372464
rect 85118 372408 85174 372464
rect 77022 372136 77078 372192
rect 80518 372272 80574 372328
rect 81898 372272 81954 372328
rect 83830 371864 83886 371920
rect 90086 372544 90142 372600
rect 92202 372544 92258 372600
rect 93582 372544 93638 372600
rect 100850 373244 100906 373280
rect 100850 373224 100852 373244
rect 100852 373224 100904 373244
rect 100904 373224 100906 373244
rect 108854 372544 108910 372600
rect 114006 372544 114062 372600
rect 183190 372544 183246 372600
rect 102782 372408 102838 372464
rect 102046 372272 102102 372328
rect 97722 371592 97778 371648
rect 99286 371592 99342 371648
rect 100114 371592 100170 371648
rect 101034 371456 101090 371512
rect 104622 371864 104678 371920
rect 117962 372272 118018 372328
rect 117962 372000 118018 372056
rect 105910 371728 105966 371784
rect 104622 369688 104678 369744
rect 105910 369552 105966 369608
rect 182822 371456 182878 371512
rect 107566 371320 107622 371376
rect 197358 477672 197414 477728
rect 196898 465704 196954 465760
rect 179786 355272 179842 355328
rect 191378 355272 191434 355328
rect 178590 354748 178646 354784
rect 178590 354728 178592 354748
rect 178592 354728 178644 354748
rect 178644 354728 178646 354748
rect 110970 269864 111026 269920
rect 148506 269864 148562 269920
rect 83094 269592 83150 269648
rect 91282 269592 91338 269648
rect 93582 269592 93638 269648
rect 94502 269592 94558 269648
rect 133418 269728 133474 269784
rect 135902 269728 135958 269784
rect 138478 269728 138534 269784
rect 140870 269728 140926 269784
rect 76010 268776 76066 268832
rect 77114 268776 77170 268832
rect 66258 267008 66314 267064
rect 77298 267008 77354 267064
rect 78678 267008 78734 267064
rect 90730 268776 90786 268832
rect 143538 269592 143594 269648
rect 145930 269592 145986 269648
rect 95882 268776 95938 268832
rect 96066 268776 96122 268832
rect 98458 268776 98514 268832
rect 99378 268776 99434 268832
rect 100758 268776 100814 268832
rect 106370 268776 106426 268832
rect 85394 268096 85450 268152
rect 92386 268096 92442 268152
rect 84198 267688 84254 267744
rect 88338 267008 88394 267064
rect 85578 266328 85634 266384
rect 86958 266328 87014 266384
rect 88338 266328 88394 266384
rect 89718 266328 89774 266384
rect 103518 268096 103574 268152
rect 96986 267688 97042 267744
rect 97998 267724 98000 267744
rect 98000 267724 98052 267744
rect 98052 267724 98054 267744
rect 97998 267688 98054 267724
rect 102690 267688 102746 267744
rect 113546 268096 113602 268152
rect 128358 268096 128414 268152
rect 104898 267164 104954 267200
rect 104898 267144 104900 267164
rect 104900 267144 104952 267164
rect 104952 267144 104954 267164
rect 100758 267028 100814 267064
rect 100758 267008 100760 267028
rect 100760 267008 100812 267028
rect 100812 267008 100814 267028
rect 104898 266464 104954 266520
rect 92478 266328 92534 266384
rect 106278 266328 106334 266384
rect 111246 267724 111248 267744
rect 111248 267724 111300 267744
rect 111300 267724 111302 267744
rect 111246 267688 111302 267724
rect 112350 267688 112406 267744
rect 107658 267280 107714 267336
rect 119066 267688 119122 267744
rect 120078 267688 120134 267744
rect 125598 267688 125654 267744
rect 150990 267688 151046 267744
rect 158534 267708 158590 267744
rect 158534 267688 158536 267708
rect 158536 267688 158588 267708
rect 158588 267688 158590 267708
rect 163502 267688 163558 267744
rect 129738 267552 129794 267608
rect 155958 267552 156014 267608
rect 160926 267552 160982 267608
rect 115938 267416 115994 267472
rect 117318 267436 117374 267472
rect 117318 267416 117320 267436
rect 117320 267416 117372 267436
rect 117372 267416 117374 267436
rect 183282 267280 183338 267336
rect 109958 267008 110014 267064
rect 107658 266328 107714 266384
rect 183466 267008 183522 267064
rect 114374 266600 114430 266656
rect 117318 266600 117374 266656
rect 113730 266328 113786 266384
rect 179326 249872 179382 249928
rect 179786 249872 179842 249928
rect 190918 249872 190974 249928
rect 85854 249056 85910 249112
rect 96066 164872 96122 164928
rect 115754 164872 115810 164928
rect 84106 164600 84162 164656
rect 103518 164600 103574 164656
rect 105910 164600 105966 164656
rect 114374 164600 114430 164656
rect 138478 164736 138534 164792
rect 140870 164736 140926 164792
rect 143538 164736 143594 164792
rect 163318 164736 163374 164792
rect 76010 162696 76066 162752
rect 77298 162696 77354 162752
rect 78678 162696 78734 162752
rect 80058 162696 80114 162752
rect 81438 162696 81494 162752
rect 82818 162696 82874 162752
rect 75918 162152 75974 162208
rect 59358 140800 59414 140856
rect 98458 164192 98514 164248
rect 101034 164192 101090 164248
rect 108210 164192 108266 164248
rect 111154 163920 111210 163976
rect 99378 163104 99434 163160
rect 84198 162696 84254 162752
rect 85578 162696 85634 162752
rect 86958 162696 87014 162752
rect 88430 162696 88486 162752
rect 89810 162696 89866 162752
rect 90730 162696 90786 162752
rect 91190 162696 91246 162752
rect 92478 162696 92534 162752
rect 93858 162696 93914 162752
rect 95238 162696 95294 162752
rect 96618 162696 96674 162752
rect 97998 162696 98054 162752
rect 84106 161608 84162 161664
rect 84290 161608 84346 161664
rect 88338 162152 88394 162208
rect 90914 162424 90970 162480
rect 91098 162424 91154 162480
rect 90914 162152 90970 162208
rect 92478 145968 92534 146024
rect 100758 162696 100814 162752
rect 102138 162696 102194 162752
rect 103794 162696 103850 162752
rect 104898 162696 104954 162752
rect 106278 162696 106334 162752
rect 107658 162696 107714 162752
rect 110510 162696 110566 162752
rect 98642 145832 98698 145888
rect 100758 162016 100814 162072
rect 100022 145696 100078 145752
rect 106370 162424 106426 162480
rect 113454 163648 113510 163704
rect 118054 164600 118110 164656
rect 153382 164600 153438 164656
rect 122746 164192 122802 164248
rect 145930 164192 145986 164248
rect 148506 164192 148562 164248
rect 150898 164192 150954 164248
rect 110970 162696 111026 162752
rect 113178 162696 113234 162752
rect 115938 162696 115994 162752
rect 118330 162696 118386 162752
rect 118698 162696 118754 162752
rect 120722 162696 120778 162752
rect 112810 162172 112866 162208
rect 112810 162152 112812 162172
rect 112812 162152 112864 162172
rect 112864 162152 112866 162172
rect 116030 162424 116086 162480
rect 165894 164600 165950 164656
rect 128358 163104 128414 163160
rect 125874 162696 125930 162752
rect 130842 162696 130898 162752
rect 133418 162716 133474 162752
rect 133418 162696 133420 162716
rect 133420 162696 133472 162716
rect 133472 162696 133474 162716
rect 135994 162732 135996 162752
rect 135996 162732 136048 162752
rect 136048 162732 136050 162752
rect 135994 162696 136050 162732
rect 155958 162696 156014 162752
rect 183466 162696 183522 162752
rect 183190 162560 183246 162616
rect 198094 394576 198150 394632
rect 198278 391992 198334 392048
rect 198186 390632 198242 390688
rect 199014 454688 199070 454744
rect 199198 390768 199254 390824
rect 200118 478252 200120 478272
rect 200120 478252 200172 478272
rect 200172 478252 200174 478272
rect 200118 478216 200174 478252
rect 200670 477672 200726 477728
rect 199658 394032 199714 394088
rect 199566 390768 199622 390824
rect 199474 372680 199530 372736
rect 198738 349560 198794 349616
rect 199014 349560 199070 349616
rect 100758 145560 100814 145616
rect 191746 145424 191802 145480
rect 179050 144880 179106 144936
rect 179694 144880 179750 144936
rect 77114 59744 77170 59800
rect 83094 59744 83150 59800
rect 99470 59744 99526 59800
rect 113546 59744 113602 59800
rect 94502 59608 94558 59664
rect 95698 59608 95754 59664
rect 102782 59608 102838 59664
rect 103886 59608 103942 59664
rect 95698 59336 95754 59392
rect 95882 59336 95938 59392
rect 96986 59336 97042 59392
rect 101770 59336 101826 59392
rect 111154 59336 111210 59392
rect 115938 59336 115994 59392
rect 148506 59200 148562 59256
rect 150898 59200 150954 59256
rect 84198 57976 84254 58032
rect 76010 57840 76066 57896
rect 78218 57840 78274 57896
rect 79506 57840 79562 57896
rect 80058 57840 80114 57896
rect 81806 57840 81862 57896
rect 85394 57840 85450 57896
rect 86498 57840 86554 57896
rect 86958 57840 87014 57896
rect 88338 57840 88394 57896
rect 88706 57840 88762 57896
rect 89718 57840 89774 57896
rect 90730 57840 90786 57896
rect 91190 57840 91246 57896
rect 92110 57840 92166 57896
rect 92478 57840 92534 57896
rect 93674 57840 93730 57896
rect 98090 57840 98146 57896
rect 106370 57840 106426 57896
rect 107382 57840 107438 57896
rect 108026 57840 108082 57896
rect 112074 57840 112130 57896
rect 113178 57840 113234 57896
rect 123482 57840 123538 57896
rect 130842 57840 130898 57896
rect 133234 57840 133290 57896
rect 145562 57860 145618 57896
rect 145562 57840 145564 57860
rect 145564 57840 145616 57860
rect 145616 57840 145618 57860
rect 98642 57432 98698 57488
rect 98642 57024 98698 57080
rect 109038 57568 109094 57624
rect 153290 57840 153346 57896
rect 157430 57840 157486 57896
rect 183282 57860 183338 57896
rect 183282 57840 183284 57860
rect 183284 57840 183336 57860
rect 183336 57840 183338 57860
rect 113270 57568 113326 57624
rect 114558 57568 114614 57624
rect 116122 57568 116178 57624
rect 117318 57568 117374 57624
rect 118698 57568 118754 57624
rect 155958 57568 156014 57624
rect 153290 56344 153346 56400
rect 199014 289720 199070 289776
rect 198830 288360 198886 288416
rect 198830 287680 198886 287736
rect 198738 244160 198794 244216
rect 198922 283056 198978 283112
rect 198830 183504 198886 183560
rect 198830 182008 198886 182064
rect 198830 181328 198886 181384
rect 198738 179424 198794 179480
rect 199382 288360 199438 288416
rect 199658 388456 199714 388512
rect 199750 373768 199806 373824
rect 201498 477944 201554 478000
rect 199566 286320 199622 286376
rect 199106 284824 199162 284880
rect 199014 184320 199070 184376
rect 198922 178608 198978 178664
rect 198830 76336 198886 76392
rect 198738 74840 198794 74896
rect 199750 289720 199806 289776
rect 199658 283056 199714 283112
rect 199198 244160 199254 244216
rect 199106 179424 199162 179480
rect 201406 375264 201462 375320
rect 199382 183504 199438 183560
rect 199382 182688 199438 182744
rect 199290 182008 199346 182064
rect 199198 139168 199254 139224
rect 199014 79328 199070 79384
rect 199382 77696 199438 77752
rect 198922 73616 198978 73672
rect 202786 375264 202842 375320
rect 204350 478524 204352 478544
rect 204352 478524 204404 478544
rect 204404 478524 204406 478544
rect 204350 478488 204406 478524
rect 203706 267552 203762 267608
rect 205638 478660 205640 478680
rect 205640 478660 205692 478680
rect 205692 478660 205694 478680
rect 205638 478624 205694 478660
rect 205638 478352 205694 478408
rect 205546 456864 205602 456920
rect 205454 373904 205510 373960
rect 205454 373632 205510 373688
rect 206834 375264 206890 375320
rect 207754 459312 207810 459368
rect 208306 407768 208362 407824
rect 208214 265512 208270 265568
rect 183466 57740 183468 57760
rect 183468 57740 183520 57760
rect 183520 57740 183522 57760
rect 183466 57704 183522 57740
rect 208490 478488 208546 478544
rect 209042 465976 209098 466032
rect 208950 369144 209006 369200
rect 209410 266736 209466 266792
rect 212538 478080 212594 478136
rect 210054 371864 210110 371920
rect 210054 371592 210110 371648
rect 210330 371864 210386 371920
rect 210330 371456 210386 371512
rect 209594 265648 209650 265704
rect 209594 265512 209650 265568
rect 211066 375264 211122 375320
rect 210974 372680 211030 372736
rect 160098 57568 160154 57624
rect 165618 57568 165674 57624
rect 211618 372136 211674 372192
rect 211986 465840 212042 465896
rect 212446 382336 212502 382392
rect 212354 375264 212410 375320
rect 212262 371728 212318 371784
rect 212078 267416 212134 267472
rect 213918 478624 213974 478680
rect 212906 374584 212962 374640
rect 213182 459040 213238 459096
rect 213274 267280 213330 267336
rect 213642 371592 213698 371648
rect 213826 369144 213882 369200
rect 213458 266192 213514 266248
rect 213366 265104 213422 265160
rect 165618 55120 165674 55176
rect 160098 54984 160154 55040
rect 155958 54848 156014 54904
rect 118698 54712 118754 54768
rect 116122 54576 116178 54632
rect 214746 459176 214802 459232
rect 214930 466248 214986 466304
rect 215482 374312 215538 374368
rect 214930 264968 214986 265024
rect 214562 145832 214618 145888
rect 215206 369824 215262 369880
rect 215022 145424 215078 145480
rect 215390 369552 215446 369608
rect 215298 266328 215354 266384
rect 216954 477536 217010 477592
rect 215758 372272 215814 372328
rect 215666 369688 215722 369744
rect 215574 266056 215630 266112
rect 215574 265104 215630 265160
rect 215850 265648 215906 265704
rect 216678 408720 216734 408776
rect 216678 407788 216734 407824
rect 216678 407768 216680 407788
rect 216680 407768 216732 407788
rect 216732 407768 216734 407788
rect 216954 411304 217010 411360
rect 217046 409944 217102 410000
rect 216862 406000 216918 406056
rect 216678 384956 216680 384976
rect 216680 384956 216732 384976
rect 216732 384956 216734 384976
rect 216678 384920 216734 384956
rect 216678 383288 216734 383344
rect 216862 383016 216918 383072
rect 216770 375264 216826 375320
rect 216770 374856 216826 374912
rect 216310 267008 216366 267064
rect 215758 145968 215814 146024
rect 216218 146240 216274 146296
rect 216218 145968 216274 146024
rect 216494 266464 216550 266520
rect 216310 145696 216366 145752
rect 216954 374992 217010 375048
rect 217046 372680 217102 372736
rect 216954 303728 217010 303784
rect 216862 302776 216918 302832
rect 217046 301008 217102 301064
rect 216770 299376 216826 299432
rect 216678 279928 216734 279984
rect 216954 278316 217010 278352
rect 216954 278296 216956 278316
rect 216956 278296 217008 278316
rect 217008 278296 217010 278316
rect 216678 278024 216734 278080
rect 216954 268776 217010 268832
rect 216678 201864 216734 201920
rect 216770 201320 216826 201376
rect 216678 173304 216734 173360
rect 216678 96872 216734 96928
rect 216862 197376 216918 197432
rect 216770 95920 216826 95976
rect 217782 477672 217838 477728
rect 217782 410896 217838 410952
rect 217782 409944 217838 410000
rect 217966 411848 218022 411904
rect 217966 411304 218022 411360
rect 217690 404232 217746 404288
rect 217874 404912 217930 404968
rect 217874 404232 217930 404288
rect 217874 403144 217930 403200
rect 217874 375264 217930 375320
rect 217782 307672 217838 307728
rect 217782 306856 217838 306912
rect 217690 305904 217746 305960
rect 217414 303728 217470 303784
rect 217322 301008 217378 301064
rect 217230 299920 217286 299976
rect 217046 196016 217102 196072
rect 217046 173032 217102 173088
rect 217506 302776 217562 302832
rect 217414 198736 217470 198792
rect 217598 299376 217654 299432
rect 217598 298152 217654 298208
rect 217506 197784 217562 197840
rect 217506 197376 217562 197432
rect 217230 194928 217286 194984
rect 216862 92792 216918 92848
rect 216678 69944 216734 70000
rect 216678 68312 216734 68368
rect 218242 374176 218298 374232
rect 218610 372408 218666 372464
rect 218334 371592 218390 371648
rect 218150 371456 218206 371512
rect 217966 307672 218022 307728
rect 217966 267960 218022 268016
rect 218426 266872 218482 266928
rect 217874 265784 217930 265840
rect 217874 264968 217930 265024
rect 217782 201864 217838 201920
rect 217690 201320 217746 201376
rect 217690 200912 217746 200968
rect 217782 198736 217838 198792
rect 217690 196016 217746 196072
rect 217598 193160 217654 193216
rect 217230 89936 217286 89992
rect 217874 161084 217930 161120
rect 217874 161064 217876 161084
rect 217876 161064 217928 161084
rect 217928 161064 217930 161084
rect 217782 93744 217838 93800
rect 217690 91024 217746 91080
rect 217598 88168 217654 88224
rect 218334 163648 218390 163704
rect 217966 68312 218022 68368
rect 218886 458904 218942 458960
rect 219254 266872 219310 266928
rect 218702 60560 218758 60616
rect 219622 374040 219678 374096
rect 219438 371320 219494 371376
rect 219254 60560 219310 60616
rect 223118 477536 223174 477592
rect 222198 476720 222254 476776
rect 226154 478216 226210 478272
rect 230570 478488 230626 478544
rect 231490 478352 231546 478408
rect 232318 478080 232374 478136
rect 231858 475496 231914 475552
rect 233698 478216 233754 478272
rect 233238 474136 233294 474192
rect 234526 477944 234582 478000
rect 235906 478760 235962 478816
rect 235446 478624 235502 478680
rect 234066 471144 234122 471200
rect 230478 468424 230534 468480
rect 229098 465704 229154 465760
rect 223762 458904 223818 458960
rect 252742 474272 252798 474328
rect 255226 476856 255282 476912
rect 256146 472504 256202 472560
rect 263690 469784 263746 469840
rect 266358 461488 266414 461544
rect 278778 460128 278834 460184
rect 295522 462848 295578 462904
rect 296810 465840 296866 465896
rect 295430 460264 295486 460320
rect 338302 460980 338304 461000
rect 338304 460980 338356 461000
rect 338356 460980 338358 461000
rect 338302 460944 338358 460980
rect 339774 460964 339830 461000
rect 339774 460944 339776 460964
rect 339776 460944 339828 460964
rect 339828 460944 339830 460964
rect 350998 460964 351054 461000
rect 350998 460944 351000 460964
rect 351000 460944 351052 460964
rect 351052 460944 351054 460964
rect 223578 458768 223634 458824
rect 244738 374992 244794 375048
rect 270498 374992 270554 375048
rect 283010 374992 283066 375048
rect 311806 374992 311862 375048
rect 244278 374448 244334 374504
rect 220726 371728 220782 371784
rect 220726 371320 220782 371376
rect 222106 374176 222162 374232
rect 222014 374040 222070 374096
rect 235998 373088 236054 373144
rect 236090 372544 236146 372600
rect 238114 372544 238170 372600
rect 239310 372544 239366 372600
rect 240414 372544 240470 372600
rect 222106 372136 222162 372192
rect 222014 372000 222070 372056
rect 247590 374448 247646 374504
rect 253478 374448 253534 374504
rect 265254 374448 265310 374504
rect 270314 374176 270370 374232
rect 270222 374040 270278 374096
rect 242898 373224 242954 373280
rect 241518 372544 241574 372600
rect 245658 372544 245714 372600
rect 248418 372544 248474 372600
rect 258078 373768 258134 373824
rect 262862 373768 262918 373824
rect 253938 373108 253994 373144
rect 253938 373088 253940 373108
rect 253940 373088 253992 373108
rect 253992 373088 253994 373108
rect 255410 373088 255466 373144
rect 261298 373244 261354 373280
rect 261298 373224 261300 373244
rect 261300 373224 261352 373244
rect 261352 373224 261354 373244
rect 251178 372544 251234 372600
rect 256698 372544 256754 372600
rect 259458 372544 259514 372600
rect 259642 372544 259698 372600
rect 247038 371592 247094 371648
rect 249890 371592 249946 371648
rect 251178 371592 251234 371648
rect 249798 371340 249854 371376
rect 249798 371320 249800 371340
rect 249800 371320 249852 371340
rect 249852 371320 249854 371340
rect 263690 373516 263746 373552
rect 263690 373496 263692 373516
rect 263692 373496 263744 373516
rect 263744 373496 263746 373516
rect 269210 373380 269266 373416
rect 269210 373360 269212 373380
rect 269212 373360 269264 373380
rect 269264 373360 269266 373380
rect 270222 372136 270278 372192
rect 271970 373088 272026 373144
rect 300858 373088 300914 373144
rect 270314 372000 270370 372056
rect 273258 372564 273314 372600
rect 273258 372544 273260 372564
rect 273260 372544 273312 372564
rect 273312 372544 273314 372564
rect 276294 372408 276350 372464
rect 271970 371864 272026 371920
rect 278686 372272 278742 372328
rect 275374 371728 275430 371784
rect 262770 371456 262826 371512
rect 264978 371456 265034 371512
rect 252558 371320 252614 371376
rect 255318 371320 255374 371376
rect 258170 371320 258226 371376
rect 260838 371320 260894 371376
rect 263598 371320 263654 371376
rect 266358 371320 266414 371376
rect 267738 371320 267794 371376
rect 273350 371456 273406 371512
rect 276018 371320 276074 371376
rect 277766 371320 277822 371376
rect 280158 371320 280214 371376
rect 285678 371320 285734 371376
rect 287242 371320 287298 371376
rect 289818 371320 289874 371376
rect 292578 371320 292634 371376
rect 295338 371320 295394 371376
rect 298098 371320 298154 371376
rect 320914 374604 320970 374640
rect 320914 374584 320916 374604
rect 320916 374584 320968 374604
rect 320968 374584 320970 374604
rect 310518 372544 310574 372600
rect 313278 372564 313334 372600
rect 313278 372544 313280 372564
rect 313280 372544 313332 372564
rect 313332 372544 313334 372564
rect 304998 372408 305054 372464
rect 317418 371728 317474 371784
rect 302238 371320 302294 371376
rect 307758 371320 307814 371376
rect 325882 371592 325938 371648
rect 322938 371320 322994 371376
rect 343086 371320 343142 371376
rect 343454 371340 343510 371376
rect 343454 371320 343456 371340
rect 343456 371320 343508 371340
rect 343508 371320 343510 371340
rect 340050 355000 340106 355056
rect 351734 355000 351790 355056
rect 338118 354764 338120 354784
rect 338120 354764 338172 354784
rect 338172 354764 338174 354784
rect 338118 354728 338174 354764
rect 250718 269728 250774 269784
rect 283470 269592 283526 269648
rect 288254 269592 288310 269648
rect 291014 269592 291070 269648
rect 293406 269592 293462 269648
rect 305918 269592 305974 269648
rect 318430 269592 318486 269648
rect 243082 268776 243138 268832
rect 258078 268776 258134 268832
rect 261666 268776 261722 268832
rect 220818 267824 220874 267880
rect 295890 268796 295946 268832
rect 295890 268776 295892 268796
rect 295892 268776 295944 268796
rect 295944 268776 295946 268796
rect 298466 268812 298468 268832
rect 298468 268812 298520 268832
rect 298520 268812 298522 268832
rect 298466 268776 298522 268812
rect 300858 268776 300914 268832
rect 303434 268776 303490 268832
rect 323306 269048 323362 269104
rect 265162 268096 265218 268152
rect 275926 268096 275982 268152
rect 255318 267708 255374 267744
rect 255318 267688 255320 267708
rect 255320 267688 255372 267708
rect 255372 267688 255374 267708
rect 258262 267688 258318 267744
rect 260838 267688 260894 267744
rect 263598 267688 263654 267744
rect 264978 267688 265034 267744
rect 255318 267008 255374 267064
rect 247038 266872 247094 266928
rect 252558 266892 252614 266928
rect 252558 266872 252560 266892
rect 252560 266872 252612 266892
rect 252612 266872 252614 266892
rect 249798 266600 249854 266656
rect 244370 266464 244426 266520
rect 244278 266328 244334 266384
rect 245658 266328 245714 266384
rect 247038 266328 247094 266384
rect 248510 266328 248566 266384
rect 251270 266464 251326 266520
rect 259550 266464 259606 266520
rect 251178 266328 251234 266384
rect 252558 266328 252614 266384
rect 253938 266328 253994 266384
rect 256698 266328 256754 266384
rect 259458 266328 259514 266384
rect 262218 266348 262274 266384
rect 262218 266328 262220 266348
rect 262220 266328 262272 266348
rect 262272 266328 262274 266348
rect 263598 266328 263654 266384
rect 267830 267688 267886 267744
rect 270498 267688 270554 267744
rect 273258 267688 273314 267744
rect 273258 267028 273314 267064
rect 276018 267688 276074 267744
rect 277030 267688 277086 267744
rect 278134 267688 278190 267744
rect 280158 267688 280214 267744
rect 343454 267416 343510 267472
rect 279146 267164 279202 267200
rect 279146 267144 279148 267164
rect 279148 267144 279200 267164
rect 279200 267144 279202 267164
rect 273258 267008 273260 267028
rect 273260 267008 273312 267028
rect 273312 267008 273314 267028
rect 343454 267008 343510 267064
rect 285678 266872 285734 266928
rect 266358 266464 266414 266520
rect 266450 266328 266506 266384
rect 267738 266328 267794 266384
rect 269118 266328 269174 266384
rect 270498 266328 270554 266384
rect 273166 266328 273222 266384
rect 338486 249872 338542 249928
rect 340050 249872 340106 249928
rect 351734 249872 351790 249928
rect 261022 164736 261078 164792
rect 288254 164600 288310 164656
rect 305918 164600 305974 164656
rect 265898 164464 265954 164520
rect 298466 164192 298522 164248
rect 300858 164192 300914 164248
rect 303434 164192 303490 164248
rect 285954 163820 285956 163840
rect 285956 163820 286008 163840
rect 286008 163820 286010 163840
rect 285954 163784 286010 163820
rect 313370 164192 313426 164248
rect 235998 163104 236054 163160
rect 264978 163104 265034 163160
rect 276110 163104 276166 163160
rect 236090 162696 236146 162752
rect 263690 162832 263746 162888
rect 237378 162696 237434 162752
rect 240138 162696 240194 162752
rect 241518 162696 241574 162752
rect 242898 162696 242954 162752
rect 244370 162696 244426 162752
rect 245658 162696 245714 162752
rect 247038 162696 247094 162752
rect 248234 162696 248290 162752
rect 248418 162696 248474 162752
rect 249798 162696 249854 162752
rect 250626 162696 250682 162752
rect 251178 162696 251234 162752
rect 252558 162696 252614 162752
rect 253570 162696 253626 162752
rect 253938 162696 253994 162752
rect 255318 162696 255374 162752
rect 256146 162696 256202 162752
rect 256698 162696 256754 162752
rect 258354 162696 258410 162752
rect 259458 162696 259514 162752
rect 260838 162696 260894 162752
rect 262218 162696 262274 162752
rect 263598 162696 263654 162752
rect 238758 161472 238814 161528
rect 237378 145832 237434 145888
rect 244278 162016 244334 162072
rect 251270 162016 251326 162072
rect 258078 161472 258134 161528
rect 259550 162016 259606 162072
rect 268290 162832 268346 162888
rect 273442 162832 273498 162888
rect 266358 162696 266414 162752
rect 267554 162696 267610 162752
rect 267738 162696 267794 162752
rect 269118 162696 269174 162752
rect 270498 162696 270554 162752
rect 271878 162696 271934 162752
rect 273258 162696 273314 162752
rect 262218 146240 262274 146296
rect 269118 145696 269174 145752
rect 274822 162696 274878 162752
rect 276018 162696 276074 162752
rect 274546 162016 274602 162072
rect 280066 162696 280122 162752
rect 280802 162716 280858 162752
rect 280802 162696 280804 162716
rect 280804 162696 280856 162716
rect 280856 162696 280858 162716
rect 278042 161472 278098 161528
rect 278226 148960 278282 149016
rect 278226 148280 278282 148336
rect 276018 146376 276074 146432
rect 283746 162696 283802 162752
rect 293222 162732 293224 162752
rect 293224 162732 293276 162752
rect 293276 162732 293278 162752
rect 293222 162696 293278 162732
rect 320914 162696 320970 162752
rect 343454 162696 343510 162752
rect 343362 162560 343418 162616
rect 357438 477808 357494 477864
rect 270498 145560 270554 145616
rect 338486 144880 338542 144936
rect 340234 144880 340290 144936
rect 351642 144880 351698 144936
rect 237102 59744 237158 59800
rect 255870 59744 255926 59800
rect 256974 59744 257030 59800
rect 261758 59744 261814 59800
rect 263874 59744 263930 59800
rect 260654 59608 260710 59664
rect 262770 59472 262826 59528
rect 305918 59608 305974 59664
rect 318430 59608 318486 59664
rect 279238 59200 279294 59256
rect 290922 59200 290978 59256
rect 298466 59200 298522 59256
rect 313370 59200 313426 59256
rect 325882 59200 325938 59256
rect 259458 58656 259514 58712
rect 235998 57840 236054 57896
rect 237378 57840 237434 57896
rect 239218 57840 239274 57896
rect 240138 57840 240194 57896
rect 241610 57840 241666 57896
rect 242898 57840 242954 57896
rect 244370 57840 244426 57896
rect 245290 57840 245346 57896
rect 245658 57840 245714 57896
rect 247038 57840 247094 57896
rect 248602 57840 248658 57896
rect 249798 57840 249854 57896
rect 251178 57840 251234 57896
rect 251362 57840 251418 57896
rect 253386 57840 253442 57896
rect 253938 57840 253994 57896
rect 264978 57840 265034 57896
rect 265898 57840 265954 57896
rect 266358 57840 266414 57896
rect 268474 57840 268530 57896
rect 271234 57840 271290 57896
rect 271878 57840 271934 57896
rect 273258 57840 273314 57896
rect 275466 57840 275522 57896
rect 287610 57840 287666 57896
rect 293314 57840 293370 57896
rect 295890 57840 295946 57896
rect 300858 57840 300914 57896
rect 303434 57840 303490 57896
rect 308494 57840 308550 57896
rect 310978 57840 311034 57896
rect 315762 57860 315818 57896
rect 315762 57840 315764 57860
rect 315764 57840 315816 57860
rect 315816 57840 315818 57860
rect 266450 57568 266506 57624
rect 269118 57568 269174 57624
rect 273350 57568 273406 57624
rect 276018 57568 276074 57624
rect 320914 57840 320970 57896
rect 323306 57876 323308 57896
rect 323308 57876 323360 57896
rect 323360 57876 323362 57896
rect 323306 57840 323362 57876
rect 343178 57876 343180 57896
rect 343180 57876 343232 57896
rect 343232 57876 343234 57896
rect 343178 57840 343234 57876
rect 343454 57860 343510 57896
rect 357714 148960 357770 149016
rect 343454 57840 343456 57860
rect 343456 57840 343508 57860
rect 343508 57840 343510 57860
rect 358634 407768 358690 407824
rect 358542 269048 358598 269104
rect 358818 454688 358874 454744
rect 358818 373224 358874 373280
rect 359094 389272 359150 389328
rect 358910 349560 358966 349616
rect 360014 393760 360070 393816
rect 359922 392128 359978 392184
rect 359830 390768 359886 390824
rect 359094 289312 359150 289368
rect 359002 288360 359058 288416
rect 359002 283056 359058 283112
rect 358910 243752 358966 243808
rect 358910 183504 358966 183560
rect 358910 182688 358966 182744
rect 359278 286320 359334 286376
rect 359186 283056 359242 283112
rect 359094 184864 359150 184920
rect 359002 178608 359058 178664
rect 358910 78240 358966 78296
rect 360106 388048 360162 388104
rect 359554 288360 359610 288416
rect 359462 284824 359518 284880
rect 359370 243752 359426 243808
rect 359278 181328 359334 181384
rect 359094 79872 359150 79928
rect 359278 179424 359334 179480
rect 359186 76880 359242 76936
rect 359554 183504 359610 183560
rect 359462 179424 359518 179480
rect 359370 139304 359426 139360
rect 359278 75384 359334 75440
rect 359002 74024 359058 74080
rect 361118 266872 361174 266928
rect 276018 55120 276074 55176
rect 136454 3984 136510 4040
rect 132958 3848 133014 3904
rect 129370 3304 129426 3360
rect 147126 3712 147182 3768
rect 143538 3576 143594 3632
rect 140042 3168 140098 3224
rect 150622 3440 150678 3496
rect 370318 269320 370374 269376
rect 369306 164056 369362 164112
rect 371606 372680 371662 372736
rect 371606 265512 371662 265568
rect 371790 265104 371846 265160
rect 370962 148416 371018 148472
rect 373078 374040 373134 374096
rect 372526 145560 372582 145616
rect 373814 371728 373870 371784
rect 373814 265512 373870 265568
rect 374458 146240 374514 146296
rect 375838 266328 375894 266384
rect 375930 146240 375986 146296
rect 375930 145696 375986 145752
rect 376206 265104 376262 265160
rect 376114 162424 376170 162480
rect 377034 411884 377036 411904
rect 377036 411884 377088 411904
rect 377088 411884 377090 411904
rect 377034 411848 377090 411884
rect 376942 384956 376944 384976
rect 376944 384956 376996 384976
rect 376996 384956 376998 384976
rect 376942 384920 376998 384956
rect 376942 383288 376998 383344
rect 376850 383016 376906 383072
rect 376574 267144 376630 267200
rect 376574 266328 376630 266384
rect 376942 368464 376998 368520
rect 377218 410896 377274 410952
rect 377218 408720 377274 408776
rect 377126 407788 377182 407824
rect 377126 407768 377128 407788
rect 377128 407768 377180 407788
rect 377180 407768 377182 407788
rect 377218 406000 377274 406056
rect 377034 306856 377090 306912
rect 376850 278296 376906 278352
rect 376758 278024 376814 278080
rect 376298 161744 376354 161800
rect 377034 303592 377090 303648
rect 376942 202816 376998 202872
rect 377494 407768 377550 407824
rect 377310 304952 377366 305008
rect 377218 301008 377274 301064
rect 377126 264968 377182 265024
rect 376942 198736 376998 198792
rect 376850 174936 376906 174992
rect 376850 173304 376906 173360
rect 377770 410896 377826 410952
rect 377586 404948 377588 404968
rect 377588 404948 377640 404968
rect 377640 404948 377642 404968
rect 377586 404912 377642 404948
rect 377494 302776 377550 302832
rect 377310 200912 377366 200968
rect 377034 196016 377090 196072
rect 377218 196016 377274 196072
rect 376942 93744 376998 93800
rect 377218 193160 377274 193216
rect 377126 173032 377182 173088
rect 377034 91024 377090 91080
rect 377678 403144 377734 403200
rect 377862 408720 377918 408776
rect 429290 583276 429346 583332
rect 391938 485016 391994 485072
rect 377770 305904 377826 305960
rect 377770 304952 377826 305008
rect 377862 303592 377918 303648
rect 377586 299920 377642 299976
rect 377770 299920 377826 299976
rect 377678 264968 377734 265024
rect 377586 202816 377642 202872
rect 377586 201864 377642 201920
rect 377494 197784 377550 197840
rect 377310 95920 377366 95976
rect 377862 298152 377918 298208
rect 377770 194928 377826 194984
rect 377586 96872 377642 96928
rect 377494 92792 377550 92848
rect 377218 88168 377274 88224
rect 376942 69944 376998 70000
rect 376942 68332 376998 68368
rect 376942 68312 376944 68332
rect 376944 68312 376996 68332
rect 376996 68312 376998 68332
rect 377862 193160 377918 193216
rect 377770 89936 377826 89992
rect 378966 267552 379022 267608
rect 378874 162288 378930 162344
rect 430762 633392 430818 633448
rect 430670 632168 430726 632224
rect 580170 683848 580226 683904
rect 430946 626456 431002 626512
rect 430854 621968 430910 622024
rect 430762 616800 430818 616856
rect 430670 612448 430726 612504
rect 456798 619656 456854 619712
rect 456798 607416 456854 607472
rect 430578 607144 430634 607200
rect 430578 587968 430634 588024
rect 429474 553424 429530 553480
rect 429382 530848 429438 530904
rect 477130 619928 477186 619984
rect 488722 619928 488778 619984
rect 506754 619928 506810 619984
rect 457534 613536 457590 613592
rect 510710 616936 510766 616992
rect 580170 630828 580226 630864
rect 580170 630808 580172 630828
rect 580172 630808 580224 630828
rect 580224 630808 580226 630828
rect 511998 610816 512054 610872
rect 510618 604016 510674 604072
rect 457626 601296 457682 601352
rect 457534 588376 457590 588432
rect 457442 582256 457498 582312
rect 430670 578312 430726 578368
rect 457442 576136 457498 576192
rect 430762 572736 430818 572792
rect 430670 524864 430726 524920
rect 430854 567704 430910 567760
rect 430946 563080 431002 563136
rect 431038 549344 431094 549400
rect 431130 543904 431186 543960
rect 431222 539552 431278 539608
rect 431314 534384 431370 534440
rect 511998 597896 512054 597952
rect 457718 594496 457774 594552
rect 483018 482160 483074 482216
rect 506478 479712 506534 479768
rect 457534 479576 457590 479632
rect 512182 591776 512238 591832
rect 512090 585656 512146 585712
rect 511998 478352 512054 478408
rect 429290 475360 429346 475416
rect 512274 579536 512330 579592
rect 580170 577632 580226 577688
rect 513286 572756 513342 572792
rect 513286 572736 513288 572756
rect 513288 572736 513340 572756
rect 513340 572736 513342 572756
rect 512090 474000 512146 474056
rect 498198 460964 498254 461000
rect 498198 460944 498200 460964
rect 498200 460944 498252 460964
rect 498252 460944 498254 460964
rect 499854 460980 499856 461000
rect 499856 460980 499908 461000
rect 499908 460980 499910 461000
rect 499854 460944 499910 460980
rect 510894 460964 510950 461000
rect 510894 460944 510896 460964
rect 510896 460944 510948 460964
rect 510948 460944 510950 460964
rect 516598 454688 516654 454744
rect 407762 374992 407818 375048
rect 425058 374992 425114 375048
rect 440330 374992 440386 375048
rect 443090 374992 443146 375048
rect 404174 374720 404230 374776
rect 410706 374584 410762 374640
rect 433614 374448 433670 374504
rect 436006 374448 436062 374504
rect 438490 374448 438546 374504
rect 379058 162560 379114 162616
rect 379150 146240 379206 146296
rect 379426 265648 379482 265704
rect 379426 264968 379482 265024
rect 379426 250960 379482 251016
rect 379150 145832 379206 145888
rect 451002 374584 451058 374640
rect 416042 373788 416098 373824
rect 416042 373768 416044 373788
rect 416044 373768 416096 373788
rect 416096 373768 416098 373788
rect 421010 373768 421066 373824
rect 423034 373768 423090 373824
rect 426898 373804 426900 373824
rect 426900 373804 426952 373824
rect 426952 373804 426954 373824
rect 426898 373768 426954 373804
rect 430578 373768 430634 373824
rect 445850 373632 445906 373688
rect 455418 373652 455474 373688
rect 455418 373632 455420 373652
rect 455420 373632 455472 373652
rect 455472 373632 455474 373652
rect 447690 373516 447746 373552
rect 447690 373496 447692 373516
rect 447692 373496 447744 373516
rect 447744 373496 447746 373516
rect 458178 373496 458234 373552
rect 452842 373380 452898 373416
rect 452842 373360 452844 373380
rect 452844 373360 452896 373380
rect 452896 373360 452898 373380
rect 485778 373360 485834 373416
rect 408498 372544 408554 372600
rect 426438 372580 426440 372600
rect 426440 372580 426492 372600
rect 426492 372580 426494 372600
rect 426438 372544 426494 372580
rect 433338 372544 433394 372600
rect 437478 372564 437534 372600
rect 437478 372544 437480 372564
rect 437480 372544 437532 372564
rect 437532 372544 437534 372564
rect 470598 372272 470654 372328
rect 404358 372136 404414 372192
rect 396078 372020 396134 372056
rect 396078 372000 396080 372020
rect 396080 372000 396132 372020
rect 396132 372000 396134 372020
rect 397458 372000 397514 372056
rect 398838 372000 398894 372056
rect 400218 372000 400274 372056
rect 381082 371864 381138 371920
rect 409878 372000 409934 372056
rect 439870 371728 439926 371784
rect 401598 371592 401654 371648
rect 411258 371612 411314 371648
rect 411258 371592 411260 371612
rect 411260 371592 411312 371612
rect 411312 371592 411314 371612
rect 418342 371592 418398 371648
rect 423678 371592 423734 371648
rect 427818 371592 427874 371648
rect 407118 371476 407174 371512
rect 407118 371456 407120 371476
rect 407120 371456 407172 371476
rect 407172 371456 407174 371476
rect 411258 371456 411314 371512
rect 418250 371456 418306 371512
rect 396078 371320 396134 371376
rect 402978 371320 403034 371376
rect 405738 371320 405794 371376
rect 412638 371320 412694 371376
rect 413190 371320 413246 371376
rect 414018 371320 414074 371376
rect 415398 371320 415454 371376
rect 416778 371320 416834 371376
rect 418158 371320 418214 371376
rect 420918 371456 420974 371512
rect 419538 371320 419594 371376
rect 422298 371320 422354 371376
rect 425058 371320 425114 371376
rect 462318 371592 462374 371648
rect 465078 371592 465134 371648
rect 427910 371320 427966 371376
rect 431958 371320 432014 371376
rect 434718 371320 434774 371376
rect 436098 371320 436154 371376
rect 460938 371320 460994 371376
rect 467838 371320 467894 371376
rect 503166 372136 503222 372192
rect 503534 372136 503590 372192
rect 477498 371592 477554 371648
rect 473358 371320 473414 371376
rect 480258 371456 480314 371512
rect 483018 371320 483074 371376
rect 498842 355000 498898 355056
rect 500866 354864 500922 354920
rect 510894 354764 510896 354784
rect 510896 354764 510948 354784
rect 510948 354764 510950 354784
rect 510894 354728 510950 354764
rect 416042 269728 416098 269784
rect 425242 269728 425298 269784
rect 433338 269728 433394 269784
rect 434350 269728 434406 269784
rect 429750 269592 429806 269648
rect 422850 268912 422906 268968
rect 425978 268912 426034 268968
rect 416962 268776 417018 268832
rect 421010 268776 421066 268832
rect 398194 268096 398250 268152
rect 401690 268096 401746 268152
rect 388442 265104 388498 265160
rect 379978 264968 380034 265024
rect 379518 146240 379574 146296
rect 389178 264968 389234 265024
rect 396078 266348 396134 266384
rect 396078 266328 396080 266348
rect 396080 266328 396132 266348
rect 396132 266328 396134 266348
rect 398838 266328 398894 266384
rect 400218 266328 400274 266384
rect 436006 269592 436062 269648
rect 468482 269592 468538 269648
rect 470966 269592 471022 269648
rect 480902 269592 480958 269648
rect 430946 268912 431002 268968
rect 432234 268912 432290 268968
rect 475842 268912 475898 268968
rect 478418 268912 478474 268968
rect 483386 268912 483442 268968
rect 455786 268096 455842 268152
rect 402978 267688 403034 267744
rect 414386 267688 414442 267744
rect 415398 267688 415454 267744
rect 418158 267144 418214 267200
rect 409878 267008 409934 267064
rect 412914 267008 412970 267064
rect 408498 266600 408554 266656
rect 403162 266328 403218 266384
rect 404358 266328 404414 266384
rect 405738 266328 405794 266384
rect 407118 266328 407174 266384
rect 411350 266464 411406 266520
rect 418250 266464 418306 266520
rect 409878 266328 409934 266384
rect 411258 266328 411314 266384
rect 413006 266328 413062 266384
rect 418158 266328 418214 266384
rect 419538 266328 419594 266384
rect 420918 266328 420974 266384
rect 426438 266328 426494 266384
rect 428646 267688 428702 267744
rect 434718 267688 434774 267744
rect 449898 267688 449954 267744
rect 452658 267688 452714 267744
rect 442998 267416 443054 267472
rect 458178 267688 458234 267744
rect 460938 267708 460994 267744
rect 460938 267688 460940 267708
rect 460940 267688 460992 267708
rect 460992 267688 460994 267708
rect 503166 267416 503222 267472
rect 503534 267416 503590 267472
rect 440054 267280 440110 267336
rect 440238 267300 440294 267336
rect 440238 267280 440240 267300
rect 440240 267280 440292 267300
rect 440292 267280 440294 267300
rect 437478 267144 437534 267200
rect 433338 267028 433394 267064
rect 447138 267280 447194 267336
rect 445758 267164 445814 267200
rect 445758 267144 445760 267164
rect 445760 267144 445812 267164
rect 445812 267144 445814 267164
rect 433338 267008 433340 267028
rect 433340 267008 433392 267028
rect 433392 267008 433394 267028
rect 437478 266600 437534 266656
rect 436098 266328 436154 266384
rect 499026 249872 499082 249928
rect 500038 249872 500094 249928
rect 510894 249908 510896 249928
rect 510896 249908 510948 249928
rect 510948 249908 510950 249928
rect 510894 249872 510950 249908
rect 412546 164872 412602 164928
rect 401598 163104 401654 163160
rect 396078 162696 396134 162752
rect 397458 162696 397514 162752
rect 398838 162696 398894 162752
rect 400218 162696 400274 162752
rect 393962 162016 394018 162072
rect 380806 148416 380862 148472
rect 379978 146240 380034 146296
rect 396170 162152 396226 162208
rect 403070 162696 403126 162752
rect 404358 162696 404414 162752
rect 405738 162696 405794 162752
rect 407210 162696 407266 162752
rect 408314 162696 408370 162752
rect 408498 162696 408554 162752
rect 409878 162696 409934 162752
rect 410614 162696 410670 162752
rect 411350 162696 411406 162752
rect 402978 162152 403034 162208
rect 411258 162152 411314 162208
rect 425978 164736 426034 164792
rect 451002 164736 451058 164792
rect 423494 164600 423550 164656
rect 418434 164192 418490 164248
rect 421010 164192 421066 164248
rect 429750 164600 429806 164656
rect 436926 164600 436982 164656
rect 428186 164192 428242 164248
rect 416042 163104 416098 163160
rect 413558 162696 413614 162752
rect 414018 162696 414074 162752
rect 415490 162696 415546 162752
rect 412546 161472 412602 161528
rect 412730 161472 412786 161528
rect 415306 162016 415362 162072
rect 414018 146240 414074 146296
rect 430946 164192 431002 164248
rect 470966 164600 471022 164656
rect 480902 164600 480958 164656
rect 473450 164192 473506 164248
rect 475842 164192 475898 164248
rect 478418 164192 478474 164248
rect 483386 164192 483442 164248
rect 580170 511264 580226 511320
rect 518898 454144 518954 454200
rect 518990 393760 519046 393816
rect 519174 392128 519230 392184
rect 519082 388048 519138 388104
rect 518898 349152 518954 349208
rect 455786 163104 455842 163160
rect 416778 162696 416834 162752
rect 418158 162696 418214 162752
rect 419538 162696 419594 162752
rect 420918 162696 420974 162752
rect 422298 162696 422354 162752
rect 423678 162696 423734 162752
rect 425058 162696 425114 162752
rect 426438 162696 426494 162752
rect 429106 162696 429162 162752
rect 430578 162696 430634 162752
rect 431958 162696 432014 162752
rect 433338 162696 433394 162752
rect 435730 162696 435786 162752
rect 435914 162696 435970 162752
rect 437478 162696 437534 162752
rect 438490 162696 438546 162752
rect 438858 162696 438914 162752
rect 440882 162696 440938 162752
rect 443458 162696 443514 162752
rect 445850 162696 445906 162752
rect 448242 162696 448298 162752
rect 453394 162716 453450 162752
rect 453394 162696 453396 162716
rect 453396 162696 453448 162716
rect 453448 162696 453450 162716
rect 415490 145832 415546 145888
rect 418250 162172 418306 162208
rect 418250 162152 418252 162172
rect 418252 162152 418304 162172
rect 418304 162152 418306 162172
rect 416778 145696 416834 145752
rect 426530 162152 426586 162208
rect 434626 162152 434682 162208
rect 433522 162016 433578 162072
rect 458362 162696 458418 162752
rect 503258 162696 503314 162752
rect 503626 162560 503682 162616
rect 438858 148280 438914 148336
rect 422298 145560 422354 145616
rect 510618 145424 510674 145480
rect 498658 144880 498714 144936
rect 500222 144880 500278 144936
rect 396078 59744 396134 59800
rect 397090 59764 397146 59800
rect 397090 59744 397092 59764
rect 397092 59744 397144 59764
rect 397144 59744 397146 59764
rect 416962 59744 417018 59800
rect 418434 59744 418490 59800
rect 423954 59744 424010 59800
rect 403070 59608 403126 59664
rect 404174 59608 404230 59664
rect 412546 59608 412602 59664
rect 397458 57840 397514 57896
rect 399482 57840 399538 57896
rect 400218 57840 400274 57896
rect 401690 57840 401746 57896
rect 404358 57840 404414 57896
rect 405830 57840 405886 57896
rect 407210 57840 407266 57896
rect 408314 57840 408370 57896
rect 408682 57840 408738 57896
rect 409878 57840 409934 57896
rect 411350 57840 411406 57896
rect 411258 56888 411314 56944
rect 418158 59472 418214 59528
rect 419446 59608 419502 59664
rect 421746 59608 421802 59664
rect 423494 59608 423550 59664
rect 420642 59472 420698 59528
rect 503258 59608 503314 59664
rect 425242 59336 425298 59392
rect 425978 59336 426034 59392
rect 428186 59336 428242 59392
rect 465906 59336 465962 59392
rect 485962 59200 486018 59256
rect 414570 57840 414626 57896
rect 415490 57840 415546 57896
rect 416042 57840 416098 57896
rect 426438 57840 426494 57896
rect 427634 57840 427690 57896
rect 427818 57840 427874 57896
rect 429198 57840 429254 57896
rect 430578 57840 430634 57896
rect 431958 57840 432014 57896
rect 433430 57840 433486 57896
rect 435914 57840 435970 57896
rect 436098 57840 436154 57896
rect 438306 57840 438362 57896
rect 438490 57840 438546 57896
rect 438858 57840 438914 57896
rect 440882 57840 440938 57896
rect 443458 57860 443514 57896
rect 443458 57840 443460 57860
rect 443460 57840 443512 57860
rect 443512 57840 443514 57860
rect 412546 56888 412602 56944
rect 412638 56752 412694 56808
rect 427818 54984 427874 55040
rect 430946 57160 431002 57216
rect 433338 57160 433394 57216
rect 433522 57160 433578 57216
rect 435730 57160 435786 57216
rect 445850 57840 445906 57896
rect 451002 57840 451058 57896
rect 478418 57876 478420 57896
rect 478420 57876 478472 57896
rect 478472 57876 478474 57896
rect 478418 57840 478474 57876
rect 503350 57876 503352 57896
rect 503352 57876 503404 57896
rect 503404 57876 503406 57896
rect 503350 57840 503406 57876
rect 518990 289312 519046 289368
rect 518990 288360 519046 288416
rect 518990 287136 519046 287192
rect 518898 244160 518954 244216
rect 519266 390768 519322 390824
rect 519358 389272 519414 389328
rect 519174 288360 519230 288416
rect 580262 458088 580318 458144
rect 580262 404912 580318 404968
rect 519266 285776 519322 285832
rect 580446 378392 580502 378448
rect 580354 351872 580410 351928
rect 580262 325216 580318 325272
rect 519542 289312 519598 289368
rect 519358 284824 519414 284880
rect 519082 284144 519138 284200
rect 518990 182688 519046 182744
rect 519358 244160 519414 244216
rect 519266 184864 519322 184920
rect 519174 182688 519230 182744
rect 518990 179424 519046 179480
rect 518898 178744 518954 178800
rect 519634 285776 519690 285832
rect 519542 184864 519598 184920
rect 520186 284824 520242 284880
rect 580354 272176 580410 272232
rect 580262 232328 580318 232384
rect 580354 192480 580410 192536
rect 520186 182688 520242 182744
rect 519542 181328 519598 181384
rect 519450 179424 519506 179480
rect 519358 139304 519414 139360
rect 519266 79872 519322 79928
rect 519174 78240 519230 78296
rect 580262 152632 580318 152688
rect 520186 79872 520242 79928
rect 519542 76744 519598 76800
rect 518990 75384 519046 75440
rect 518898 74160 518954 74216
rect 438858 55120 438914 55176
rect 580446 112784 580502 112840
rect 580354 72936 580410 72992
rect 580262 33088 580318 33144
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect 280654 633388 280660 633452
rect 280724 633450 280730 633452
rect 430757 633450 430823 633453
rect 280724 633448 430823 633450
rect 280724 633392 430762 633448
rect 430818 633392 430823 633448
rect 280724 633390 430823 633392
rect 280724 633388 280730 633390
rect 430757 633387 430823 633390
rect 319529 632362 319595 632365
rect 392117 632362 392183 632365
rect 319529 632360 392183 632362
rect 319529 632304 319534 632360
rect 319590 632304 392122 632360
rect 392178 632304 392183 632360
rect 319529 632302 392183 632304
rect 319529 632299 319595 632302
rect 392117 632299 392183 632302
rect 281073 632226 281139 632229
rect 430665 632226 430731 632229
rect 281073 632224 430731 632226
rect -960 632090 480 632180
rect 281073 632168 281078 632224
rect 281134 632168 430670 632224
rect 430726 632168 430731 632224
rect 281073 632166 430731 632168
rect 281073 632163 281139 632166
rect 430665 632163 430731 632166
rect 3509 632090 3575 632093
rect -960 632088 3575 632090
rect -960 632032 3514 632088
rect 3570 632032 3575 632088
rect -960 632030 3575 632032
rect -960 631940 480 632030
rect 3509 632027 3575 632030
rect 42057 632090 42123 632093
rect 346393 632090 346459 632093
rect 42057 632088 346459 632090
rect 42057 632032 42062 632088
rect 42118 632032 346398 632088
rect 346454 632032 346459 632088
rect 42057 632030 346459 632032
rect 42057 632027 42123 632030
rect 346393 632027 346459 632030
rect 53046 630804 53052 630868
rect 53116 630866 53122 630868
rect 328085 630866 328151 630869
rect 53116 630864 328151 630866
rect 53116 630808 328090 630864
rect 328146 630808 328151 630864
rect 53116 630806 328151 630808
rect 53116 630804 53122 630806
rect 328085 630803 328151 630806
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 54334 630668 54340 630732
rect 54404 630730 54410 630732
rect 405365 630730 405431 630733
rect 54404 630728 405431 630730
rect 54404 630672 405370 630728
rect 405426 630672 405431 630728
rect 583520 630716 584960 630806
rect 54404 630670 405431 630672
rect 54404 630668 54410 630670
rect 405365 630667 405431 630670
rect 317781 629642 317847 629645
rect 320038 629642 320098 630224
rect 317781 629640 320098 629642
rect 317781 629584 317786 629640
rect 317842 629584 320098 629640
rect 317781 629582 320098 629584
rect 317781 629579 317847 629582
rect 430941 626514 431007 626517
rect 428782 626512 431007 626514
rect 428782 626456 430946 626512
rect 431002 626456 431007 626512
rect 428782 626454 431007 626456
rect 428782 626144 428842 626454
rect 430941 626451 431007 626454
rect 317597 625290 317663 625293
rect 320038 625290 320098 625464
rect 317597 625288 320098 625290
rect 317597 625232 317602 625288
rect 317658 625232 320098 625288
rect 317597 625230 320098 625232
rect 317597 625227 317663 625230
rect 430849 622026 430915 622029
rect 428782 622024 430915 622026
rect 428782 621968 430854 622024
rect 430910 621968 430915 622024
rect 428782 621966 430915 621968
rect 428782 621384 428842 621966
rect 430849 621963 430915 621966
rect 57697 620666 57763 620669
rect 137369 620666 137435 620669
rect 216673 620666 216739 620669
rect 57697 620664 60076 620666
rect 57697 620608 57702 620664
rect 57758 620608 60076 620664
rect 57697 620606 60076 620608
rect 137369 620664 140116 620666
rect 137369 620608 137374 620664
rect 137430 620608 140116 620664
rect 137369 620606 140116 620608
rect 216673 620664 220156 620666
rect 216673 620608 216678 620664
rect 216734 620608 220156 620664
rect 216673 620606 220156 620608
rect 57697 620603 57763 620606
rect 137369 620603 137435 620606
rect 216673 620603 216739 620606
rect 317965 620122 318031 620125
rect 320038 620122 320098 620704
rect 317965 620120 320098 620122
rect 317965 620064 317970 620120
rect 318026 620064 320098 620120
rect 317965 620062 320098 620064
rect 317965 620059 318031 620062
rect 122925 619986 122991 619989
rect 201585 619986 201651 619989
rect 281901 619986 281967 619989
rect 120796 619984 122991 619986
rect 120796 619928 122930 619984
rect 122986 619928 122991 619984
rect 120796 619926 122991 619928
rect 200836 619984 201651 619986
rect 200836 619928 201590 619984
rect 201646 619928 201651 619984
rect 200836 619926 201651 619928
rect 280876 619984 281967 619986
rect 280876 619928 281906 619984
rect 281962 619928 281967 619984
rect 280876 619926 281967 619928
rect 122925 619923 122991 619926
rect 201585 619923 201651 619926
rect 281901 619923 281967 619926
rect 476062 619924 476068 619988
rect 476132 619986 476138 619988
rect 477125 619986 477191 619989
rect 476132 619984 477191 619986
rect 476132 619928 477130 619984
rect 477186 619928 477191 619984
rect 476132 619926 477191 619928
rect 476132 619924 476138 619926
rect 477125 619923 477191 619926
rect 488574 619924 488580 619988
rect 488644 619986 488650 619988
rect 488717 619986 488783 619989
rect 488644 619984 488783 619986
rect 488644 619928 488722 619984
rect 488778 619928 488783 619984
rect 488644 619926 488783 619928
rect 488644 619924 488650 619926
rect 488717 619923 488783 619926
rect 506606 619924 506612 619988
rect 506676 619986 506682 619988
rect 506749 619986 506815 619989
rect 506676 619984 506815 619986
rect 506676 619928 506754 619984
rect 506810 619928 506815 619984
rect 506676 619926 506815 619928
rect 506676 619924 506682 619926
rect 506749 619923 506815 619926
rect 456793 619714 456859 619717
rect 456793 619712 460092 619714
rect 456793 619656 456798 619712
rect 456854 619656 460092 619712
rect 456793 619654 460092 619656
rect 456793 619651 456859 619654
rect -960 619020 480 619260
rect 59261 617810 59327 617813
rect 59494 617810 60076 617870
rect 139350 617818 140032 617878
rect 219390 617818 220064 617878
rect 139025 617810 139091 617813
rect 139350 617810 139410 617818
rect 59261 617808 59554 617810
rect 59261 617752 59266 617808
rect 59322 617752 59554 617808
rect 59261 617750 59554 617752
rect 139025 617808 139410 617810
rect 139025 617752 139030 617808
rect 139086 617752 139410 617808
rect 139025 617750 139410 617752
rect 216673 617810 216739 617813
rect 219390 617810 219450 617818
rect 216673 617808 219450 617810
rect 216673 617752 216678 617808
rect 216734 617752 219450 617808
rect 216673 617750 219450 617752
rect 59261 617747 59327 617750
rect 139025 617747 139091 617750
rect 216673 617747 216739 617750
rect 583520 617388 584960 617628
rect 123109 617266 123175 617269
rect 202873 617266 202939 617269
rect 120796 617264 123175 617266
rect 120796 617208 123114 617264
rect 123170 617208 123175 617264
rect 120796 617206 123175 617208
rect 200836 617264 202939 617266
rect 200836 617208 202878 617264
rect 202934 617208 202939 617264
rect 200836 617206 202939 617208
rect 123109 617203 123175 617206
rect 202873 617203 202939 617206
rect 280846 616997 280906 617236
rect 280846 616992 280955 616997
rect 510705 616994 510771 616997
rect 280846 616936 280894 616992
rect 280950 616936 280955 616992
rect 280846 616934 280955 616936
rect 509956 616992 510771 616994
rect 509956 616936 510710 616992
rect 510766 616936 510771 616992
rect 509956 616934 510771 616936
rect 280889 616931 280955 616934
rect 510705 616931 510771 616934
rect 430757 616858 430823 616861
rect 428782 616856 430823 616858
rect 428782 616800 430762 616856
rect 430818 616800 430823 616856
rect 428782 616798 430823 616800
rect 428782 616624 428842 616798
rect 430757 616795 430823 616798
rect 317965 615634 318031 615637
rect 320038 615634 320098 615944
rect 317965 615632 320098 615634
rect 317965 615576 317970 615632
rect 318026 615576 320098 615632
rect 317965 615574 320098 615576
rect 317965 615571 318031 615574
rect 57513 614410 57579 614413
rect 59494 614410 60076 614470
rect 139350 614418 140032 614478
rect 219390 614418 220064 614478
rect 139209 614410 139275 614413
rect 139350 614410 139410 614418
rect 57513 614408 59554 614410
rect 57513 614352 57518 614408
rect 57574 614352 59554 614408
rect 57513 614350 59554 614352
rect 139209 614408 139410 614410
rect 139209 614352 139214 614408
rect 139270 614352 139410 614408
rect 139209 614350 139410 614352
rect 217685 614410 217751 614413
rect 219390 614410 219450 614418
rect 217685 614408 219450 614410
rect 217685 614352 217690 614408
rect 217746 614352 219450 614408
rect 217685 614350 219450 614352
rect 57513 614347 57579 614350
rect 139209 614347 139275 614350
rect 217685 614347 217751 614350
rect 121729 613866 121795 613869
rect 201769 613866 201835 613869
rect 282913 613866 282979 613869
rect 120796 613864 121795 613866
rect 120796 613808 121734 613864
rect 121790 613808 121795 613864
rect 120796 613806 121795 613808
rect 200836 613864 201835 613866
rect 200836 613808 201774 613864
rect 201830 613808 201835 613864
rect 200836 613806 201835 613808
rect 280876 613864 282979 613866
rect 280876 613808 282918 613864
rect 282974 613808 282979 613864
rect 280876 613806 282979 613808
rect 121729 613803 121795 613806
rect 201769 613803 201835 613806
rect 282913 613803 282979 613806
rect 457529 613594 457595 613597
rect 457529 613592 460092 613594
rect 457529 613536 457534 613592
rect 457590 613536 460092 613592
rect 457529 613534 460092 613536
rect 457529 613531 457595 613534
rect 430665 612506 430731 612509
rect 428782 612504 430731 612506
rect 428782 612448 430670 612504
rect 430726 612448 430731 612504
rect 428782 612446 430731 612448
rect 428782 611864 428842 612446
rect 430665 612443 430731 612446
rect 59077 611690 59143 611693
rect 59494 611690 60076 611750
rect 139350 611698 140032 611758
rect 219390 611698 220064 611758
rect 137645 611690 137711 611693
rect 139350 611690 139410 611698
rect 59077 611688 59554 611690
rect 59077 611632 59082 611688
rect 59138 611632 59554 611688
rect 59077 611630 59554 611632
rect 137645 611688 139410 611690
rect 137645 611632 137650 611688
rect 137706 611632 139410 611688
rect 137645 611630 139410 611632
rect 215937 611690 216003 611693
rect 219390 611690 219450 611698
rect 215937 611688 219450 611690
rect 215937 611632 215942 611688
rect 215998 611632 219450 611688
rect 215937 611630 219450 611632
rect 59077 611627 59143 611630
rect 137645 611627 137711 611630
rect 215937 611627 216003 611630
rect 121913 611146 121979 611149
rect 203057 611146 203123 611149
rect 281625 611146 281691 611149
rect 120796 611144 121979 611146
rect 120796 611088 121918 611144
rect 121974 611088 121979 611144
rect 120796 611086 121979 611088
rect 200836 611144 203123 611146
rect 200836 611088 203062 611144
rect 203118 611088 203123 611144
rect 200836 611086 203123 611088
rect 280876 611144 281691 611146
rect 280876 611088 281630 611144
rect 281686 611088 281691 611144
rect 280876 611086 281691 611088
rect 121913 611083 121979 611086
rect 203057 611083 203123 611086
rect 281625 611083 281691 611086
rect 317873 610602 317939 610605
rect 320038 610602 320098 611184
rect 511993 610874 512059 610877
rect 509956 610872 512059 610874
rect 509956 610816 511998 610872
rect 512054 610816 512059 610872
rect 509956 610814 512059 610816
rect 511993 610811 512059 610814
rect 317873 610600 320098 610602
rect 317873 610544 317878 610600
rect 317934 610544 320098 610600
rect 317873 610542 320098 610544
rect 317873 610539 317939 610542
rect 58893 608290 58959 608293
rect 59494 608290 60076 608350
rect 139350 608298 140032 608358
rect 219390 608298 220064 608358
rect 136725 608290 136791 608293
rect 139350 608290 139410 608298
rect 58893 608288 59554 608290
rect 58893 608232 58898 608288
rect 58954 608232 59554 608288
rect 58893 608230 59554 608232
rect 136725 608288 139410 608290
rect 136725 608232 136730 608288
rect 136786 608232 139410 608288
rect 136725 608230 139410 608232
rect 216673 608290 216739 608293
rect 219390 608290 219450 608298
rect 216673 608288 219450 608290
rect 216673 608232 216678 608288
rect 216734 608232 219450 608288
rect 216673 608230 219450 608232
rect 58893 608227 58959 608230
rect 136725 608227 136791 608230
rect 216673 608227 216739 608230
rect 123017 607746 123083 607749
rect 202965 607746 203031 607749
rect 283005 607746 283071 607749
rect 120796 607744 123083 607746
rect 120796 607688 123022 607744
rect 123078 607688 123083 607744
rect 120796 607686 123083 607688
rect 200836 607744 203031 607746
rect 200836 607688 202970 607744
rect 203026 607688 203031 607744
rect 200836 607686 203031 607688
rect 280876 607744 283071 607746
rect 280876 607688 283010 607744
rect 283066 607688 283071 607744
rect 280876 607686 283071 607688
rect 123017 607683 123083 607686
rect 202965 607683 203031 607686
rect 283005 607683 283071 607686
rect 456793 607474 456859 607477
rect 456793 607472 460092 607474
rect 456793 607416 456798 607472
rect 456854 607416 460092 607472
rect 456793 607414 460092 607416
rect 456793 607411 456859 607414
rect 430573 607202 430639 607205
rect 428782 607200 430639 607202
rect 428782 607144 430578 607200
rect 430634 607144 430639 607200
rect 428782 607142 430639 607144
rect 428782 607104 428842 607142
rect 430573 607139 430639 607142
rect -960 605964 480 606204
rect 317965 606114 318031 606117
rect 320038 606114 320098 606424
rect 317965 606112 320098 606114
rect 317965 606056 317970 606112
rect 318026 606056 320098 606112
rect 317965 606054 320098 606056
rect 317965 606051 318031 606054
rect 59169 605570 59235 605573
rect 59494 605570 60076 605630
rect 139350 605578 140032 605638
rect 219390 605578 220064 605638
rect 138841 605570 138907 605573
rect 139350 605570 139410 605578
rect 59169 605568 59554 605570
rect 59169 605512 59174 605568
rect 59230 605512 59554 605568
rect 59169 605510 59554 605512
rect 138841 605568 139410 605570
rect 138841 605512 138846 605568
rect 138902 605512 139410 605568
rect 138841 605510 139410 605512
rect 219249 605570 219315 605573
rect 219390 605570 219450 605578
rect 219249 605568 219450 605570
rect 219249 605512 219254 605568
rect 219310 605512 219450 605568
rect 219249 605510 219450 605512
rect 59169 605507 59235 605510
rect 138841 605507 138907 605510
rect 219249 605507 219315 605510
rect 123201 605026 123267 605029
rect 201861 605026 201927 605029
rect 283189 605026 283255 605029
rect 120796 605024 123267 605026
rect 120796 604968 123206 605024
rect 123262 604968 123267 605024
rect 120796 604966 123267 604968
rect 200836 605024 201927 605026
rect 200836 604968 201866 605024
rect 201922 604968 201927 605024
rect 200836 604966 201927 604968
rect 280876 605024 283255 605026
rect 280876 604968 283194 605024
rect 283250 604968 283255 605024
rect 280876 604966 283255 604968
rect 123201 604963 123267 604966
rect 201861 604963 201927 604966
rect 283189 604963 283255 604966
rect 510613 604074 510679 604077
rect 509956 604072 510679 604074
rect 509956 604016 510618 604072
rect 510674 604016 510679 604072
rect 583520 604060 584960 604300
rect 509956 604014 510679 604016
rect 510613 604011 510679 604014
rect 58985 602170 59051 602173
rect 59494 602170 60076 602230
rect 139350 602178 140032 602238
rect 219390 602178 220064 602238
rect 138933 602170 138999 602173
rect 139350 602170 139410 602178
rect 58985 602168 59554 602170
rect 58985 602112 58990 602168
rect 59046 602112 59554 602168
rect 58985 602110 59554 602112
rect 138933 602168 139410 602170
rect 138933 602112 138938 602168
rect 138994 602112 139410 602168
rect 138933 602110 139410 602112
rect 217225 602170 217291 602173
rect 219390 602170 219450 602178
rect 217225 602168 219450 602170
rect 217225 602112 217230 602168
rect 217286 602112 219450 602168
rect 217225 602110 219450 602112
rect 58985 602107 59051 602110
rect 138933 602107 138999 602110
rect 217225 602107 217291 602110
rect 428782 601762 428842 602344
rect 430614 601762 430620 601764
rect 428782 601702 430620 601762
rect 430614 601700 430620 601702
rect 430684 601700 430690 601764
rect 121821 601626 121887 601629
rect 203149 601626 203215 601629
rect 283097 601626 283163 601629
rect 120796 601624 121887 601626
rect 120796 601568 121826 601624
rect 121882 601568 121887 601624
rect 120796 601566 121887 601568
rect 200836 601624 203215 601626
rect 200836 601568 203154 601624
rect 203210 601568 203215 601624
rect 200836 601566 203215 601568
rect 280876 601624 283163 601626
rect 280876 601568 283102 601624
rect 283158 601568 283163 601624
rect 280876 601566 283163 601568
rect 121821 601563 121887 601566
rect 203149 601563 203215 601566
rect 283097 601563 283163 601566
rect 317597 601082 317663 601085
rect 320038 601082 320098 601664
rect 457621 601354 457687 601357
rect 457621 601352 460092 601354
rect 457621 601296 457626 601352
rect 457682 601296 460092 601352
rect 457621 601294 460092 601296
rect 457621 601291 457687 601294
rect 317597 601080 320098 601082
rect 317597 601024 317602 601080
rect 317658 601024 320098 601080
rect 317597 601022 320098 601024
rect 317597 601019 317663 601022
rect 57881 599586 57947 599589
rect 137829 599586 137895 599589
rect 217777 599586 217843 599589
rect 57881 599584 59554 599586
rect 57881 599528 57886 599584
rect 57942 599566 59554 599584
rect 137829 599584 139594 599586
rect 57942 599528 60076 599566
rect 57881 599526 60076 599528
rect 57881 599523 57947 599526
rect 59494 599506 60076 599526
rect 137829 599528 137834 599584
rect 137890 599566 139594 599584
rect 217777 599584 219818 599586
rect 137890 599528 140116 599566
rect 137829 599526 140116 599528
rect 137829 599523 137895 599526
rect 139534 599506 140116 599526
rect 217777 599528 217782 599584
rect 217838 599566 219818 599584
rect 217838 599528 220156 599566
rect 217777 599526 220156 599528
rect 217777 599523 217843 599526
rect 219758 599506 220156 599526
rect 283281 598906 283347 598909
rect 280876 598904 283347 598906
rect 120766 598365 120826 598876
rect 200806 598365 200866 598876
rect 280876 598848 283286 598904
rect 283342 598848 283347 598904
rect 280876 598846 283347 598848
rect 283281 598843 283347 598846
rect 120766 598360 120875 598365
rect 120766 598304 120814 598360
rect 120870 598304 120875 598360
rect 120766 598302 120875 598304
rect 120809 598299 120875 598302
rect 200757 598360 200866 598365
rect 200757 598304 200762 598360
rect 200818 598304 200866 598360
rect 200757 598302 200866 598304
rect 200757 598299 200823 598302
rect 511993 597954 512059 597957
rect 509956 597952 512059 597954
rect 509956 597896 511998 597952
rect 512054 597896 512059 597952
rect 509956 597894 512059 597896
rect 511993 597891 512059 597894
rect 430798 597682 430804 597684
rect 428782 597622 430804 597682
rect 428782 597584 428842 597622
rect 430798 597620 430804 597622
rect 430868 597620 430874 597684
rect 317597 596458 317663 596461
rect 320038 596458 320098 596904
rect 317597 596456 320098 596458
rect 317597 596400 317602 596456
rect 317658 596400 320098 596456
rect 317597 596398 320098 596400
rect 317597 596395 317663 596398
rect 137921 596186 137987 596189
rect 218697 596186 218763 596189
rect 137921 596184 139594 596186
rect 137921 596128 137926 596184
rect 137982 596160 139594 596184
rect 218697 596184 219818 596186
rect 137982 596128 140116 596160
rect 137921 596126 140116 596128
rect 137921 596123 137987 596126
rect 57881 596050 57947 596053
rect 59494 596050 60076 596110
rect 139534 596100 140116 596126
rect 218697 596128 218702 596184
rect 218758 596166 219818 596184
rect 218758 596128 220156 596166
rect 218697 596126 220156 596128
rect 218697 596123 218763 596126
rect 219758 596106 220156 596126
rect 57881 596048 59554 596050
rect 57881 595992 57886 596048
rect 57942 595992 59554 596048
rect 57881 595990 59554 595992
rect 57881 595987 57947 595990
rect 123385 595506 123451 595509
rect 203057 595506 203123 595509
rect 120796 595504 123451 595506
rect 120796 595448 123390 595504
rect 123446 595448 123451 595504
rect 120796 595446 123451 595448
rect 200836 595504 203123 595506
rect 200836 595448 203062 595504
rect 203118 595448 203123 595504
rect 200836 595446 203123 595448
rect 123385 595443 123451 595446
rect 203057 595443 203123 595446
rect 280846 594962 280906 595476
rect 280981 594962 281047 594965
rect 280846 594960 281047 594962
rect 280846 594904 280986 594960
rect 281042 594904 281047 594960
rect 280846 594902 281047 594904
rect 280981 594899 281047 594902
rect 137277 594826 137343 594829
rect 137921 594826 137987 594829
rect 137277 594824 137987 594826
rect 137277 594768 137282 594824
rect 137338 594768 137926 594824
rect 137982 594768 137987 594824
rect 137277 594766 137987 594768
rect 137277 594763 137343 594766
rect 137921 594763 137987 594766
rect 457713 594554 457779 594557
rect 457713 594552 460092 594554
rect 457713 594496 457718 594552
rect 457774 594496 460092 594552
rect 457713 594494 460092 594496
rect 457713 594491 457779 594494
rect 57605 593466 57671 593469
rect 137921 593466 137987 593469
rect 216673 593466 216739 593469
rect 57605 593464 59554 593466
rect 57605 593408 57610 593464
rect 57666 593446 59554 593464
rect 137921 593464 139594 593466
rect 57666 593408 60076 593446
rect 57605 593406 60076 593408
rect 57605 593403 57671 593406
rect 59494 593386 60076 593406
rect 137921 593408 137926 593464
rect 137982 593446 139594 593464
rect 216673 593464 219818 593466
rect 137982 593408 140116 593446
rect 137921 593406 140116 593408
rect 137921 593403 137987 593406
rect 139534 593386 140116 593406
rect 216673 593408 216678 593464
rect 216734 593446 219818 593464
rect 216734 593408 220156 593446
rect 216673 593406 220156 593408
rect 216673 593403 216739 593406
rect 219758 593386 220156 593406
rect -960 592908 480 593148
rect 123293 592786 123359 592789
rect 201953 592786 202019 592789
rect 281165 592786 281231 592789
rect 120796 592784 123359 592786
rect 120796 592728 123298 592784
rect 123354 592728 123359 592784
rect 120796 592726 123359 592728
rect 200836 592784 202019 592786
rect 200836 592728 201958 592784
rect 202014 592728 202019 592784
rect 200836 592726 202019 592728
rect 280876 592784 281231 592786
rect 280876 592728 281170 592784
rect 281226 592728 281231 592784
rect 280876 592726 281231 592728
rect 123293 592723 123359 592726
rect 201953 592723 202019 592726
rect 281165 592723 281231 592726
rect 318793 592786 318859 592789
rect 318793 592784 320098 592786
rect 318793 592728 318798 592784
rect 318854 592728 320098 592784
rect 318793 592726 320098 592728
rect 318793 592723 318859 592726
rect 320038 592144 320098 592726
rect 428782 592242 428842 592824
rect 430982 592242 430988 592244
rect 428782 592182 430988 592242
rect 430982 592180 430988 592182
rect 431052 592180 431058 592244
rect 512177 591834 512243 591837
rect 509956 591832 512243 591834
rect 509956 591776 512182 591832
rect 512238 591776 512243 591832
rect 509956 591774 512243 591776
rect 512177 591771 512243 591774
rect 583520 590868 584960 591108
rect 57421 589930 57487 589933
rect 59494 589930 60076 589990
rect 139350 589938 140032 589998
rect 219390 589938 220064 589998
rect 136725 589930 136791 589933
rect 139350 589930 139410 589938
rect 57421 589928 59554 589930
rect 57421 589872 57426 589928
rect 57482 589872 59554 589928
rect 57421 589870 59554 589872
rect 136725 589928 139410 589930
rect 136725 589872 136730 589928
rect 136786 589872 139410 589928
rect 136725 589870 139410 589872
rect 216673 589930 216739 589933
rect 219390 589930 219450 589938
rect 216673 589928 219450 589930
rect 216673 589872 216678 589928
rect 216734 589872 219450 589928
rect 216673 589870 219450 589872
rect 57421 589867 57487 589870
rect 136725 589867 136791 589870
rect 216673 589867 216739 589870
rect 124121 589386 124187 589389
rect 203241 589386 203307 589389
rect 283649 589386 283715 589389
rect 120796 589384 124187 589386
rect 120796 589328 124126 589384
rect 124182 589328 124187 589384
rect 120796 589326 124187 589328
rect 200836 589384 203307 589386
rect 200836 589328 203246 589384
rect 203302 589328 203307 589384
rect 200836 589326 203307 589328
rect 280876 589384 283715 589386
rect 280876 589328 283654 589384
rect 283710 589328 283715 589384
rect 280876 589326 283715 589328
rect 124121 589323 124187 589326
rect 203241 589323 203307 589326
rect 283649 589323 283715 589326
rect 457529 588434 457595 588437
rect 457529 588432 460092 588434
rect 457529 588376 457534 588432
rect 457590 588376 460092 588432
rect 457529 588374 460092 588376
rect 457529 588371 457595 588374
rect 428782 588026 428842 588064
rect 430573 588026 430639 588029
rect 428782 588024 430639 588026
rect 428782 587968 430578 588024
rect 430634 587968 430639 588024
rect 428782 587966 430639 587968
rect 430573 587963 430639 587966
rect 59494 587210 60076 587270
rect 139350 587218 140032 587278
rect 219390 587218 220064 587278
rect 138749 587210 138815 587213
rect 139350 587210 139410 587218
rect 57329 586394 57395 586397
rect 59494 586394 59554 587210
rect 138749 587208 139410 587210
rect 138749 587152 138754 587208
rect 138810 587152 139410 587208
rect 138749 587150 139410 587152
rect 216673 587210 216739 587213
rect 219390 587210 219450 587218
rect 216673 587208 219450 587210
rect 216673 587152 216678 587208
rect 216734 587152 219450 587208
rect 216673 587150 219450 587152
rect 138749 587147 138815 587150
rect 216673 587147 216739 587150
rect 122189 586666 122255 586669
rect 202137 586666 202203 586669
rect 281717 586666 281783 586669
rect 120796 586664 122255 586666
rect 120796 586608 122194 586664
rect 122250 586608 122255 586664
rect 120796 586606 122255 586608
rect 200836 586664 202203 586666
rect 200836 586608 202142 586664
rect 202198 586608 202203 586664
rect 200836 586606 202203 586608
rect 280876 586664 281783 586666
rect 280876 586608 281722 586664
rect 281778 586608 281783 586664
rect 280876 586606 281783 586608
rect 122189 586603 122255 586606
rect 202137 586603 202203 586606
rect 281717 586603 281783 586606
rect 317413 586530 317479 586533
rect 317413 586528 317522 586530
rect 317413 586472 317418 586528
rect 317474 586472 317522 586528
rect 317413 586467 317522 586472
rect 57329 586392 59554 586394
rect 57329 586336 57334 586392
rect 57390 586336 59554 586392
rect 57329 586334 59554 586336
rect 317462 586394 317522 586467
rect 320038 586394 320098 587384
rect 317462 586334 320098 586394
rect 57329 586331 57395 586334
rect 512085 585714 512151 585717
rect 509956 585712 512151 585714
rect 509956 585656 512090 585712
rect 512146 585656 512151 585712
rect 509956 585654 512151 585656
rect 512085 585651 512151 585654
rect 59494 583810 60076 583870
rect 139350 583818 140032 583878
rect 219390 583818 220064 583878
rect 137829 583810 137895 583813
rect 139350 583810 139410 583818
rect 57470 583750 59554 583810
rect 137829 583808 139410 583810
rect 137829 583752 137834 583808
rect 137890 583752 139410 583808
rect 137829 583750 139410 583752
rect 217409 583810 217475 583813
rect 219390 583810 219450 583818
rect 217409 583808 219450 583810
rect 217409 583752 217414 583808
rect 217470 583752 219450 583808
rect 217409 583750 219450 583752
rect 57470 583677 57530 583750
rect 137829 583747 137895 583750
rect 217409 583747 217475 583750
rect 57470 583672 57579 583677
rect 57470 583616 57518 583672
rect 57574 583616 57579 583672
rect 57470 583614 57579 583616
rect 57513 583611 57579 583614
rect 429285 583334 429351 583337
rect 428812 583332 429351 583334
rect 428812 583276 429290 583332
rect 429346 583276 429351 583332
rect 428812 583274 429351 583276
rect 429285 583271 429351 583274
rect 122097 583266 122163 583269
rect 202045 583266 202111 583269
rect 283373 583266 283439 583269
rect 120796 583264 122163 583266
rect 120796 583208 122102 583264
rect 122158 583208 122163 583264
rect 120796 583206 122163 583208
rect 200836 583264 202111 583266
rect 200836 583208 202050 583264
rect 202106 583208 202111 583264
rect 200836 583206 202111 583208
rect 280876 583264 283439 583266
rect 280876 583208 283378 583264
rect 283434 583208 283439 583264
rect 280876 583206 283439 583208
rect 122097 583203 122163 583206
rect 202045 583203 202111 583206
rect 283373 583203 283439 583206
rect 317965 582586 318031 582589
rect 320038 582586 320098 582624
rect 317965 582584 320098 582586
rect 317965 582528 317970 582584
rect 318026 582528 320098 582584
rect 317965 582526 320098 582528
rect 317965 582523 318031 582526
rect 457437 582314 457503 582317
rect 457437 582312 460092 582314
rect 457437 582256 457442 582312
rect 457498 582256 460092 582312
rect 457437 582254 460092 582256
rect 457437 582251 457503 582254
rect 58801 581090 58867 581093
rect 59494 581090 60076 581150
rect 139350 581098 140032 581158
rect 219390 581098 220064 581158
rect 138657 581090 138723 581093
rect 139350 581090 139410 581098
rect 58801 581088 59554 581090
rect 58801 581032 58806 581088
rect 58862 581032 59554 581088
rect 58801 581030 59554 581032
rect 138657 581088 139410 581090
rect 138657 581032 138662 581088
rect 138718 581032 139410 581088
rect 138657 581030 139410 581032
rect 217685 581090 217751 581093
rect 219390 581090 219450 581098
rect 217685 581088 219450 581090
rect 217685 581032 217690 581088
rect 217746 581032 219450 581088
rect 217685 581030 219450 581032
rect 58801 581027 58867 581030
rect 138657 581027 138723 581030
rect 217685 581027 217751 581030
rect 122005 580546 122071 580549
rect 202321 580546 202387 580549
rect 281809 580546 281875 580549
rect 120796 580544 122071 580546
rect 120796 580488 122010 580544
rect 122066 580488 122071 580544
rect 120796 580486 122071 580488
rect 200836 580544 202387 580546
rect 200836 580488 202326 580544
rect 202382 580488 202387 580544
rect 200836 580486 202387 580488
rect 280876 580544 281875 580546
rect 280876 580488 281814 580544
rect 281870 580488 281875 580544
rect 280876 580486 281875 580488
rect 122005 580483 122071 580486
rect 202321 580483 202387 580486
rect 281809 580483 281875 580486
rect -960 580002 480 580092
rect 3417 580002 3483 580005
rect -960 580000 3483 580002
rect -960 579944 3422 580000
rect 3478 579944 3483 580000
rect -960 579942 3483 579944
rect -960 579852 480 579942
rect 3417 579939 3483 579942
rect 512269 579594 512335 579597
rect 509956 579592 512335 579594
rect 509956 579536 512274 579592
rect 512330 579536 512335 579592
rect 509956 579534 512335 579536
rect 512269 579531 512335 579534
rect 428782 578370 428842 578544
rect 430665 578370 430731 578373
rect 428782 578368 430731 578370
rect 428782 578312 430670 578368
rect 430726 578312 430731 578368
rect 428782 578310 430731 578312
rect 430665 578307 430731 578310
rect 57053 577690 57119 577693
rect 59494 577690 60076 577750
rect 139350 577698 140032 577758
rect 219390 577698 220064 577758
rect 136725 577690 136791 577693
rect 139350 577690 139410 577698
rect 57053 577688 59554 577690
rect 57053 577632 57058 577688
rect 57114 577632 59554 577688
rect 57053 577630 59554 577632
rect 136725 577688 139410 577690
rect 136725 577632 136730 577688
rect 136786 577632 139410 577688
rect 136725 577630 139410 577632
rect 216029 577690 216095 577693
rect 219390 577690 219450 577698
rect 216029 577688 219450 577690
rect 216029 577632 216034 577688
rect 216090 577632 219450 577688
rect 216029 577630 219450 577632
rect 57053 577627 57119 577630
rect 136725 577627 136791 577630
rect 216029 577627 216095 577630
rect 317873 577282 317939 577285
rect 320038 577282 320098 577864
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect 317873 577280 320098 577282
rect 317873 577224 317878 577280
rect 317934 577224 320098 577280
rect 317873 577222 320098 577224
rect 317873 577219 317939 577222
rect 203333 577146 203399 577149
rect 283557 577146 283623 577149
rect 200836 577144 203399 577146
rect 120766 576874 120826 577116
rect 200836 577088 203338 577144
rect 203394 577088 203399 577144
rect 200836 577086 203399 577088
rect 280876 577144 283623 577146
rect 280876 577088 283562 577144
rect 283618 577088 283623 577144
rect 280876 577086 283623 577088
rect 203333 577083 203399 577086
rect 283557 577083 283623 577086
rect 120993 576874 121059 576877
rect 120766 576872 121059 576874
rect 120766 576816 120998 576872
rect 121054 576816 121059 576872
rect 120766 576814 121059 576816
rect 120993 576811 121059 576814
rect 457437 576194 457503 576197
rect 457437 576192 460092 576194
rect 457437 576136 457442 576192
rect 457498 576136 460092 576192
rect 457437 576134 460092 576136
rect 457437 576131 457503 576134
rect 57145 574970 57211 574973
rect 59494 574970 60076 575030
rect 139350 574978 140032 575038
rect 219390 574978 220064 575038
rect 137461 574970 137527 574973
rect 139350 574970 139410 574978
rect 57145 574968 59554 574970
rect 57145 574912 57150 574968
rect 57206 574912 59554 574968
rect 57145 574910 59554 574912
rect 137461 574968 139410 574970
rect 137461 574912 137466 574968
rect 137522 574912 139410 574968
rect 137461 574910 139410 574912
rect 216673 574970 216739 574973
rect 219390 574970 219450 574978
rect 216673 574968 219450 574970
rect 216673 574912 216678 574968
rect 216734 574912 219450 574968
rect 216673 574910 219450 574912
rect 57145 574907 57211 574910
rect 137461 574907 137527 574910
rect 216673 574907 216739 574910
rect 123477 574426 123543 574429
rect 203241 574426 203307 574429
rect 283465 574426 283531 574429
rect 120796 574424 123543 574426
rect 120796 574368 123482 574424
rect 123538 574368 123543 574424
rect 120796 574366 123543 574368
rect 200836 574424 203307 574426
rect 200836 574368 203246 574424
rect 203302 574368 203307 574424
rect 200836 574366 203307 574368
rect 280876 574424 283531 574426
rect 280876 574368 283470 574424
rect 283526 574368 283531 574424
rect 280876 574366 283531 574368
rect 123477 574363 123543 574366
rect 203241 574363 203307 574366
rect 283465 574363 283531 574366
rect 428782 572794 428842 573104
rect 430757 572794 430823 572797
rect 513281 572794 513347 572797
rect 428782 572792 430823 572794
rect 428782 572736 430762 572792
rect 430818 572736 430823 572792
rect 428782 572734 430823 572736
rect 509956 572792 513347 572794
rect 509956 572736 513286 572792
rect 513342 572736 513347 572792
rect 509956 572734 513347 572736
rect 430757 572731 430823 572734
rect 513281 572731 513347 572734
rect 317965 571842 318031 571845
rect 320038 571842 320098 572424
rect 317965 571840 320098 571842
rect 317965 571784 317970 571840
rect 318026 571784 320098 571840
rect 317965 571782 320098 571784
rect 317965 571779 318031 571782
rect 57329 571570 57395 571573
rect 59494 571570 60076 571630
rect 139350 571578 140032 571638
rect 219390 571578 220064 571638
rect 137553 571570 137619 571573
rect 139350 571570 139410 571578
rect 57329 571568 59554 571570
rect 57329 571512 57334 571568
rect 57390 571512 59554 571568
rect 57329 571510 59554 571512
rect 137553 571568 139410 571570
rect 137553 571512 137558 571568
rect 137614 571512 139410 571568
rect 137553 571510 139410 571512
rect 216673 571570 216739 571573
rect 219390 571570 219450 571578
rect 216673 571568 219450 571570
rect 216673 571512 216678 571568
rect 216734 571512 219450 571568
rect 216673 571510 219450 571512
rect 57329 571507 57395 571510
rect 137553 571507 137619 571510
rect 216673 571507 216739 571510
rect 121453 571026 121519 571029
rect 201493 571026 201559 571029
rect 283649 571026 283715 571029
rect 120796 571024 121519 571026
rect 120796 570968 121458 571024
rect 121514 570968 121519 571024
rect 120796 570966 121519 570968
rect 200836 571024 201559 571026
rect 200836 570968 201498 571024
rect 201554 570968 201559 571024
rect 200836 570966 201559 570968
rect 280876 571024 283715 571026
rect 280876 570968 283654 571024
rect 283710 570968 283715 571024
rect 280876 570966 283715 570968
rect 121453 570963 121519 570966
rect 201493 570963 201559 570966
rect 283649 570963 283715 570966
rect 58525 568850 58591 568853
rect 59494 568850 60076 568910
rect 139350 568858 140032 568918
rect 219390 568858 220064 568918
rect 138565 568850 138631 568853
rect 139350 568850 139410 568858
rect 58525 568848 59554 568850
rect 58525 568792 58530 568848
rect 58586 568792 59554 568848
rect 58525 568790 59554 568792
rect 138565 568848 139410 568850
rect 138565 568792 138570 568848
rect 138626 568792 139410 568848
rect 138565 568790 139410 568792
rect 219157 568850 219223 568853
rect 219390 568850 219450 568858
rect 219157 568848 219450 568850
rect 219157 568792 219162 568848
rect 219218 568792 219450 568848
rect 219157 568790 219450 568792
rect 58525 568787 58591 568790
rect 138565 568787 138631 568790
rect 219157 568787 219223 568790
rect 123569 568306 123635 568309
rect 201125 568306 201191 568309
rect 281533 568306 281599 568309
rect 120796 568304 123635 568306
rect 120796 568248 123574 568304
rect 123630 568248 123635 568304
rect 120796 568246 123635 568248
rect 200836 568304 201191 568306
rect 200836 568248 201130 568304
rect 201186 568248 201191 568304
rect 200836 568246 201191 568248
rect 280876 568304 281599 568306
rect 280876 568248 281538 568304
rect 281594 568248 281599 568304
rect 280876 568246 281599 568248
rect 123569 568243 123635 568246
rect 201125 568243 201191 568246
rect 281533 568243 281599 568246
rect 317045 568306 317111 568309
rect 317045 568304 320098 568306
rect 317045 568248 317050 568304
rect 317106 568248 320098 568304
rect 317045 568246 320098 568248
rect 317045 568243 317111 568246
rect 320038 567664 320098 568246
rect 428782 567762 428842 568344
rect 430849 567762 430915 567765
rect 428782 567760 430915 567762
rect 428782 567704 430854 567760
rect 430910 567704 430915 567760
rect 428782 567702 430915 567704
rect 430849 567699 430915 567702
rect -960 566796 480 567036
rect 57237 565450 57303 565453
rect 59494 565450 60076 565510
rect 139350 565458 140032 565518
rect 219390 565458 220064 565518
rect 138473 565450 138539 565453
rect 139350 565450 139410 565458
rect 57237 565448 59554 565450
rect 57237 565392 57242 565448
rect 57298 565392 59554 565448
rect 57237 565390 59554 565392
rect 138473 565448 139410 565450
rect 138473 565392 138478 565448
rect 138534 565392 139410 565448
rect 138473 565390 139410 565392
rect 217593 565450 217659 565453
rect 219390 565450 219450 565458
rect 217593 565448 219450 565450
rect 217593 565392 217598 565448
rect 217654 565392 219450 565448
rect 217593 565390 219450 565392
rect 57237 565387 57303 565390
rect 138473 565387 138539 565390
rect 217593 565387 217659 565390
rect 121085 564906 121151 564909
rect 203425 564906 203491 564909
rect 281257 564906 281323 564909
rect 120796 564904 121151 564906
rect 120796 564848 121090 564904
rect 121146 564848 121151 564904
rect 120796 564846 121151 564848
rect 200836 564904 203491 564906
rect 200836 564848 203430 564904
rect 203486 564848 203491 564904
rect 200836 564846 203491 564848
rect 280876 564904 281323 564906
rect 280876 564848 281262 564904
rect 281318 564848 281323 564904
rect 280876 564846 281323 564848
rect 121085 564843 121151 564846
rect 203425 564843 203491 564846
rect 281257 564843 281323 564846
rect 583520 564212 584960 564452
rect 428782 563138 428842 563584
rect 430941 563138 431007 563141
rect 428782 563136 431007 563138
rect 428782 563080 430946 563136
rect 431002 563080 431007 563136
rect 428782 563078 431007 563080
rect 430941 563075 431007 563078
rect 139393 562798 139459 562801
rect 139393 562796 140032 562798
rect 59537 562790 59603 562793
rect 59537 562788 60076 562790
rect 59537 562732 59542 562788
rect 59598 562732 60076 562788
rect 139393 562740 139398 562796
rect 139454 562740 140032 562796
rect 139393 562738 140032 562740
rect 219390 562738 220064 562798
rect 139393 562735 139459 562738
rect 59537 562730 60076 562732
rect 217133 562730 217199 562733
rect 219390 562730 219450 562738
rect 59537 562727 59603 562730
rect 217133 562728 219450 562730
rect 217133 562672 217138 562728
rect 217194 562672 219450 562728
rect 217133 562670 219450 562672
rect 217133 562667 217199 562670
rect 318333 562322 318399 562325
rect 320038 562322 320098 562904
rect 318333 562320 320098 562322
rect 318333 562264 318338 562320
rect 318394 562264 320098 562320
rect 318333 562262 320098 562264
rect 318333 562259 318399 562262
rect 121177 562186 121243 562189
rect 201217 562186 201283 562189
rect 281993 562186 282059 562189
rect 120796 562184 121243 562186
rect 120796 562128 121182 562184
rect 121238 562128 121243 562184
rect 120796 562126 121243 562128
rect 200836 562184 201283 562186
rect 200836 562128 201222 562184
rect 201278 562128 201283 562184
rect 200836 562126 201283 562128
rect 280876 562184 282059 562186
rect 280876 562128 281998 562184
rect 282054 562128 282059 562184
rect 280876 562126 282059 562128
rect 121177 562123 121243 562126
rect 201217 562123 201283 562126
rect 281993 562123 282059 562126
rect 428414 558245 428474 558824
rect 428365 558240 428474 558245
rect 428365 558184 428370 558240
rect 428426 558184 428474 558240
rect 428365 558182 428474 558184
rect 428365 558179 428431 558182
rect 317413 557698 317479 557701
rect 320038 557698 320098 558144
rect 317413 557696 320098 557698
rect 317413 557640 317418 557696
rect 317474 557640 320098 557696
rect 317413 557638 320098 557640
rect 317413 557635 317479 557638
rect -960 553740 480 553980
rect 317965 553482 318031 553485
rect 428782 553482 428842 554064
rect 429469 553482 429535 553485
rect 317965 553480 320098 553482
rect 317965 553424 317970 553480
rect 318026 553424 320098 553480
rect 317965 553422 320098 553424
rect 428782 553480 429535 553482
rect 428782 553424 429474 553480
rect 429530 553424 429535 553480
rect 428782 553422 429535 553424
rect 317965 553419 318031 553422
rect 320038 553384 320098 553422
rect 429469 553419 429535 553422
rect 583520 551020 584960 551260
rect 431033 549402 431099 549405
rect 428782 549400 431099 549402
rect 428782 549344 431038 549400
rect 431094 549344 431099 549400
rect 428782 549342 431099 549344
rect 428782 549304 428842 549342
rect 431033 549339 431099 549342
rect 317965 549130 318031 549133
rect 317965 549128 320098 549130
rect 317965 549072 317970 549128
rect 318026 549072 320098 549128
rect 317965 549070 320098 549072
rect 317965 549067 318031 549070
rect 320038 548624 320098 549070
rect 428782 543962 428842 544544
rect 431125 543962 431191 543965
rect 428782 543960 431191 543962
rect 428782 543904 431130 543960
rect 431186 543904 431191 543960
rect 428782 543902 431191 543904
rect 431125 543899 431191 543902
rect 317965 543826 318031 543829
rect 320038 543826 320098 543864
rect 317965 543824 320098 543826
rect 317965 543768 317970 543824
rect 318026 543768 320098 543824
rect 317965 543766 320098 543768
rect 317965 543763 318031 543766
rect 255129 543282 255195 543285
rect 318241 543282 318307 543285
rect 255129 543280 318307 543282
rect 255129 543224 255134 543280
rect 255190 543224 318246 543280
rect 318302 543224 318307 543280
rect 255129 543222 318307 543224
rect 255129 543219 255195 543222
rect 318241 543219 318307 543222
rect 256509 543146 256575 543149
rect 285029 543146 285095 543149
rect 256509 543144 285095 543146
rect 256509 543088 256514 543144
rect 256570 543088 285034 543144
rect 285090 543088 285095 543144
rect 256509 543086 285095 543088
rect 256509 543083 256575 543086
rect 285029 543083 285095 543086
rect 239397 543010 239463 543013
rect 280654 543010 280660 543012
rect 239397 543008 280660 543010
rect 239397 542952 239402 543008
rect 239458 542952 280660 543008
rect 239397 542950 280660 542952
rect 239397 542947 239463 542950
rect 280654 542948 280660 542950
rect 280724 542948 280730 543012
rect 285949 542874 286015 542877
rect 317045 542874 317111 542877
rect 285949 542872 317111 542874
rect 285949 542816 285954 542872
rect 286010 542816 317050 542872
rect 317106 542816 317111 542872
rect 285949 542814 317111 542816
rect 285949 542811 286015 542814
rect 317045 542811 317111 542814
rect 248689 542738 248755 542741
rect 300209 542738 300275 542741
rect 248689 542736 300275 542738
rect 248689 542680 248694 542736
rect 248750 542680 300214 542736
rect 300270 542680 300275 542736
rect 248689 542678 300275 542680
rect 248689 542675 248755 542678
rect 300209 542675 300275 542678
rect 241513 542602 241579 542605
rect 299974 542602 299980 542604
rect 241513 542600 299980 542602
rect 241513 542544 241518 542600
rect 241574 542544 299980 542600
rect 241513 542542 299980 542544
rect 241513 542539 241579 542542
rect 299974 542540 299980 542542
rect 300044 542540 300050 542604
rect 286685 542466 286751 542469
rect 301497 542466 301563 542469
rect 286685 542464 301563 542466
rect 286685 542408 286690 542464
rect 286746 542408 301502 542464
rect 301558 542408 301563 542464
rect 286685 542406 301563 542408
rect 286685 542403 286751 542406
rect 301497 542403 301563 542406
rect 284293 541650 284359 541653
rect 316769 541650 316835 541653
rect 284293 541648 316835 541650
rect 284293 541592 284298 541648
rect 284354 541592 316774 541648
rect 316830 541592 316835 541648
rect 284293 541590 316835 541592
rect 284293 541587 284359 541590
rect 316769 541587 316835 541590
rect 291653 541378 291719 541381
rect 314193 541378 314259 541381
rect 291653 541376 314259 541378
rect 291653 541320 291658 541376
rect 291714 541320 314198 541376
rect 314254 541320 314259 541376
rect 291653 541318 314259 541320
rect 291653 541315 291719 541318
rect 314193 541315 314259 541318
rect 294505 541242 294571 541245
rect 316953 541242 317019 541245
rect 294505 541240 317019 541242
rect 294505 541184 294510 541240
rect 294566 541184 316958 541240
rect 317014 541184 317019 541240
rect 294505 541182 317019 541184
rect 294505 541179 294571 541182
rect 316953 541179 317019 541182
rect 264421 541106 264487 541109
rect 320582 541106 320588 541108
rect 264421 541104 320588 541106
rect 264421 541048 264426 541104
rect 264482 541048 320588 541104
rect 264421 541046 320588 541048
rect 264421 541043 264487 541046
rect 320582 541044 320588 541046
rect 320652 541044 320658 541108
rect -960 540684 480 540924
rect 428782 539610 428842 539784
rect 431217 539610 431283 539613
rect 428782 539608 431283 539610
rect 428782 539552 431222 539608
rect 431278 539552 431283 539608
rect 428782 539550 431283 539552
rect 431217 539547 431283 539550
rect 318057 539338 318123 539341
rect 318057 539336 320098 539338
rect 318057 539280 318062 539336
rect 318118 539280 320098 539336
rect 318057 539278 320098 539280
rect 318057 539275 318123 539278
rect 320038 539104 320098 539278
rect 583520 537692 584960 537932
rect 317597 534986 317663 534989
rect 317597 534984 320098 534986
rect 317597 534928 317602 534984
rect 317658 534928 320098 534984
rect 317597 534926 320098 534928
rect 317597 534923 317663 534926
rect 320038 534344 320098 534926
rect 428782 534442 428842 535024
rect 431309 534442 431375 534445
rect 428782 534440 431375 534442
rect 428782 534384 431314 534440
rect 431370 534384 431375 534440
rect 428782 534382 431375 534384
rect 431309 534379 431375 534382
rect 302325 532402 302391 532405
rect 299828 532400 302391 532402
rect 299828 532344 302330 532400
rect 302386 532344 302391 532400
rect 299828 532342 302391 532344
rect 302325 532339 302391 532342
rect 429377 530906 429443 530909
rect 428782 530904 429443 530906
rect 428782 530848 429382 530904
rect 429438 530848 429443 530904
rect 428782 530846 429443 530848
rect 428782 530264 428842 530846
rect 429377 530843 429443 530846
rect 317597 529818 317663 529821
rect 317597 529816 320098 529818
rect 317597 529760 317602 529816
rect 317658 529760 320098 529816
rect 317597 529758 320098 529760
rect 317597 529755 317663 529758
rect 320038 529584 320098 529758
rect -960 527764 480 528004
rect 317689 525466 317755 525469
rect 317689 525464 320098 525466
rect 317689 525408 317694 525464
rect 317750 525408 320098 525464
rect 317689 525406 320098 525408
rect 317689 525403 317755 525406
rect 320038 524824 320098 525406
rect 428782 524922 428842 525504
rect 430665 524922 430731 524925
rect 428782 524920 430731 524922
rect 428782 524864 430670 524920
rect 430726 524864 430731 524920
rect 428782 524862 430731 524864
rect 430665 524859 430731 524862
rect 583520 524364 584960 524604
rect 427813 520298 427879 520301
rect 428230 520298 428290 520744
rect 427813 520296 428290 520298
rect 427813 520240 427818 520296
rect 427874 520240 428290 520296
rect 427813 520238 428290 520240
rect 427813 520235 427879 520238
rect 318241 520162 318307 520165
rect 430614 520162 430620 520164
rect 318241 520160 430620 520162
rect 318241 520104 318246 520160
rect 318302 520104 430620 520160
rect 318241 520102 430620 520104
rect 318241 520099 318307 520102
rect 430614 520100 430620 520102
rect 430684 520100 430690 520164
rect 300209 518802 300275 518805
rect 430798 518802 430804 518804
rect 300209 518800 430804 518802
rect 300209 518744 300214 518800
rect 300270 518744 430804 518800
rect 300209 518742 430804 518744
rect 300209 518739 300275 518742
rect 430798 518740 430804 518742
rect 430868 518740 430874 518804
rect 320766 518604 320772 518668
rect 320836 518666 320842 518668
rect 374453 518666 374519 518669
rect 320836 518664 374519 518666
rect 320836 518608 374458 518664
rect 374514 518608 374519 518664
rect 320836 518606 374519 518608
rect 320836 518604 320842 518606
rect 374453 518603 374519 518606
rect 312537 518530 312603 518533
rect 356237 518530 356303 518533
rect 312537 518528 356303 518530
rect 312537 518472 312542 518528
rect 312598 518472 356242 518528
rect 356298 518472 356303 518528
rect 312537 518470 356303 518472
rect 312537 518467 312603 518470
rect 356237 518467 356303 518470
rect 319713 518394 319779 518397
rect 337653 518394 337719 518397
rect 319713 518392 337719 518394
rect 319713 518336 319718 518392
rect 319774 518336 337658 518392
rect 337714 518336 337719 518392
rect 319713 518334 337719 518336
rect 319713 518331 319779 518334
rect 337653 518331 337719 518334
rect 302601 517442 302667 517445
rect 299828 517440 302667 517442
rect 299828 517384 302606 517440
rect 302662 517384 302667 517440
rect 299828 517382 302667 517384
rect 302601 517379 302667 517382
rect 299974 517244 299980 517308
rect 300044 517306 300050 517308
rect 430982 517306 430988 517308
rect 300044 517246 430988 517306
rect 300044 517244 300050 517246
rect 430982 517244 430988 517246
rect 431052 517244 431058 517308
rect -960 514858 480 514948
rect 3601 514858 3667 514861
rect -960 514856 3667 514858
rect -960 514800 3606 514856
rect 3662 514800 3667 514856
rect -960 514798 3667 514800
rect -960 514708 480 514798
rect 3601 514795 3667 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect 57697 509962 57763 509965
rect 57881 509962 57947 509965
rect 57697 509960 60076 509962
rect 57697 509904 57702 509960
rect 57758 509904 57886 509960
rect 57942 509904 60076 509960
rect 57697 509902 60076 509904
rect 57697 509899 57763 509902
rect 57881 509899 57947 509902
rect 302233 502482 302299 502485
rect 299828 502480 302299 502482
rect 299828 502424 302238 502480
rect 302294 502424 302299 502480
rect 299828 502422 302299 502424
rect 302233 502419 302299 502422
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 302877 487522 302943 487525
rect 299828 487520 302943 487522
rect 299828 487464 302882 487520
rect 302938 487464 302943 487520
rect 299828 487462 302943 487464
rect 302877 487459 302943 487462
rect 360878 485012 360884 485076
rect 360948 485074 360954 485076
rect 391933 485074 391999 485077
rect 360948 485072 391999 485074
rect 360948 485016 391938 485072
rect 391994 485016 391999 485072
rect 360948 485014 391999 485016
rect 360948 485012 360954 485014
rect 391933 485011 391999 485014
rect 583520 484516 584960 484756
rect 363454 483652 363460 483716
rect 363524 483714 363530 483716
rect 488574 483714 488580 483716
rect 363524 483654 488580 483714
rect 363524 483652 363530 483654
rect 488574 483652 488580 483654
rect 488644 483652 488650 483716
rect 364926 482156 364932 482220
rect 364996 482218 365002 482220
rect 483013 482218 483079 482221
rect 364996 482216 483079 482218
rect 364996 482160 483018 482216
rect 483074 482160 483079 482216
rect 364996 482158 483079 482160
rect 364996 482156 365002 482158
rect 483013 482155 483079 482158
rect 366357 480858 366423 480861
rect 506606 480858 506612 480860
rect 366357 480856 506612 480858
rect 366357 480800 366362 480856
rect 366418 480800 506612 480856
rect 366357 480798 506612 480800
rect 366357 480795 366423 480798
rect 506606 480796 506612 480798
rect 506676 480796 506682 480860
rect 365110 479708 365116 479772
rect 365180 479770 365186 479772
rect 506473 479770 506539 479773
rect 365180 479768 506539 479770
rect 365180 479712 506478 479768
rect 506534 479712 506539 479768
rect 365180 479710 506539 479712
rect 365180 479708 365186 479710
rect 506473 479707 506539 479710
rect 208894 479572 208900 479636
rect 208964 479634 208970 479636
rect 457529 479634 457595 479637
rect 208964 479632 457595 479634
rect 208964 479576 457534 479632
rect 457590 479576 457595 479632
rect 208964 479574 457595 479576
rect 208964 479572 208970 479574
rect 457529 479571 457595 479574
rect 206134 479436 206140 479500
rect 206204 479498 206210 479500
rect 476062 479498 476068 479500
rect 206204 479438 476068 479498
rect 206204 479436 206210 479438
rect 476062 479436 476068 479438
rect 476132 479436 476138 479500
rect 73429 478954 73495 478957
rect 72926 478952 73495 478954
rect 72926 478896 73434 478952
rect 73490 478896 73495 478952
rect 72926 478894 73495 478896
rect 55070 478756 55076 478820
rect 55140 478818 55146 478820
rect 72049 478818 72115 478821
rect 55140 478816 72115 478818
rect 55140 478760 72054 478816
rect 72110 478760 72115 478816
rect 55140 478758 72115 478760
rect 55140 478756 55146 478758
rect 72049 478755 72115 478758
rect 54886 478620 54892 478684
rect 54956 478682 54962 478684
rect 72926 478682 72986 478894
rect 73429 478891 73495 478894
rect 107745 478954 107811 478957
rect 198774 478954 198780 478956
rect 107745 478952 198780 478954
rect 107745 478896 107750 478952
rect 107806 478896 198780 478952
rect 107745 478894 198780 478896
rect 107745 478891 107811 478894
rect 198774 478892 198780 478894
rect 198844 478892 198850 478956
rect 73153 478818 73219 478821
rect 79501 478818 79567 478821
rect 73153 478816 79567 478818
rect 73153 478760 73158 478816
rect 73214 478760 79506 478816
rect 79562 478760 79567 478816
rect 73153 478758 79567 478760
rect 73153 478755 73219 478758
rect 79501 478755 79567 478758
rect 170213 478818 170279 478821
rect 198222 478818 198228 478820
rect 170213 478816 198228 478818
rect 170213 478760 170218 478816
rect 170274 478760 198228 478816
rect 170213 478758 198228 478760
rect 170213 478755 170279 478758
rect 198222 478756 198228 478758
rect 198292 478756 198298 478820
rect 235901 478818 235967 478821
rect 360694 478818 360700 478820
rect 235901 478816 360700 478818
rect 235901 478760 235906 478816
rect 235962 478760 360700 478816
rect 235901 478758 360700 478760
rect 235901 478755 235967 478758
rect 360694 478756 360700 478758
rect 360764 478756 360770 478820
rect 54956 478622 72986 478682
rect 73153 478682 73219 478685
rect 77753 478682 77819 478685
rect 73153 478680 77819 478682
rect 73153 478624 73158 478680
rect 73214 478624 77758 478680
rect 77814 478624 77819 478680
rect 73153 478622 77819 478624
rect 54956 478620 54962 478622
rect 73153 478619 73219 478622
rect 77753 478619 77819 478622
rect 163589 478682 163655 478685
rect 196566 478682 196572 478684
rect 163589 478680 196572 478682
rect 163589 478624 163594 478680
rect 163650 478624 196572 478680
rect 163589 478622 196572 478624
rect 163589 478619 163655 478622
rect 196566 478620 196572 478622
rect 196636 478620 196642 478684
rect 205633 478682 205699 478685
rect 206870 478682 206876 478684
rect 205633 478680 206876 478682
rect 205633 478624 205638 478680
rect 205694 478624 206876 478680
rect 205633 478622 206876 478624
rect 205633 478619 205699 478622
rect 206870 478620 206876 478622
rect 206940 478620 206946 478684
rect 213913 478682 213979 478685
rect 214782 478682 214788 478684
rect 213913 478680 214788 478682
rect 213913 478624 213918 478680
rect 213974 478624 214788 478680
rect 213913 478622 214788 478624
rect 213913 478619 213979 478622
rect 214782 478620 214788 478622
rect 214852 478620 214858 478684
rect 235441 478682 235507 478685
rect 371734 478682 371740 478684
rect 235441 478680 371740 478682
rect 235441 478624 235446 478680
rect 235502 478624 371740 478680
rect 235441 478622 371740 478624
rect 235441 478619 235507 478622
rect 371734 478620 371740 478622
rect 371804 478620 371810 478684
rect 55438 478484 55444 478548
rect 55508 478546 55514 478548
rect 147305 478546 147371 478549
rect 198038 478546 198044 478548
rect 55508 478486 74550 478546
rect 55508 478484 55514 478486
rect 54702 478348 54708 478412
rect 54772 478410 54778 478412
rect 74490 478410 74550 478486
rect 147305 478544 198044 478546
rect 147305 478488 147310 478544
rect 147366 478488 198044 478544
rect 147305 478486 198044 478488
rect 147305 478483 147371 478486
rect 198038 478484 198044 478486
rect 198108 478484 198114 478548
rect 204345 478546 204411 478549
rect 205398 478546 205404 478548
rect 204345 478544 205404 478546
rect 204345 478488 204350 478544
rect 204406 478488 205404 478544
rect 204345 478486 205404 478488
rect 204345 478483 204411 478486
rect 205398 478484 205404 478486
rect 205468 478484 205474 478548
rect 208485 478546 208551 478549
rect 209262 478546 209268 478548
rect 208485 478544 209268 478546
rect 208485 478488 208490 478544
rect 208546 478488 209268 478544
rect 208485 478486 209268 478488
rect 208485 478483 208551 478486
rect 209262 478484 209268 478486
rect 209332 478484 209338 478548
rect 230565 478546 230631 478549
rect 367686 478546 367692 478548
rect 230565 478544 367692 478546
rect 230565 478488 230570 478544
rect 230626 478488 367692 478544
rect 230565 478486 367692 478488
rect 230565 478483 230631 478486
rect 367686 478484 367692 478486
rect 367756 478484 367762 478548
rect 74625 478410 74691 478413
rect 54772 478350 69674 478410
rect 74490 478408 74691 478410
rect 74490 478352 74630 478408
rect 74686 478352 74691 478408
rect 74490 478350 74691 478352
rect 54772 478348 54778 478350
rect 52310 478212 52316 478276
rect 52380 478274 52386 478276
rect 66253 478274 66319 478277
rect 52380 478272 66319 478274
rect 52380 478216 66258 478272
rect 66314 478216 66319 478272
rect 52380 478214 66319 478216
rect 69614 478274 69674 478350
rect 74625 478347 74691 478350
rect 148225 478410 148291 478413
rect 200614 478410 200620 478412
rect 148225 478408 200620 478410
rect 148225 478352 148230 478408
rect 148286 478352 200620 478408
rect 148225 478350 200620 478352
rect 148225 478347 148291 478350
rect 200614 478348 200620 478350
rect 200684 478348 200690 478412
rect 205633 478410 205699 478413
rect 206502 478410 206508 478412
rect 205633 478408 206508 478410
rect 205633 478352 205638 478408
rect 205694 478352 206508 478408
rect 205633 478350 206508 478352
rect 205633 478347 205699 478350
rect 206502 478348 206508 478350
rect 206572 478348 206578 478412
rect 231485 478410 231551 478413
rect 370446 478410 370452 478412
rect 231485 478408 370452 478410
rect 231485 478352 231490 478408
rect 231546 478352 370452 478408
rect 231485 478350 370452 478352
rect 231485 478347 231551 478350
rect 370446 478348 370452 478350
rect 370516 478348 370522 478412
rect 374494 478348 374500 478412
rect 374564 478410 374570 478412
rect 511993 478410 512059 478413
rect 374564 478408 512059 478410
rect 374564 478352 511998 478408
rect 512054 478352 512059 478408
rect 374564 478350 512059 478352
rect 374564 478348 374570 478350
rect 511993 478347 512059 478350
rect 76005 478274 76071 478277
rect 69614 478272 76071 478274
rect 69614 478216 76010 478272
rect 76066 478216 76071 478272
rect 69614 478214 76071 478216
rect 52380 478212 52386 478214
rect 66253 478211 66319 478214
rect 76005 478211 76071 478214
rect 145557 478274 145623 478277
rect 197854 478274 197860 478276
rect 145557 478272 197860 478274
rect 145557 478216 145562 478272
rect 145618 478216 197860 478272
rect 145557 478214 197860 478216
rect 145557 478211 145623 478214
rect 197854 478212 197860 478214
rect 197924 478212 197930 478276
rect 200113 478274 200179 478277
rect 200982 478274 200988 478276
rect 200113 478272 200988 478274
rect 200113 478216 200118 478272
rect 200174 478216 200988 478272
rect 200113 478214 200988 478216
rect 200113 478211 200179 478214
rect 200982 478212 200988 478214
rect 201052 478212 201058 478276
rect 219198 478212 219204 478276
rect 219268 478274 219274 478276
rect 226149 478274 226215 478277
rect 219268 478272 226215 478274
rect 219268 478216 226154 478272
rect 226210 478216 226215 478272
rect 219268 478214 226215 478216
rect 219268 478212 219274 478214
rect 226149 478211 226215 478214
rect 233693 478274 233759 478277
rect 375966 478274 375972 478276
rect 233693 478272 375972 478274
rect 233693 478216 233698 478272
rect 233754 478216 375972 478272
rect 233693 478214 375972 478216
rect 233693 478211 233759 478214
rect 375966 478212 375972 478214
rect 376036 478212 376042 478276
rect 46790 478076 46796 478140
rect 46860 478138 46866 478140
rect 80789 478138 80855 478141
rect 46860 478136 80855 478138
rect 46860 478080 80794 478136
rect 80850 478080 80855 478136
rect 46860 478078 80855 478080
rect 46860 478076 46866 478078
rect 80789 478075 80855 478078
rect 145097 478138 145163 478141
rect 202086 478138 202092 478140
rect 145097 478136 202092 478138
rect 145097 478080 145102 478136
rect 145158 478080 202092 478136
rect 145097 478078 202092 478080
rect 145097 478075 145163 478078
rect 202086 478076 202092 478078
rect 202156 478076 202162 478140
rect 212533 478138 212599 478141
rect 213678 478138 213684 478140
rect 212533 478136 213684 478138
rect 212533 478080 212538 478136
rect 212594 478080 213684 478136
rect 212533 478078 213684 478080
rect 212533 478075 212599 478078
rect 213678 478076 213684 478078
rect 213748 478076 213754 478140
rect 232313 478138 232379 478141
rect 374678 478138 374684 478140
rect 232313 478136 374684 478138
rect 232313 478080 232318 478136
rect 232374 478080 374684 478136
rect 232313 478078 374684 478080
rect 232313 478075 232379 478078
rect 374678 478076 374684 478078
rect 374748 478076 374754 478140
rect 59302 477940 59308 478004
rect 59372 478002 59378 478004
rect 72509 478002 72575 478005
rect 59372 478000 72575 478002
rect 59372 477944 72514 478000
rect 72570 477944 72575 478000
rect 59372 477942 72575 477944
rect 59372 477940 59378 477942
rect 72509 477939 72575 477942
rect 185669 478002 185735 478005
rect 196750 478002 196756 478004
rect 185669 478000 196756 478002
rect 185669 477944 185674 478000
rect 185730 477944 196756 478000
rect 185669 477942 196756 477944
rect 185669 477939 185735 477942
rect 196750 477940 196756 477942
rect 196820 477940 196826 478004
rect 201493 478002 201559 478005
rect 202638 478002 202644 478004
rect 201493 478000 202644 478002
rect 201493 477944 201498 478000
rect 201554 477944 202644 478000
rect 201493 477942 202644 477944
rect 201493 477939 201559 477942
rect 202638 477940 202644 477942
rect 202708 477940 202714 478004
rect 234521 478002 234587 478005
rect 357934 478002 357940 478004
rect 234521 478000 357940 478002
rect 234521 477944 234526 478000
rect 234582 477944 357940 478000
rect 234521 477942 357940 477944
rect 234521 477939 234587 477942
rect 357934 477940 357940 477942
rect 358004 477940 358010 478004
rect 66253 477866 66319 477869
rect 76465 477866 76531 477869
rect 66253 477864 76531 477866
rect 66253 477808 66258 477864
rect 66314 477808 76470 477864
rect 76526 477808 76531 477864
rect 66253 477806 76531 477808
rect 66253 477803 66319 477806
rect 76465 477803 76531 477806
rect 357433 477866 357499 477869
rect 358118 477866 358124 477868
rect 357433 477864 358124 477866
rect 357433 477808 357438 477864
rect 357494 477808 358124 477864
rect 357433 477806 358124 477808
rect 357433 477803 357499 477806
rect 358118 477804 358124 477806
rect 358188 477804 358194 477868
rect 197353 477730 197419 477733
rect 198590 477730 198596 477732
rect 197353 477728 198596 477730
rect 197353 477672 197358 477728
rect 197414 477672 198596 477728
rect 197353 477670 198596 477672
rect 197353 477667 197419 477670
rect 198590 477668 198596 477670
rect 198660 477668 198666 477732
rect 200665 477730 200731 477733
rect 201350 477730 201356 477732
rect 200665 477728 201356 477730
rect 200665 477672 200670 477728
rect 200726 477672 201356 477728
rect 200665 477670 201356 477672
rect 200665 477667 200731 477670
rect 201350 477668 201356 477670
rect 201420 477668 201426 477732
rect 216990 477668 216996 477732
rect 217060 477730 217066 477732
rect 217777 477730 217843 477733
rect 217060 477728 217843 477730
rect 217060 477672 217782 477728
rect 217838 477672 217843 477728
rect 217060 477670 217843 477672
rect 217060 477668 217066 477670
rect 217777 477667 217843 477670
rect 50889 477596 50955 477597
rect 50838 477594 50844 477596
rect 50798 477534 50844 477594
rect 50908 477592 50955 477596
rect 50950 477536 50955 477592
rect 50838 477532 50844 477534
rect 50908 477532 50955 477536
rect 53230 477532 53236 477596
rect 53300 477594 53306 477596
rect 53465 477594 53531 477597
rect 53300 477592 53531 477594
rect 53300 477536 53470 477592
rect 53526 477536 53531 477592
rect 53300 477534 53531 477536
rect 53300 477532 53306 477534
rect 50889 477531 50955 477532
rect 53465 477531 53531 477534
rect 216949 477594 217015 477597
rect 217542 477594 217548 477596
rect 216949 477592 217548 477594
rect 216949 477536 216954 477592
rect 217010 477536 217548 477592
rect 216949 477534 217548 477536
rect 216949 477531 217015 477534
rect 217542 477532 217548 477534
rect 217612 477532 217618 477596
rect 219934 477532 219940 477596
rect 220004 477594 220010 477596
rect 223113 477594 223179 477597
rect 220004 477592 223179 477594
rect 220004 477536 223118 477592
rect 223174 477536 223179 477592
rect 220004 477534 223179 477536
rect 220004 477532 220010 477534
rect 223113 477531 223179 477534
rect 255221 476914 255287 476917
rect 359406 476914 359412 476916
rect 255221 476912 359412 476914
rect 255221 476856 255226 476912
rect 255282 476856 359412 476912
rect 255221 476854 359412 476856
rect 255221 476851 255287 476854
rect 359406 476852 359412 476854
rect 359476 476852 359482 476916
rect 153101 476778 153167 476781
rect 209814 476778 209820 476780
rect 153101 476776 209820 476778
rect 153101 476720 153106 476776
rect 153162 476720 209820 476776
rect 153101 476718 209820 476720
rect 153101 476715 153167 476718
rect 209814 476716 209820 476718
rect 209884 476716 209890 476780
rect 222193 476778 222259 476781
rect 367870 476778 367876 476780
rect 222193 476776 367876 476778
rect 222193 476720 222198 476776
rect 222254 476720 367876 476776
rect 222193 476718 367876 476720
rect 222193 476715 222259 476718
rect 367870 476716 367876 476718
rect 367940 476716 367946 476780
rect 46841 475962 46907 475965
rect 66345 475962 66411 475965
rect 46841 475960 66411 475962
rect 46841 475904 46846 475960
rect 46902 475904 66350 475960
rect 66406 475904 66411 475960
rect 46841 475902 66411 475904
rect 46841 475899 46907 475902
rect 66345 475899 66411 475902
rect -960 475540 480 475780
rect 57094 475764 57100 475828
rect 57164 475826 57170 475828
rect 121361 475826 121427 475829
rect 57164 475824 121427 475826
rect 57164 475768 121366 475824
rect 121422 475768 121427 475824
rect 57164 475766 121427 475768
rect 57164 475764 57170 475766
rect 121361 475763 121427 475766
rect 50337 475690 50403 475693
rect 120901 475690 120967 475693
rect 50337 475688 120967 475690
rect 50337 475632 50342 475688
rect 50398 475632 120906 475688
rect 120962 475632 120967 475688
rect 50337 475630 120967 475632
rect 50337 475627 50403 475630
rect 120901 475627 120967 475630
rect 46473 475554 46539 475557
rect 120441 475554 120507 475557
rect 46473 475552 120507 475554
rect 46473 475496 46478 475552
rect 46534 475496 120446 475552
rect 120502 475496 120507 475552
rect 46473 475494 120507 475496
rect 46473 475491 46539 475494
rect 120441 475491 120507 475494
rect 155677 475554 155743 475557
rect 215334 475554 215340 475556
rect 155677 475552 215340 475554
rect 155677 475496 155682 475552
rect 155738 475496 215340 475552
rect 155677 475494 215340 475496
rect 155677 475491 155743 475494
rect 215334 475492 215340 475494
rect 215404 475492 215410 475556
rect 231853 475554 231919 475557
rect 371918 475554 371924 475556
rect 231853 475552 371924 475554
rect 231853 475496 231858 475552
rect 231914 475496 371924 475552
rect 231853 475494 371924 475496
rect 231853 475491 231919 475494
rect 371918 475492 371924 475494
rect 371988 475492 371994 475556
rect 3601 475418 3667 475421
rect 429285 475418 429351 475421
rect 3601 475416 429351 475418
rect 3601 475360 3606 475416
rect 3662 475360 429290 475416
rect 429346 475360 429351 475416
rect 3601 475358 429351 475360
rect 3601 475355 3667 475358
rect 429285 475355 429351 475358
rect 171593 474330 171659 474333
rect 213310 474330 213316 474332
rect 171593 474328 213316 474330
rect 171593 474272 171598 474328
rect 171654 474272 213316 474328
rect 171593 474270 213316 474272
rect 171593 474267 171659 474270
rect 213310 474268 213316 474270
rect 213380 474268 213386 474332
rect 252737 474330 252803 474333
rect 377254 474330 377260 474332
rect 252737 474328 377260 474330
rect 252737 474272 252742 474328
rect 252798 474272 377260 474328
rect 252737 474270 377260 474272
rect 252737 474267 252803 474270
rect 377254 474268 377260 474270
rect 377324 474268 377330 474332
rect 150433 474194 150499 474197
rect 214414 474194 214420 474196
rect 150433 474192 214420 474194
rect 150433 474136 150438 474192
rect 150494 474136 214420 474192
rect 150433 474134 214420 474136
rect 150433 474131 150499 474134
rect 214414 474132 214420 474134
rect 214484 474132 214490 474196
rect 233233 474194 233299 474197
rect 363638 474194 363644 474196
rect 233233 474192 363644 474194
rect 233233 474136 233238 474192
rect 233294 474136 363644 474192
rect 233233 474134 363644 474136
rect 233233 474131 233299 474134
rect 363638 474132 363644 474134
rect 363708 474132 363714 474196
rect 116301 474058 116367 474061
rect 198958 474058 198964 474060
rect 116301 474056 198964 474058
rect 116301 474000 116306 474056
rect 116362 474000 198964 474056
rect 116301 473998 198964 474000
rect 116301 473995 116367 473998
rect 198958 473996 198964 473998
rect 199028 473996 199034 474060
rect 210366 473996 210372 474060
rect 210436 474058 210442 474060
rect 512085 474058 512151 474061
rect 210436 474056 512151 474058
rect 210436 474000 512090 474056
rect 512146 474000 512151 474056
rect 210436 473998 512151 474000
rect 210436 473996 210442 473998
rect 512085 473995 512151 473998
rect 43989 472970 44055 472973
rect 81249 472970 81315 472973
rect 43989 472968 81315 472970
rect 43989 472912 43994 472968
rect 44050 472912 81254 472968
rect 81310 472912 81315 472968
rect 43989 472910 81315 472912
rect 43989 472907 44055 472910
rect 81249 472907 81315 472910
rect 58985 472834 59051 472837
rect 95785 472834 95851 472837
rect 58985 472832 95851 472834
rect 58985 472776 58990 472832
rect 59046 472776 95790 472832
rect 95846 472776 95851 472832
rect 58985 472774 95851 472776
rect 58985 472771 59051 472774
rect 95785 472771 95851 472774
rect 57278 472636 57284 472700
rect 57348 472698 57354 472700
rect 122649 472698 122715 472701
rect 57348 472696 122715 472698
rect 57348 472640 122654 472696
rect 122710 472640 122715 472696
rect 57348 472638 122715 472640
rect 57348 472636 57354 472638
rect 122649 472635 122715 472638
rect 179965 472698 180031 472701
rect 217174 472698 217180 472700
rect 179965 472696 217180 472698
rect 179965 472640 179970 472696
rect 180026 472640 217180 472696
rect 179965 472638 217180 472640
rect 179965 472635 180031 472638
rect 217174 472636 217180 472638
rect 217244 472636 217250 472700
rect 55857 472562 55923 472565
rect 121821 472562 121887 472565
rect 55857 472560 121887 472562
rect 55857 472504 55862 472560
rect 55918 472504 121826 472560
rect 121882 472504 121887 472560
rect 55857 472502 121887 472504
rect 55857 472499 55923 472502
rect 121821 472499 121887 472502
rect 152641 472562 152707 472565
rect 212022 472562 212028 472564
rect 152641 472560 212028 472562
rect 152641 472504 152646 472560
rect 152702 472504 212028 472560
rect 152641 472502 212028 472504
rect 152641 472499 152707 472502
rect 212022 472500 212028 472502
rect 212092 472500 212098 472564
rect 256141 472562 256207 472565
rect 379462 472562 379468 472564
rect 256141 472560 379468 472562
rect 256141 472504 256146 472560
rect 256202 472504 379468 472560
rect 256141 472502 379468 472504
rect 256141 472499 256207 472502
rect 379462 472500 379468 472502
rect 379532 472500 379538 472564
rect 146017 471338 146083 471341
rect 204846 471338 204852 471340
rect 146017 471336 204852 471338
rect 146017 471280 146022 471336
rect 146078 471280 204852 471336
rect 146017 471278 204852 471280
rect 146017 471275 146083 471278
rect 204846 471276 204852 471278
rect 204916 471276 204922 471340
rect 583520 471324 584960 471564
rect 151721 471202 151787 471205
rect 215518 471202 215524 471204
rect 151721 471200 215524 471202
rect 151721 471144 151726 471200
rect 151782 471144 215524 471200
rect 151721 471142 215524 471144
rect 151721 471139 151787 471142
rect 215518 471140 215524 471142
rect 215588 471140 215594 471204
rect 234061 471202 234127 471205
rect 378726 471202 378732 471204
rect 234061 471200 378732 471202
rect 234061 471144 234066 471200
rect 234122 471144 378732 471200
rect 234061 471142 378732 471144
rect 234061 471139 234127 471142
rect 378726 471140 378732 471142
rect 378796 471140 378802 471204
rect 172697 470114 172763 470117
rect 206318 470114 206324 470116
rect 172697 470112 206324 470114
rect 172697 470056 172702 470112
rect 172758 470056 206324 470112
rect 172697 470054 206324 470056
rect 172697 470051 172763 470054
rect 206318 470052 206324 470054
rect 206388 470052 206394 470116
rect 44766 469916 44772 469980
rect 44836 469978 44842 469980
rect 124305 469978 124371 469981
rect 44836 469976 124371 469978
rect 44836 469920 124310 469976
rect 124366 469920 124371 469976
rect 44836 469918 124371 469920
rect 44836 469916 44842 469918
rect 124305 469915 124371 469918
rect 155953 469978 156019 469981
rect 211838 469978 211844 469980
rect 155953 469976 211844 469978
rect 155953 469920 155958 469976
rect 156014 469920 211844 469976
rect 155953 469918 211844 469920
rect 155953 469915 156019 469918
rect 211838 469916 211844 469918
rect 211908 469916 211914 469980
rect 44950 469780 44956 469844
rect 45020 469842 45026 469844
rect 128537 469842 128603 469845
rect 45020 469840 128603 469842
rect 45020 469784 128542 469840
rect 128598 469784 128603 469840
rect 45020 469782 128603 469784
rect 45020 469780 45026 469782
rect 128537 469779 128603 469782
rect 153285 469842 153351 469845
rect 212574 469842 212580 469844
rect 153285 469840 212580 469842
rect 153285 469784 153290 469840
rect 153346 469784 212580 469840
rect 153285 469782 212580 469784
rect 153285 469779 153351 469782
rect 212574 469780 212580 469782
rect 212644 469780 212650 469844
rect 263685 469842 263751 469845
rect 359590 469842 359596 469844
rect 263685 469840 359596 469842
rect 263685 469784 263690 469840
rect 263746 469784 359596 469840
rect 263685 469782 359596 469784
rect 263685 469779 263751 469782
rect 359590 469780 359596 469782
rect 359660 469780 359666 469844
rect 157425 468754 157491 468757
rect 209998 468754 210004 468756
rect 157425 468752 210004 468754
rect 157425 468696 157430 468752
rect 157486 468696 210004 468752
rect 157425 468694 210004 468696
rect 157425 468691 157491 468694
rect 209998 468692 210004 468694
rect 210068 468692 210074 468756
rect 150433 468618 150499 468621
rect 214598 468618 214604 468620
rect 150433 468616 214604 468618
rect 150433 468560 150438 468616
rect 150494 468560 214604 468616
rect 150433 468558 214604 468560
rect 150433 468555 150499 468558
rect 214598 468556 214604 468558
rect 214668 468556 214674 468620
rect 143625 468482 143691 468485
rect 211654 468482 211660 468484
rect 143625 468480 211660 468482
rect 143625 468424 143630 468480
rect 143686 468424 211660 468480
rect 143625 468422 211660 468424
rect 143625 468419 143691 468422
rect 211654 468420 211660 468422
rect 211724 468420 211730 468484
rect 230473 468482 230539 468485
rect 378910 468482 378916 468484
rect 230473 468480 378916 468482
rect 230473 468424 230478 468480
rect 230534 468424 378916 468480
rect 230473 468422 378916 468424
rect 230473 468419 230539 468422
rect 378910 468420 378916 468422
rect 378980 468420 378986 468484
rect 154573 467258 154639 467261
rect 207054 467258 207060 467260
rect 154573 467256 207060 467258
rect 154573 467200 154578 467256
rect 154634 467200 207060 467256
rect 154573 467198 207060 467200
rect 154573 467195 154639 467198
rect 207054 467196 207060 467198
rect 207124 467196 207130 467260
rect 147673 467122 147739 467125
rect 209078 467122 209084 467124
rect 147673 467120 209084 467122
rect 147673 467064 147678 467120
rect 147734 467064 209084 467120
rect 147673 467062 209084 467064
rect 147673 467059 147739 467062
rect 209078 467060 209084 467062
rect 209148 467060 209154 467124
rect 42609 466306 42675 466309
rect 70577 466306 70643 466309
rect 42609 466304 70643 466306
rect 42609 466248 42614 466304
rect 42670 466248 70582 466304
rect 70638 466248 70643 466304
rect 42609 466246 70643 466248
rect 42609 466243 42675 466246
rect 70577 466243 70643 466246
rect 187877 466306 187943 466309
rect 214925 466306 214991 466309
rect 187877 466304 214991 466306
rect 187877 466248 187882 466304
rect 187938 466248 214930 466304
rect 214986 466248 214991 466304
rect 187877 466246 214991 466248
rect 187877 466243 187943 466246
rect 214925 466243 214991 466246
rect 53465 466170 53531 466173
rect 85757 466170 85823 466173
rect 53465 466168 85823 466170
rect 53465 466112 53470 466168
rect 53526 466112 85762 466168
rect 85818 466112 85823 466168
rect 53465 466110 85823 466112
rect 53465 466107 53531 466110
rect 85757 466107 85823 466110
rect 169845 466170 169911 466173
rect 203190 466170 203196 466172
rect 169845 466168 203196 466170
rect 169845 466112 169850 466168
rect 169906 466112 203196 466168
rect 169845 466110 203196 466112
rect 169845 466107 169911 466110
rect 203190 466108 203196 466110
rect 203260 466108 203266 466172
rect 50797 466034 50863 466037
rect 84285 466034 84351 466037
rect 50797 466032 84351 466034
rect 50797 465976 50802 466032
rect 50858 465976 84290 466032
rect 84346 465976 84351 466032
rect 50797 465974 84351 465976
rect 50797 465971 50863 465974
rect 84285 465971 84351 465974
rect 160093 466034 160159 466037
rect 209037 466034 209103 466037
rect 160093 466032 209103 466034
rect 160093 465976 160098 466032
rect 160154 465976 209042 466032
rect 209098 465976 209103 466032
rect 160093 465974 209103 465976
rect 160093 465971 160159 465974
rect 209037 465971 209103 465974
rect 47894 465836 47900 465900
rect 47964 465898 47970 465900
rect 81525 465898 81591 465901
rect 47964 465896 81591 465898
rect 47964 465840 81530 465896
rect 81586 465840 81591 465896
rect 47964 465838 81591 465840
rect 47964 465836 47970 465838
rect 81525 465835 81591 465838
rect 161657 465898 161723 465901
rect 211981 465898 212047 465901
rect 161657 465896 212047 465898
rect 161657 465840 161662 465896
rect 161718 465840 211986 465896
rect 212042 465840 212047 465896
rect 161657 465838 212047 465840
rect 161657 465835 161723 465838
rect 211981 465835 212047 465838
rect 296805 465898 296871 465901
rect 377438 465898 377444 465900
rect 296805 465896 377444 465898
rect 296805 465840 296810 465896
rect 296866 465840 377444 465896
rect 296805 465838 377444 465840
rect 296805 465835 296871 465838
rect 377438 465836 377444 465838
rect 377508 465836 377514 465900
rect 57830 465700 57836 465764
rect 57900 465762 57906 465764
rect 102225 465762 102291 465765
rect 57900 465760 102291 465762
rect 57900 465704 102230 465760
rect 102286 465704 102291 465760
rect 57900 465702 102291 465704
rect 57900 465700 57906 465702
rect 102225 465699 102291 465702
rect 124213 465762 124279 465765
rect 196893 465762 196959 465765
rect 124213 465760 196959 465762
rect 124213 465704 124218 465760
rect 124274 465704 196898 465760
rect 196954 465704 196959 465760
rect 124213 465702 196959 465704
rect 124213 465699 124279 465702
rect 196893 465699 196959 465702
rect 229093 465762 229159 465765
rect 376150 465762 376156 465764
rect 229093 465760 376156 465762
rect 229093 465704 229098 465760
rect 229154 465704 376156 465760
rect 229093 465702 376156 465704
rect 229093 465699 229159 465702
rect 376150 465700 376156 465702
rect 376220 465700 376226 465764
rect 172605 464402 172671 464405
rect 207974 464402 207980 464404
rect 172605 464400 207980 464402
rect 172605 464344 172610 464400
rect 172666 464344 207980 464400
rect 172605 464342 207980 464344
rect 172605 464339 172671 464342
rect 207974 464340 207980 464342
rect 208044 464340 208050 464404
rect 52126 463388 52132 463452
rect 52196 463450 52202 463452
rect 70485 463450 70551 463453
rect 52196 463448 70551 463450
rect 52196 463392 70490 463448
rect 70546 463392 70551 463448
rect 52196 463390 70551 463392
rect 52196 463388 52202 463390
rect 70485 463387 70551 463390
rect 59077 463314 59143 463317
rect 91185 463314 91251 463317
rect 59077 463312 91251 463314
rect 59077 463256 59082 463312
rect 59138 463256 91190 463312
rect 91246 463256 91251 463312
rect 59077 463254 91251 463256
rect 59077 463251 59143 463254
rect 91185 463251 91251 463254
rect 186313 463314 186379 463317
rect 217358 463314 217364 463316
rect 186313 463312 217364 463314
rect 186313 463256 186318 463312
rect 186374 463256 217364 463312
rect 186313 463254 217364 463256
rect 186313 463251 186379 463254
rect 217358 463252 217364 463254
rect 217428 463252 217434 463316
rect 59997 463178 60063 463181
rect 92657 463178 92723 463181
rect 59997 463176 92723 463178
rect 59997 463120 60002 463176
rect 60058 463120 92662 463176
rect 92718 463120 92723 463176
rect 59997 463118 92723 463120
rect 59997 463115 60063 463118
rect 92657 463115 92723 463118
rect 171225 463178 171291 463181
rect 203006 463178 203012 463180
rect 171225 463176 203012 463178
rect 171225 463120 171230 463176
rect 171286 463120 203012 463176
rect 171225 463118 203012 463120
rect 171225 463115 171291 463118
rect 203006 463116 203012 463118
rect 203076 463116 203082 463180
rect 50981 463042 51047 463045
rect 93945 463042 94011 463045
rect 50981 463040 94011 463042
rect 50981 462984 50986 463040
rect 51042 462984 93950 463040
rect 94006 462984 94011 463040
rect 50981 462982 94011 462984
rect 50981 462979 51047 462982
rect 93945 462979 94011 462982
rect 146477 463042 146543 463045
rect 202270 463042 202276 463044
rect 146477 463040 202276 463042
rect 146477 462984 146482 463040
rect 146538 462984 202276 463040
rect 146477 462982 202276 462984
rect 146477 462979 146543 462982
rect 202270 462980 202276 462982
rect 202340 462980 202346 463044
rect 47710 462844 47716 462908
rect 47780 462906 47786 462908
rect 94037 462906 94103 462909
rect 47780 462904 94103 462906
rect 47780 462848 94042 462904
rect 94098 462848 94103 462904
rect 47780 462846 94103 462848
rect 47780 462844 47786 462846
rect 94037 462843 94103 462846
rect 146293 462906 146359 462909
rect 213126 462906 213132 462908
rect 146293 462904 213132 462906
rect 146293 462848 146298 462904
rect 146354 462848 213132 462904
rect 146293 462846 213132 462848
rect 146293 462843 146359 462846
rect 213126 462844 213132 462846
rect 213196 462844 213202 462908
rect 295517 462906 295583 462909
rect 376886 462906 376892 462908
rect 295517 462904 376892 462906
rect 295517 462848 295522 462904
rect 295578 462848 376892 462904
rect 295517 462846 376892 462848
rect 295517 462843 295583 462846
rect 376886 462844 376892 462846
rect 376956 462844 376962 462908
rect -960 462634 480 462724
rect 3601 462634 3667 462637
rect -960 462632 3667 462634
rect -960 462576 3606 462632
rect 3662 462576 3667 462632
rect -960 462574 3667 462576
rect -960 462484 480 462574
rect 3601 462571 3667 462574
rect 59118 461620 59124 461684
rect 59188 461682 59194 461684
rect 67909 461682 67975 461685
rect 59188 461680 67975 461682
rect 59188 461624 67914 461680
rect 67970 461624 67975 461680
rect 59188 461622 67975 461624
rect 59188 461620 59194 461622
rect 67909 461619 67975 461622
rect 179505 461682 179571 461685
rect 179638 461682 179644 461684
rect 179505 461680 179644 461682
rect 179505 461624 179510 461680
rect 179566 461624 179644 461680
rect 179505 461622 179644 461624
rect 179505 461619 179571 461622
rect 179638 461620 179644 461622
rect 179708 461620 179714 461684
rect 60222 461484 60228 461548
rect 60292 461546 60298 461548
rect 73245 461546 73311 461549
rect 60292 461544 73311 461546
rect 60292 461488 73250 461544
rect 73306 461488 73311 461544
rect 60292 461486 73311 461488
rect 60292 461484 60298 461486
rect 73245 461483 73311 461486
rect 266353 461546 266419 461549
rect 359774 461546 359780 461548
rect 266353 461544 359780 461546
rect 266353 461488 266358 461544
rect 266414 461488 359780 461544
rect 266353 461486 359780 461488
rect 266353 461483 266419 461486
rect 359774 461484 359780 461486
rect 359844 461484 359850 461548
rect 178309 461412 178375 461413
rect 178309 461408 178356 461412
rect 178420 461410 178426 461412
rect 178309 461352 178314 461408
rect 178309 461348 178356 461352
rect 178420 461350 178466 461410
rect 178420 461348 178426 461350
rect 178309 461347 178375 461348
rect 190913 461004 190979 461005
rect 338297 461004 338363 461005
rect 339769 461004 339835 461005
rect 350993 461004 351059 461005
rect 190862 461002 190868 461004
rect 190822 460942 190868 461002
rect 190932 461000 190979 461004
rect 338246 461002 338252 461004
rect 190974 460944 190979 461000
rect 190862 460940 190868 460942
rect 190932 460940 190979 460944
rect 338206 460942 338252 461002
rect 338316 461000 338363 461004
rect 339718 461002 339724 461004
rect 338358 460944 338363 461000
rect 338246 460940 338252 460942
rect 338316 460940 338363 460944
rect 339678 460942 339724 461002
rect 339788 461000 339835 461004
rect 350942 461002 350948 461004
rect 339830 460944 339835 461000
rect 339718 460940 339724 460942
rect 339788 460940 339835 460944
rect 350902 460942 350948 461002
rect 351012 461000 351059 461004
rect 351054 460944 351059 461000
rect 350942 460940 350948 460942
rect 351012 460940 351059 460944
rect 190913 460939 190979 460940
rect 338297 460939 338363 460940
rect 339769 460939 339835 460940
rect 350993 460939 351059 460940
rect 498193 461002 498259 461005
rect 499849 461004 499915 461005
rect 510889 461004 510955 461005
rect 498510 461002 498516 461004
rect 498193 461000 498516 461002
rect 498193 460944 498198 461000
rect 498254 460944 498516 461000
rect 498193 460942 498516 460944
rect 498193 460939 498259 460942
rect 498510 460940 498516 460942
rect 498580 460940 498586 461004
rect 499798 461002 499804 461004
rect 499758 460942 499804 461002
rect 499868 461000 499915 461004
rect 510838 461002 510844 461004
rect 499910 460944 499915 461000
rect 499798 460940 499804 460942
rect 499868 460940 499915 460944
rect 510798 460942 510844 461002
rect 510908 461000 510955 461004
rect 510950 460944 510955 461000
rect 510838 460940 510844 460942
rect 510908 460940 510955 460944
rect 499849 460939 499915 460940
rect 510889 460939 510955 460940
rect 48078 460804 48084 460868
rect 48148 460866 48154 460868
rect 69197 460866 69263 460869
rect 48148 460864 69263 460866
rect 48148 460808 69202 460864
rect 69258 460808 69263 460864
rect 48148 460806 69263 460808
rect 48148 460804 48154 460806
rect 69197 460803 69263 460806
rect 167177 460866 167243 460869
rect 202454 460866 202460 460868
rect 167177 460864 202460 460866
rect 167177 460808 167182 460864
rect 167238 460808 202460 460864
rect 167177 460806 202460 460808
rect 167177 460803 167243 460806
rect 202454 460804 202460 460806
rect 202524 460804 202530 460868
rect 46606 460668 46612 460732
rect 46676 460730 46682 460732
rect 67817 460730 67883 460733
rect 46676 460728 67883 460730
rect 46676 460672 67822 460728
rect 67878 460672 67883 460728
rect 46676 460670 67883 460672
rect 46676 460668 46682 460670
rect 67817 460667 67883 460670
rect 166993 460730 167059 460733
rect 205214 460730 205220 460732
rect 166993 460728 205220 460730
rect 166993 460672 166998 460728
rect 167054 460672 205220 460728
rect 166993 460670 205220 460672
rect 166993 460667 167059 460670
rect 205214 460668 205220 460670
rect 205284 460668 205290 460732
rect 55622 460532 55628 460596
rect 55692 460594 55698 460596
rect 77385 460594 77451 460597
rect 55692 460592 77451 460594
rect 55692 460536 77390 460592
rect 77446 460536 77451 460592
rect 55692 460534 77451 460536
rect 55692 460532 55698 460534
rect 77385 460531 77451 460534
rect 164325 460594 164391 460597
rect 215886 460594 215892 460596
rect 164325 460592 215892 460594
rect 164325 460536 164330 460592
rect 164386 460536 215892 460592
rect 164325 460534 215892 460536
rect 164325 460531 164391 460534
rect 215886 460532 215892 460534
rect 215956 460532 215962 460596
rect 51942 460396 51948 460460
rect 52012 460458 52018 460460
rect 74625 460458 74691 460461
rect 52012 460456 74691 460458
rect 52012 460400 74630 460456
rect 74686 460400 74691 460456
rect 52012 460398 74691 460400
rect 52012 460396 52018 460398
rect 74625 460395 74691 460398
rect 157333 460458 157399 460461
rect 218646 460458 218652 460460
rect 157333 460456 218652 460458
rect 157333 460400 157338 460456
rect 157394 460400 218652 460456
rect 157333 460398 218652 460400
rect 157333 460395 157399 460398
rect 218646 460396 218652 460398
rect 218716 460396 218722 460460
rect 51758 460260 51764 460324
rect 51828 460322 51834 460324
rect 75913 460322 75979 460325
rect 51828 460320 75979 460322
rect 51828 460264 75918 460320
rect 75974 460264 75979 460320
rect 51828 460262 75979 460264
rect 51828 460260 51834 460262
rect 75913 460259 75979 460262
rect 143717 460322 143783 460325
rect 205030 460322 205036 460324
rect 143717 460320 205036 460322
rect 143717 460264 143722 460320
rect 143778 460264 205036 460320
rect 143717 460262 205036 460264
rect 143717 460259 143783 460262
rect 205030 460260 205036 460262
rect 205100 460260 205106 460324
rect 295425 460322 295491 460325
rect 359958 460322 359964 460324
rect 295425 460320 359964 460322
rect 295425 460264 295430 460320
rect 295486 460264 359964 460320
rect 295425 460262 359964 460264
rect 295425 460259 295491 460262
rect 359958 460260 359964 460262
rect 360028 460260 360034 460324
rect 50654 460124 50660 460188
rect 50724 460186 50730 460188
rect 78673 460186 78739 460189
rect 50724 460184 78739 460186
rect 50724 460128 78678 460184
rect 78734 460128 78739 460184
rect 50724 460126 78739 460128
rect 50724 460124 50730 460126
rect 78673 460123 78739 460126
rect 153193 460186 153259 460189
rect 218830 460186 218836 460188
rect 153193 460184 218836 460186
rect 153193 460128 153198 460184
rect 153254 460128 218836 460184
rect 153193 460126 218836 460128
rect 153193 460123 153259 460126
rect 218830 460124 218836 460126
rect 218900 460124 218906 460188
rect 278773 460186 278839 460189
rect 377622 460186 377628 460188
rect 278773 460184 377628 460186
rect 278773 460128 278778 460184
rect 278834 460128 377628 460184
rect 278773 460126 377628 460128
rect 278773 460123 278839 460126
rect 377622 460124 377628 460126
rect 377692 460124 377698 460188
rect 53414 459988 53420 460052
rect 53484 460050 53490 460052
rect 74533 460050 74599 460053
rect 53484 460048 74599 460050
rect 53484 459992 74538 460048
rect 74594 459992 74599 460048
rect 53484 459990 74599 459992
rect 53484 459988 53490 459990
rect 74533 459987 74599 459990
rect 50470 459580 50476 459644
rect 50540 459642 50546 459644
rect 50705 459642 50771 459645
rect 50540 459640 50771 459642
rect 50540 459584 50710 459640
rect 50766 459584 50771 459640
rect 50540 459582 50771 459584
rect 50540 459580 50546 459582
rect 50705 459579 50771 459582
rect 53598 459580 53604 459644
rect 53668 459642 53674 459644
rect 53741 459642 53807 459645
rect 53668 459640 53807 459642
rect 53668 459584 53746 459640
rect 53802 459584 53807 459640
rect 53668 459582 53807 459584
rect 53668 459580 53674 459582
rect 53741 459579 53807 459582
rect 172513 459506 172579 459509
rect 200798 459506 200804 459508
rect 172513 459504 200804 459506
rect 172513 459448 172518 459504
rect 172574 459448 200804 459504
rect 172513 459446 200804 459448
rect 172513 459443 172579 459446
rect 200798 459444 200804 459446
rect 200868 459444 200874 459508
rect 168557 459370 168623 459373
rect 207749 459370 207815 459373
rect 168557 459368 207815 459370
rect 168557 459312 168562 459368
rect 168618 459312 207754 459368
rect 207810 459312 207815 459368
rect 168557 459310 207815 459312
rect 168557 459307 168623 459310
rect 207749 459307 207815 459310
rect 171133 459234 171199 459237
rect 214741 459234 214807 459237
rect 171133 459232 214807 459234
rect 171133 459176 171138 459232
rect 171194 459176 214746 459232
rect 214802 459176 214807 459232
rect 171133 459174 214807 459176
rect 171133 459171 171199 459174
rect 214741 459171 214807 459174
rect 58566 459036 58572 459100
rect 58636 459098 58642 459100
rect 67633 459098 67699 459101
rect 58636 459096 67699 459098
rect 58636 459040 67638 459096
rect 67694 459040 67699 459096
rect 58636 459038 67699 459040
rect 58636 459036 58642 459038
rect 67633 459035 67699 459038
rect 168373 459098 168439 459101
rect 213177 459098 213243 459101
rect 168373 459096 213243 459098
rect 168373 459040 168378 459096
rect 168434 459040 213182 459096
rect 213238 459040 213243 459096
rect 168373 459038 213243 459040
rect 168373 459035 168439 459038
rect 213177 459035 213243 459038
rect 58934 458900 58940 458964
rect 59004 458962 59010 458964
rect 69105 458962 69171 458965
rect 59004 458960 69171 458962
rect 59004 458904 69110 458960
rect 69166 458904 69171 458960
rect 59004 458902 69171 458904
rect 59004 458900 59010 458902
rect 69105 458899 69171 458902
rect 164233 458962 164299 458965
rect 218881 458962 218947 458965
rect 164233 458960 218947 458962
rect 164233 458904 164238 458960
rect 164294 458904 218886 458960
rect 218942 458904 218947 458960
rect 164233 458902 218947 458904
rect 164233 458899 164299 458902
rect 218881 458899 218947 458902
rect 223757 458962 223823 458965
rect 379094 458962 379100 458964
rect 223757 458960 379100 458962
rect 223757 458904 223762 458960
rect 223818 458904 379100 458960
rect 223757 458902 379100 458904
rect 223757 458899 223823 458902
rect 379094 458900 379100 458902
rect 379164 458900 379170 458964
rect 58750 458764 58756 458828
rect 58820 458826 58826 458828
rect 69013 458826 69079 458829
rect 58820 458824 69079 458826
rect 58820 458768 69018 458824
rect 69074 458768 69079 458824
rect 58820 458766 69079 458768
rect 58820 458764 58826 458766
rect 69013 458763 69079 458766
rect 125685 458826 125751 458829
rect 199142 458826 199148 458828
rect 125685 458824 199148 458826
rect 125685 458768 125690 458824
rect 125746 458768 199148 458824
rect 125685 458766 199148 458768
rect 125685 458763 125751 458766
rect 199142 458764 199148 458766
rect 199212 458764 199218 458828
rect 223573 458826 223639 458829
rect 379278 458826 379284 458828
rect 223573 458824 379284 458826
rect 223573 458768 223578 458824
rect 223634 458768 379284 458824
rect 223573 458766 379284 458768
rect 223573 458763 223639 458766
rect 379278 458764 379284 458766
rect 379348 458764 379354 458828
rect 580257 458146 580323 458149
rect 583520 458146 584960 458236
rect 580257 458144 584960 458146
rect 580257 458088 580262 458144
rect 580318 458088 584960 458144
rect 580257 458086 584960 458088
rect 580257 458083 580323 458086
rect 583520 457996 584960 458086
rect 205398 456860 205404 456924
rect 205468 456922 205474 456924
rect 205541 456922 205607 456925
rect 205468 456920 205607 456922
rect 205468 456864 205546 456920
rect 205602 456864 205607 456920
rect 205468 456862 205607 456864
rect 205468 456860 205474 456862
rect 205541 456859 205607 456862
rect 199009 454746 199075 454749
rect 358813 454746 358879 454749
rect 516593 454746 516659 454749
rect 196558 454744 199075 454746
rect 196558 454688 199014 454744
rect 199070 454688 199075 454744
rect 196558 454686 199075 454688
rect 196558 454190 196618 454686
rect 199009 454683 199075 454686
rect 356562 454744 358879 454746
rect 356562 454688 358818 454744
rect 358874 454688 358879 454744
rect 356562 454686 358879 454688
rect 356562 454190 356622 454686
rect 358813 454683 358879 454686
rect 516558 454744 516659 454746
rect 516558 454688 516598 454744
rect 516654 454688 516659 454744
rect 516558 454683 516659 454688
rect 516558 454202 516618 454683
rect 518893 454202 518959 454205
rect 516558 454200 518959 454202
rect 516558 454144 518898 454200
rect 518954 454144 518959 454200
rect 516558 454142 518959 454144
rect 518893 454139 518959 454142
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect 55673 415306 55739 415309
rect 56542 415306 56548 415308
rect 55673 415304 56548 415306
rect 55673 415248 55678 415304
rect 55734 415248 56548 415304
rect 55673 415246 56548 415248
rect 55673 415243 55739 415246
rect 56542 415244 56548 415246
rect 56612 415244 56618 415308
rect 56961 412314 57027 412317
rect 56961 412312 60062 412314
rect 56961 412256 56966 412312
rect 57022 412256 60062 412312
rect 56961 412254 60062 412256
rect 56961 412251 57027 412254
rect 60002 411894 60062 412254
rect 217961 411906 218027 411909
rect 219390 411906 220064 411924
rect 217961 411904 220064 411906
rect 217961 411848 217966 411904
rect 218022 411864 220064 411904
rect 377029 411906 377095 411909
rect 379470 411906 380052 411924
rect 377029 411904 380052 411906
rect 218022 411848 219450 411864
rect 217961 411846 219450 411848
rect 377029 411848 377034 411904
rect 377090 411864 380052 411904
rect 377090 411848 379530 411864
rect 377029 411846 379530 411848
rect 217961 411843 218027 411846
rect 377029 411843 377095 411846
rect 216949 411362 217015 411365
rect 217961 411362 218027 411365
rect 216949 411360 218027 411362
rect 216949 411304 216954 411360
rect 217010 411304 217966 411360
rect 218022 411304 218027 411360
rect 216949 411302 218027 411304
rect 216949 411299 217015 411302
rect 217961 411299 218027 411302
rect 217777 410954 217843 410957
rect 219390 410954 220064 410972
rect 217777 410952 220064 410954
rect -960 410546 480 410636
rect 2957 410546 3023 410549
rect -960 410544 3023 410546
rect -960 410488 2962 410544
rect 3018 410488 3023 410544
rect -960 410486 3023 410488
rect -960 410396 480 410486
rect 2957 410483 3023 410486
rect 57053 410410 57119 410413
rect 60002 410410 60062 410942
rect 217777 410896 217782 410952
rect 217838 410912 220064 410952
rect 377213 410954 377279 410957
rect 377765 410954 377831 410957
rect 379470 410954 380052 410972
rect 377213 410952 380052 410954
rect 217838 410896 219450 410912
rect 217777 410894 219450 410896
rect 377213 410896 377218 410952
rect 377274 410896 377770 410952
rect 377826 410912 380052 410952
rect 377826 410896 379530 410912
rect 377213 410894 379530 410896
rect 217777 410891 217843 410894
rect 377213 410891 377279 410894
rect 377765 410891 377831 410894
rect 57053 410408 60062 410410
rect 57053 410352 57058 410408
rect 57114 410352 60062 410408
rect 57053 410350 60062 410352
rect 57053 410347 57119 410350
rect 217041 410002 217107 410005
rect 217777 410002 217843 410005
rect 217041 410000 217843 410002
rect 217041 409944 217046 410000
rect 217102 409944 217782 410000
rect 217838 409944 217843 410000
rect 217041 409942 217843 409944
rect 217041 409939 217107 409942
rect 217777 409939 217843 409942
rect 216673 408778 216739 408781
rect 219390 408778 220064 408796
rect 216673 408776 220064 408778
rect 57053 408642 57119 408645
rect 60002 408642 60062 408766
rect 216673 408720 216678 408776
rect 216734 408736 220064 408776
rect 377213 408778 377279 408781
rect 377857 408778 377923 408781
rect 379470 408778 380052 408796
rect 377213 408776 380052 408778
rect 216734 408720 219450 408736
rect 216673 408718 219450 408720
rect 377213 408720 377218 408776
rect 377274 408720 377862 408776
rect 377918 408736 380052 408776
rect 377918 408720 379530 408736
rect 377213 408718 379530 408720
rect 216673 408715 216739 408718
rect 377213 408715 377279 408718
rect 377857 408715 377923 408718
rect 57053 408640 60062 408642
rect 57053 408584 57058 408640
rect 57114 408584 60062 408640
rect 57053 408582 60062 408584
rect 57053 408579 57119 408582
rect 56542 407764 56548 407828
rect 56612 407826 56618 407828
rect 59353 407826 59419 407829
rect 56612 407824 59419 407826
rect 56612 407768 59358 407824
rect 59414 407768 59419 407824
rect 56612 407766 59419 407768
rect 56612 407764 56618 407766
rect 59353 407763 59419 407766
rect 56961 407418 57027 407421
rect 60002 407418 60062 407814
rect 207054 407764 207060 407828
rect 207124 407826 207130 407828
rect 208301 407826 208367 407829
rect 207124 407824 208367 407826
rect 207124 407768 208306 407824
rect 208362 407768 208367 407824
rect 207124 407766 208367 407768
rect 207124 407764 207130 407766
rect 208301 407763 208367 407766
rect 216673 407826 216739 407829
rect 219390 407826 220064 407844
rect 216673 407824 220064 407826
rect 216673 407768 216678 407824
rect 216734 407784 220064 407824
rect 216734 407768 219450 407784
rect 216673 407766 219450 407768
rect 216673 407763 216739 407766
rect 358118 407764 358124 407828
rect 358188 407826 358194 407828
rect 358629 407826 358695 407829
rect 358188 407824 358695 407826
rect 358188 407768 358634 407824
rect 358690 407768 358695 407824
rect 358188 407766 358695 407768
rect 358188 407764 358194 407766
rect 358629 407763 358695 407766
rect 377121 407826 377187 407829
rect 377489 407826 377555 407829
rect 379470 407826 380052 407844
rect 377121 407824 380052 407826
rect 377121 407768 377126 407824
rect 377182 407768 377494 407824
rect 377550 407784 380052 407824
rect 377550 407768 379530 407784
rect 377121 407766 379530 407768
rect 377121 407763 377187 407766
rect 377489 407763 377555 407766
rect 56961 407416 60062 407418
rect 56961 407360 56966 407416
rect 57022 407360 60062 407416
rect 56961 407358 60062 407360
rect 56961 407355 57027 407358
rect 216857 406058 216923 406061
rect 219390 406058 220064 406076
rect 216857 406056 220064 406058
rect 57053 405786 57119 405789
rect 60002 405786 60062 406046
rect 216857 406000 216862 406056
rect 216918 406016 220064 406056
rect 377213 406058 377279 406061
rect 379470 406058 380052 406076
rect 377213 406056 380052 406058
rect 216918 406000 219450 406016
rect 216857 405998 219450 406000
rect 377213 406000 377218 406056
rect 377274 406016 380052 406056
rect 377274 406000 379530 406016
rect 377213 405998 379530 406000
rect 216857 405995 216923 405998
rect 377213 405995 377279 405998
rect 57053 405784 60062 405786
rect 57053 405728 57058 405784
rect 57114 405728 60062 405784
rect 57053 405726 60062 405728
rect 57053 405723 57119 405726
rect 217869 404970 217935 404973
rect 219390 404970 220064 404988
rect 217869 404968 220064 404970
rect 57053 404426 57119 404429
rect 60002 404426 60062 404958
rect 217869 404912 217874 404968
rect 217930 404928 220064 404968
rect 377581 404970 377647 404973
rect 379470 404970 380052 404988
rect 377581 404968 380052 404970
rect 217930 404912 219450 404928
rect 217869 404910 219450 404912
rect 377581 404912 377586 404968
rect 377642 404928 380052 404968
rect 580257 404970 580323 404973
rect 583520 404970 584960 405060
rect 580257 404968 584960 404970
rect 377642 404912 379530 404928
rect 377581 404910 379530 404912
rect 580257 404912 580262 404968
rect 580318 404912 584960 404968
rect 580257 404910 584960 404912
rect 217869 404907 217935 404910
rect 377581 404907 377647 404910
rect 580257 404907 580323 404910
rect 583520 404820 584960 404910
rect 57053 404424 60062 404426
rect 57053 404368 57058 404424
rect 57114 404368 60062 404424
rect 57053 404366 60062 404368
rect 57053 404363 57119 404366
rect 217685 404290 217751 404293
rect 217869 404290 217935 404293
rect 217685 404288 217935 404290
rect 217685 404232 217690 404288
rect 217746 404232 217874 404288
rect 217930 404232 217935 404288
rect 217685 404230 217935 404232
rect 217685 404227 217751 404230
rect 217869 404227 217935 404230
rect 217869 403202 217935 403205
rect 219390 403202 220064 403220
rect 217869 403200 220064 403202
rect 56961 403066 57027 403069
rect 60002 403066 60062 403190
rect 217869 403144 217874 403200
rect 217930 403160 220064 403200
rect 377673 403202 377739 403205
rect 379470 403202 380052 403220
rect 377673 403200 380052 403202
rect 217930 403144 219450 403160
rect 217869 403142 219450 403144
rect 377673 403144 377678 403200
rect 377734 403160 380052 403200
rect 377734 403144 379530 403160
rect 377673 403142 379530 403144
rect 217869 403139 217935 403142
rect 377673 403139 377739 403142
rect 56961 403064 60062 403066
rect 56961 403008 56966 403064
rect 57022 403008 60062 403064
rect 56961 403006 60062 403008
rect 56961 403003 57027 403006
rect -960 397340 480 397580
rect 198089 394634 198155 394637
rect 198774 394634 198780 394636
rect 198089 394632 198780 394634
rect 198089 394576 198094 394632
rect 198150 394576 198780 394632
rect 198089 394574 198780 394576
rect 198089 394571 198155 394574
rect 198774 394572 198780 394574
rect 198844 394572 198850 394636
rect 196558 394090 196618 394350
rect 199653 394090 199719 394093
rect 196558 394088 199719 394090
rect 196558 394032 199658 394088
rect 199714 394032 199719 394088
rect 196558 394030 199719 394032
rect 199653 394027 199719 394030
rect 356562 393818 356622 394350
rect 360009 393818 360075 393821
rect 356562 393816 360075 393818
rect 356562 393760 360014 393816
rect 360070 393760 360075 393816
rect 356562 393758 360075 393760
rect 516558 393818 516618 394350
rect 518985 393818 519051 393821
rect 516558 393816 519051 393818
rect 516558 393760 518990 393816
rect 519046 393760 519051 393816
rect 516558 393758 519051 393760
rect 360009 393755 360075 393758
rect 518985 393755 519051 393758
rect 196558 392186 196618 392718
rect 199326 392186 199332 392188
rect 196558 392126 199332 392186
rect 199326 392124 199332 392126
rect 199396 392124 199402 392188
rect 356562 392186 356622 392718
rect 359917 392186 359983 392189
rect 356562 392184 359983 392186
rect 356562 392128 359922 392184
rect 359978 392128 359983 392184
rect 356562 392126 359983 392128
rect 516558 392186 516618 392718
rect 519169 392186 519235 392189
rect 516558 392184 519235 392186
rect 516558 392128 519174 392184
rect 519230 392128 519235 392184
rect 516558 392126 519235 392128
rect 359917 392123 359983 392126
rect 519169 392123 519235 392126
rect 198273 392050 198339 392053
rect 198774 392050 198780 392052
rect 198273 392048 198780 392050
rect 198273 391992 198278 392048
rect 198334 391992 198780 392048
rect 198273 391990 198780 391992
rect 198273 391987 198339 391990
rect 198774 391988 198780 391990
rect 198844 391988 198850 392052
rect 583520 391628 584960 391868
rect 196558 390826 196618 391358
rect 199193 390826 199259 390829
rect 199561 390826 199627 390829
rect 196558 390824 199627 390826
rect 196558 390768 199198 390824
rect 199254 390768 199566 390824
rect 199622 390768 199627 390824
rect 196558 390766 199627 390768
rect 356562 390826 356622 391358
rect 359825 390826 359891 390829
rect 356562 390824 359891 390826
rect 356562 390768 359830 390824
rect 359886 390768 359891 390824
rect 356562 390766 359891 390768
rect 516558 390826 516618 391358
rect 519261 390826 519327 390829
rect 516558 390824 519327 390826
rect 516558 390768 519266 390824
rect 519322 390768 519327 390824
rect 516558 390766 519327 390768
rect 199193 390763 199259 390766
rect 199561 390763 199627 390766
rect 359825 390763 359891 390766
rect 519261 390763 519327 390766
rect 198181 390690 198247 390693
rect 199142 390690 199148 390692
rect 198181 390688 199148 390690
rect 198181 390632 198186 390688
rect 198242 390632 199148 390688
rect 198181 390630 199148 390632
rect 198181 390627 198247 390630
rect 199142 390628 199148 390630
rect 199212 390628 199218 390692
rect 196558 389194 196618 389862
rect 356562 389330 356622 389862
rect 359089 389330 359155 389333
rect 356562 389328 359155 389330
rect 356562 389272 359094 389328
rect 359150 389272 359155 389328
rect 356562 389270 359155 389272
rect 516558 389330 516618 389862
rect 519353 389330 519419 389333
rect 516558 389328 519419 389330
rect 516558 389272 519358 389328
rect 519414 389272 519419 389328
rect 516558 389270 519419 389272
rect 359089 389267 359155 389270
rect 519353 389267 519419 389270
rect 196558 389134 199210 389194
rect 199150 389060 199210 389134
rect 199142 388996 199148 389060
rect 199212 388996 199218 389060
rect 196558 388514 196618 388638
rect 198958 388514 198964 388516
rect 196558 388454 198964 388514
rect 198958 388452 198964 388454
rect 199028 388514 199034 388516
rect 199653 388514 199719 388517
rect 199028 388512 199719 388514
rect 199028 388456 199658 388512
rect 199714 388456 199719 388512
rect 199028 388454 199719 388456
rect 199028 388452 199034 388454
rect 199653 388451 199719 388454
rect 356562 388106 356622 388638
rect 360101 388106 360167 388109
rect 356562 388104 360167 388106
rect 356562 388048 360106 388104
rect 360162 388048 360167 388104
rect 356562 388046 360167 388048
rect 516558 388106 516618 388638
rect 519077 388106 519143 388109
rect 516558 388104 519143 388106
rect 516558 388048 519082 388104
rect 519138 388048 519143 388104
rect 516558 388046 519143 388048
rect 360101 388043 360167 388046
rect 519077 388043 519143 388046
rect 56961 384978 57027 384981
rect 216673 384978 216739 384981
rect 219390 384978 220064 384996
rect 56961 384976 60062 384978
rect 56961 384920 56966 384976
rect 57022 384920 60062 384976
rect 56961 384918 60062 384920
rect 216673 384976 220064 384978
rect 216673 384920 216678 384976
rect 216734 384936 220064 384976
rect 376937 384978 377003 384981
rect 379470 384978 380052 384996
rect 376937 384976 380052 384978
rect 216734 384920 219450 384936
rect 216673 384918 219450 384920
rect 376937 384920 376942 384976
rect 376998 384936 380052 384976
rect 376998 384920 379530 384936
rect 376937 384918 379530 384920
rect 56961 384915 57027 384918
rect 216673 384915 216739 384918
rect 376937 384915 377003 384918
rect -960 384284 480 384524
rect 56869 383346 56935 383349
rect 59494 383346 60032 383364
rect 56869 383344 60032 383346
rect 56869 383288 56874 383344
rect 56930 383304 60032 383344
rect 216673 383346 216739 383349
rect 219390 383346 220064 383364
rect 216673 383344 220064 383346
rect 56930 383288 59554 383304
rect 56869 383286 59554 383288
rect 216673 383288 216678 383344
rect 216734 383304 220064 383344
rect 376937 383346 377003 383349
rect 379470 383346 380052 383364
rect 376937 383344 380052 383346
rect 216734 383288 219450 383304
rect 216673 383286 219450 383288
rect 376937 383288 376942 383344
rect 376998 383304 380052 383344
rect 376998 383288 379530 383304
rect 376937 383286 379530 383288
rect 56869 383283 56935 383286
rect 216673 383283 216739 383286
rect 376937 383283 377003 383286
rect 57145 383074 57211 383077
rect 216857 383074 216923 383077
rect 219390 383074 220064 383092
rect 57145 383072 60062 383074
rect 57145 383016 57150 383072
rect 57206 383016 60062 383072
rect 57145 383014 60062 383016
rect 216857 383072 220064 383074
rect 216857 383016 216862 383072
rect 216918 383032 220064 383072
rect 376845 383074 376911 383077
rect 379470 383074 380052 383092
rect 376845 383072 380052 383074
rect 216918 383016 219450 383032
rect 216857 383014 219450 383016
rect 376845 383016 376850 383072
rect 376906 383032 380052 383072
rect 376906 383016 379530 383032
rect 376845 383014 379530 383016
rect 57145 383011 57211 383014
rect 216857 383011 216923 383014
rect 376845 383011 376911 383014
rect 212022 382332 212028 382396
rect 212092 382394 212098 382396
rect 212441 382394 212507 382397
rect 212092 382392 212507 382394
rect 212092 382336 212446 382392
rect 212502 382336 212507 382392
rect 212092 382334 212507 382336
rect 212092 382332 212098 382334
rect 212441 382331 212507 382334
rect 580441 378450 580507 378453
rect 583520 378450 584960 378540
rect 580441 378448 584960 378450
rect 580441 378392 580446 378448
rect 580502 378392 584960 378448
rect 580441 378390 584960 378392
rect 580441 378387 580507 378390
rect 583520 378300 584960 378390
rect 51758 375260 51764 375324
rect 51828 375322 51834 375324
rect 52361 375322 52427 375325
rect 51828 375320 52427 375322
rect 51828 375264 52366 375320
rect 52422 375264 52427 375320
rect 51828 375262 52427 375264
rect 51828 375260 51834 375262
rect 52361 375259 52427 375262
rect 53230 375260 53236 375324
rect 53300 375322 53306 375324
rect 53557 375322 53623 375325
rect 55489 375324 55555 375325
rect 55438 375322 55444 375324
rect 53300 375320 53623 375322
rect 53300 375264 53562 375320
rect 53618 375264 53623 375320
rect 53300 375262 53623 375264
rect 55398 375262 55444 375322
rect 55508 375320 55555 375324
rect 55550 375264 55555 375320
rect 53300 375260 53306 375262
rect 53557 375259 53623 375262
rect 55438 375260 55444 375262
rect 55508 375260 55555 375264
rect 200982 375260 200988 375324
rect 201052 375322 201058 375324
rect 201401 375322 201467 375325
rect 201052 375320 201467 375322
rect 201052 375264 201406 375320
rect 201462 375264 201467 375320
rect 201052 375262 201467 375264
rect 201052 375260 201058 375262
rect 55489 375259 55555 375260
rect 201401 375259 201467 375262
rect 202638 375260 202644 375324
rect 202708 375322 202714 375324
rect 202781 375322 202847 375325
rect 202708 375320 202847 375322
rect 202708 375264 202786 375320
rect 202842 375264 202847 375320
rect 202708 375262 202847 375264
rect 202708 375260 202714 375262
rect 202781 375259 202847 375262
rect 206502 375260 206508 375324
rect 206572 375322 206578 375324
rect 206829 375322 206895 375325
rect 206572 375320 206895 375322
rect 206572 375264 206834 375320
rect 206890 375264 206895 375320
rect 206572 375262 206895 375264
rect 206572 375260 206578 375262
rect 206829 375259 206895 375262
rect 209814 375260 209820 375324
rect 209884 375322 209890 375324
rect 211061 375322 211127 375325
rect 209884 375320 211127 375322
rect 209884 375264 211066 375320
rect 211122 375264 211127 375320
rect 209884 375262 211127 375264
rect 209884 375260 209890 375262
rect 211061 375259 211127 375262
rect 211838 375260 211844 375324
rect 211908 375322 211914 375324
rect 212349 375322 212415 375325
rect 211908 375320 212415 375322
rect 211908 375264 212354 375320
rect 212410 375264 212415 375320
rect 211908 375262 212415 375264
rect 211908 375260 211914 375262
rect 212349 375259 212415 375262
rect 216765 375322 216831 375325
rect 217869 375322 217935 375325
rect 216765 375320 217935 375322
rect 216765 375264 216770 375320
rect 216826 375264 217874 375320
rect 217930 375264 217935 375320
rect 216765 375262 217935 375264
rect 216765 375259 216831 375262
rect 217869 375259 217935 375262
rect 47485 375050 47551 375053
rect 216949 375050 217015 375053
rect 244733 375052 244799 375053
rect 270493 375052 270559 375053
rect 283005 375052 283071 375053
rect 244733 375050 244780 375052
rect 47485 375048 217015 375050
rect 47485 374992 47490 375048
rect 47546 374992 216954 375048
rect 217010 374992 217015 375048
rect 47485 374990 217015 374992
rect 244688 375048 244780 375050
rect 244688 374992 244738 375048
rect 244688 374990 244780 374992
rect 47485 374987 47551 374990
rect 216949 374987 217015 374990
rect 244733 374988 244780 374990
rect 244844 374988 244850 375052
rect 270493 375050 270540 375052
rect 270448 375048 270540 375050
rect 270448 374992 270498 375048
rect 270448 374990 270540 374992
rect 270493 374988 270540 374990
rect 270604 374988 270610 375052
rect 283005 375050 283052 375052
rect 282960 375048 283052 375050
rect 282960 374992 283010 375048
rect 282960 374990 283052 374992
rect 283005 374988 283052 374990
rect 283116 374988 283122 375052
rect 311801 375050 311867 375053
rect 407757 375052 407823 375053
rect 425053 375052 425119 375053
rect 440325 375052 440391 375053
rect 443085 375052 443151 375053
rect 315246 375050 315252 375052
rect 311801 375048 315252 375050
rect 311801 374992 311806 375048
rect 311862 374992 315252 375048
rect 311801 374990 315252 374992
rect 244733 374987 244799 374988
rect 270493 374987 270559 374988
rect 283005 374987 283071 374988
rect 311801 374987 311867 374990
rect 315246 374988 315252 374990
rect 315316 374988 315322 375052
rect 407757 375050 407804 375052
rect 407712 375048 407804 375050
rect 407712 374992 407762 375048
rect 407712 374990 407804 374992
rect 407757 374988 407804 374990
rect 407868 374988 407874 375052
rect 425053 375050 425100 375052
rect 425008 375048 425100 375050
rect 425008 374992 425058 375048
rect 425008 374990 425100 374992
rect 425053 374988 425100 374990
rect 425164 374988 425170 375052
rect 440325 375050 440372 375052
rect 440280 375048 440372 375050
rect 440280 374992 440330 375048
rect 440280 374990 440372 374992
rect 440325 374988 440372 374990
rect 440436 374988 440442 375052
rect 443085 375050 443132 375052
rect 443040 375048 443132 375050
rect 443040 374992 443090 375048
rect 443040 374990 443132 374992
rect 443085 374988 443132 374990
rect 443196 374988 443202 375052
rect 407757 374987 407823 374988
rect 425053 374987 425119 374988
rect 440325 374987 440391 374988
rect 443085 374987 443151 374988
rect 52453 374914 52519 374917
rect 216765 374914 216831 374917
rect 52453 374912 216831 374914
rect 52453 374856 52458 374912
rect 52514 374856 216770 374912
rect 216826 374856 216831 374912
rect 52453 374854 216831 374856
rect 52453 374851 52519 374854
rect 216765 374851 216831 374854
rect 404169 374780 404235 374781
rect 404169 374778 404214 374780
rect 404122 374776 404214 374778
rect 404122 374720 404174 374776
rect 404122 374718 404214 374720
rect 404169 374716 404214 374718
rect 404278 374716 404284 374780
rect 404169 374715 404235 374716
rect 158529 374644 158595 374645
rect 165981 374644 166047 374645
rect 158478 374580 158484 374644
rect 158548 374642 158595 374644
rect 158548 374640 158640 374642
rect 158590 374584 158640 374640
rect 158548 374582 158640 374584
rect 158548 374580 158595 374582
rect 165944 374580 165950 374644
rect 166014 374642 166047 374644
rect 195881 374642 195947 374645
rect 212901 374642 212967 374645
rect 320909 374644 320975 374645
rect 410701 374644 410767 374645
rect 450997 374644 451063 374645
rect 320909 374642 320918 374644
rect 166014 374640 166106 374642
rect 166042 374584 166106 374640
rect 166014 374582 166106 374584
rect 195881 374640 212967 374642
rect 195881 374584 195886 374640
rect 195942 374584 212906 374640
rect 212962 374584 212967 374640
rect 195881 374582 212967 374584
rect 320826 374640 320918 374642
rect 320826 374584 320914 374640
rect 320826 374582 320918 374584
rect 166014 374580 166047 374582
rect 158529 374579 158595 374580
rect 165981 374579 166047 374580
rect 195881 374579 195947 374582
rect 212901 374579 212967 374582
rect 320909 374580 320918 374582
rect 320982 374580 320988 374644
rect 359958 374580 359964 374644
rect 360028 374642 360034 374644
rect 410701 374642 410742 374644
rect 360028 374582 369870 374642
rect 410650 374640 410742 374642
rect 410650 374584 410706 374640
rect 410650 374582 410742 374584
rect 360028 374580 360034 374582
rect 320909 374579 320975 374580
rect 105445 374508 105511 374509
rect 116025 374508 116091 374509
rect 140957 374508 141023 374509
rect 143533 374508 143599 374509
rect 156505 374508 156571 374509
rect 160921 374508 160987 374509
rect 163405 374508 163471 374509
rect 244273 374508 244339 374509
rect 105445 374506 105492 374508
rect 105400 374504 105492 374506
rect 105400 374448 105450 374504
rect 105400 374446 105492 374448
rect 105445 374444 105492 374446
rect 105556 374444 105562 374508
rect 116025 374506 116038 374508
rect 115946 374504 116038 374506
rect 115946 374448 116030 374504
rect 115946 374446 116038 374448
rect 116025 374444 116038 374446
rect 116102 374444 116108 374508
rect 140920 374444 140926 374508
rect 140990 374506 141023 374508
rect 140990 374504 141082 374506
rect 141018 374448 141082 374504
rect 140990 374446 141082 374448
rect 140990 374444 141023 374446
rect 143504 374444 143510 374508
rect 143574 374506 143599 374508
rect 143574 374504 143666 374506
rect 143594 374448 143666 374504
rect 143574 374446 143666 374448
rect 143574 374444 143599 374446
rect 156454 374444 156460 374508
rect 156524 374506 156571 374508
rect 156524 374504 156616 374506
rect 156566 374448 156616 374504
rect 156524 374446 156616 374448
rect 156524 374444 156571 374446
rect 160912 374444 160918 374508
rect 160982 374506 160988 374508
rect 160982 374446 161074 374506
rect 160982 374444 160988 374446
rect 163360 374444 163366 374508
rect 163430 374506 163471 374508
rect 163430 374504 163522 374506
rect 163466 374448 163522 374504
rect 163430 374446 163522 374448
rect 163430 374444 163471 374446
rect 244222 374444 244228 374508
rect 244292 374506 244339 374508
rect 247585 374508 247651 374509
rect 253473 374508 253539 374509
rect 247585 374506 247614 374508
rect 244292 374504 244384 374506
rect 244334 374448 244384 374504
rect 244292 374446 244384 374448
rect 247522 374504 247614 374506
rect 247522 374448 247590 374504
rect 247522 374446 247614 374448
rect 244292 374444 244339 374446
rect 105445 374443 105511 374444
rect 116025 374443 116091 374444
rect 140957 374443 141023 374444
rect 143533 374443 143599 374444
rect 156505 374443 156571 374444
rect 160921 374443 160987 374444
rect 163405 374443 163471 374444
rect 244273 374443 244339 374444
rect 247585 374444 247614 374446
rect 247678 374444 247684 374508
rect 253456 374444 253462 374508
rect 253526 374506 253539 374508
rect 265249 374508 265315 374509
rect 265249 374506 265294 374508
rect 253526 374504 253618 374506
rect 253534 374448 253618 374504
rect 253526 374446 253618 374448
rect 265202 374504 265294 374506
rect 265202 374448 265254 374504
rect 265202 374446 265294 374448
rect 253526 374444 253539 374446
rect 247585 374443 247651 374444
rect 253473 374443 253539 374444
rect 265249 374444 265294 374446
rect 265358 374444 265364 374508
rect 265249 374443 265315 374444
rect 146201 374372 146267 374373
rect 148961 374372 149027 374373
rect 146150 374308 146156 374372
rect 146220 374370 146267 374372
rect 146220 374368 146312 374370
rect 146262 374312 146312 374368
rect 146220 374310 146312 374312
rect 146220 374308 146267 374310
rect 148910 374308 148916 374372
rect 148980 374370 149027 374372
rect 215477 374370 215543 374373
rect 262254 374370 262260 374372
rect 148980 374368 149072 374370
rect 149022 374312 149072 374368
rect 148980 374310 149072 374312
rect 215477 374368 262260 374370
rect 215477 374312 215482 374368
rect 215538 374312 262260 374368
rect 215477 374310 262260 374312
rect 148980 374308 149027 374310
rect 146201 374307 146267 374308
rect 148961 374307 149027 374308
rect 215477 374307 215543 374310
rect 262254 374308 262260 374310
rect 262324 374308 262330 374372
rect 218237 374234 218303 374237
rect 222101 374234 222167 374237
rect 218237 374232 222167 374234
rect 218237 374176 218242 374232
rect 218298 374176 222106 374232
rect 222162 374176 222167 374232
rect 218237 374174 222167 374176
rect 218237 374171 218303 374174
rect 222101 374171 222167 374174
rect 270309 374234 270375 374237
rect 273846 374234 273852 374236
rect 270309 374232 273852 374234
rect 270309 374176 270314 374232
rect 270370 374176 273852 374232
rect 270309 374174 273852 374176
rect 270309 374171 270375 374174
rect 273846 374172 273852 374174
rect 273916 374172 273922 374236
rect 139209 374100 139275 374101
rect 139158 374036 139164 374100
rect 139228 374098 139275 374100
rect 219617 374098 219683 374101
rect 222009 374098 222075 374101
rect 139228 374096 139320 374098
rect 139270 374040 139320 374096
rect 139228 374038 139320 374040
rect 219617 374096 222075 374098
rect 219617 374040 219622 374096
rect 219678 374040 222014 374096
rect 222070 374040 222075 374096
rect 219617 374038 222075 374040
rect 139228 374036 139275 374038
rect 139209 374035 139275 374036
rect 219617 374035 219683 374038
rect 222009 374035 222075 374038
rect 270217 374098 270283 374101
rect 271270 374098 271276 374100
rect 270217 374096 271276 374098
rect 270217 374040 270222 374096
rect 270278 374040 271276 374096
rect 270217 374038 271276 374040
rect 270217 374035 270283 374038
rect 271270 374036 271276 374038
rect 271340 374036 271346 374100
rect 369810 374098 369870 374582
rect 410701 374580 410742 374582
rect 410806 374580 410812 374644
rect 450992 374642 450998 374644
rect 450906 374582 450998 374642
rect 450992 374580 450998 374582
rect 451062 374580 451068 374644
rect 410701 374579 410767 374580
rect 450997 374579 451063 374580
rect 433609 374508 433675 374509
rect 433584 374444 433590 374508
rect 433654 374506 433675 374508
rect 436001 374508 436067 374509
rect 438485 374508 438551 374509
rect 436001 374506 436038 374508
rect 433654 374504 433746 374506
rect 433670 374448 433746 374504
rect 433654 374446 433746 374448
rect 435946 374504 436038 374506
rect 435946 374448 436006 374504
rect 435946 374446 436038 374448
rect 433654 374444 433675 374446
rect 433609 374443 433675 374444
rect 436001 374444 436038 374446
rect 436102 374444 436108 374508
rect 438480 374506 438486 374508
rect 438394 374446 438486 374506
rect 438480 374444 438486 374446
rect 438550 374444 438556 374508
rect 436001 374443 436067 374444
rect 438485 374443 438551 374444
rect 373073 374098 373139 374101
rect 429142 374098 429148 374100
rect 369810 374096 429148 374098
rect 369810 374040 373078 374096
rect 373134 374040 429148 374096
rect 369810 374038 429148 374040
rect 373073 374035 373139 374038
rect 429142 374036 429148 374038
rect 429212 374036 429218 374100
rect 42149 373962 42215 373965
rect 199142 373962 199148 373964
rect 42149 373960 199148 373962
rect 42149 373904 42154 373960
rect 42210 373904 199148 373960
rect 42149 373902 199148 373904
rect 42149 373899 42215 373902
rect 199142 373900 199148 373902
rect 199212 373900 199218 373964
rect 205449 373962 205515 373965
rect 279182 373962 279188 373964
rect 205449 373960 279188 373962
rect 205449 373904 205454 373960
rect 205510 373904 279188 373960
rect 205449 373902 279188 373904
rect 205449 373899 205515 373902
rect 279182 373900 279188 373902
rect 279252 373900 279258 373964
rect 377622 373900 377628 373964
rect 377692 373962 377698 373964
rect 475326 373962 475332 373964
rect 377692 373902 475332 373962
rect 377692 373900 377698 373902
rect 475326 373900 475332 373902
rect 475396 373900 475402 373964
rect 43253 373826 43319 373829
rect 199326 373826 199332 373828
rect 43253 373824 199332 373826
rect 43253 373768 43258 373824
rect 43314 373768 199332 373824
rect 43253 373766 199332 373768
rect 43253 373763 43319 373766
rect 199326 373764 199332 373766
rect 199396 373826 199402 373828
rect 199745 373826 199811 373829
rect 258073 373828 258139 373829
rect 199396 373824 199811 373826
rect 199396 373768 199750 373824
rect 199806 373768 199811 373824
rect 199396 373766 199811 373768
rect 199396 373764 199402 373766
rect 199745 373763 199811 373766
rect 258022 373764 258028 373828
rect 258092 373826 258139 373828
rect 262857 373826 262923 373829
rect 416037 373828 416103 373829
rect 421005 373828 421071 373829
rect 423029 373828 423095 373829
rect 426893 373828 426959 373829
rect 430573 373828 430639 373829
rect 268510 373826 268516 373828
rect 258092 373824 258184 373826
rect 258134 373768 258184 373824
rect 258092 373766 258184 373768
rect 262857 373824 268516 373826
rect 262857 373768 262862 373824
rect 262918 373768 268516 373824
rect 262857 373766 268516 373768
rect 258092 373764 258139 373766
rect 258073 373763 258139 373764
rect 262857 373763 262923 373766
rect 268510 373764 268516 373766
rect 268580 373764 268586 373828
rect 416037 373826 416084 373828
rect 415992 373824 416084 373826
rect 415992 373768 416042 373824
rect 415992 373766 416084 373768
rect 416037 373764 416084 373766
rect 416148 373764 416154 373828
rect 421005 373826 421052 373828
rect 420960 373824 421052 373826
rect 420960 373768 421010 373824
rect 420960 373766 421052 373768
rect 421005 373764 421052 373766
rect 421116 373764 421122 373828
rect 423029 373826 423076 373828
rect 422984 373824 423076 373826
rect 422984 373768 423034 373824
rect 422984 373766 423076 373768
rect 423029 373764 423076 373766
rect 423140 373764 423146 373828
rect 426893 373826 426940 373828
rect 426848 373824 426940 373826
rect 426848 373768 426898 373824
rect 426848 373766 426940 373768
rect 426893 373764 426940 373766
rect 427004 373764 427010 373828
rect 430573 373826 430620 373828
rect 430528 373824 430620 373826
rect 430528 373768 430578 373824
rect 430528 373766 430620 373768
rect 430573 373764 430620 373766
rect 430684 373764 430690 373828
rect 416037 373763 416103 373764
rect 421005 373763 421071 373764
rect 423029 373763 423095 373764
rect 426893 373763 426959 373764
rect 430573 373763 430639 373764
rect 95049 373692 95115 373693
rect 94998 373690 95004 373692
rect 94958 373630 95004 373690
rect 95068 373688 95115 373692
rect 96061 373692 96127 373693
rect 96061 373690 96108 373692
rect 95110 373632 95115 373688
rect 94998 373628 95004 373630
rect 95068 373628 95115 373632
rect 96016 373688 96108 373690
rect 96016 373632 96066 373688
rect 96016 373630 96108 373632
rect 95049 373627 95115 373628
rect 96061 373628 96108 373630
rect 96172 373628 96178 373692
rect 103278 373628 103284 373692
rect 103348 373690 103354 373692
rect 103513 373690 103579 373693
rect 107837 373692 107903 373693
rect 113541 373692 113607 373693
rect 118325 373692 118391 373693
rect 121361 373692 121427 373693
rect 107837 373690 107884 373692
rect 103348 373688 103579 373690
rect 103348 373632 103518 373688
rect 103574 373632 103579 373688
rect 103348 373630 103579 373632
rect 107792 373688 107884 373690
rect 107792 373632 107842 373688
rect 107792 373630 107884 373632
rect 103348 373628 103354 373630
rect 96061 373627 96127 373628
rect 103513 373627 103579 373630
rect 107837 373628 107884 373630
rect 107948 373628 107954 373692
rect 113541 373690 113588 373692
rect 113496 373688 113588 373690
rect 113496 373632 113546 373688
rect 113496 373630 113588 373632
rect 113541 373628 113588 373630
rect 113652 373628 113658 373692
rect 118325 373690 118372 373692
rect 118280 373688 118372 373690
rect 118280 373632 118330 373688
rect 118280 373630 118372 373632
rect 118325 373628 118372 373630
rect 118436 373628 118442 373692
rect 121310 373690 121316 373692
rect 121270 373630 121316 373690
rect 121380 373688 121427 373692
rect 205449 373690 205515 373693
rect 445845 373692 445911 373693
rect 455413 373692 455479 373693
rect 121422 373632 121427 373688
rect 121310 373628 121316 373630
rect 121380 373628 121427 373632
rect 107837 373627 107903 373628
rect 113541 373627 113607 373628
rect 118325 373627 118391 373628
rect 121361 373627 121427 373628
rect 122790 373688 205515 373690
rect 122790 373632 205454 373688
rect 205510 373632 205515 373688
rect 122790 373630 205515 373632
rect 110413 373556 110479 373557
rect 110413 373554 110460 373556
rect 110368 373552 110460 373554
rect 110368 373496 110418 373552
rect 110368 373494 110460 373496
rect 110413 373492 110460 373494
rect 110524 373492 110530 373556
rect 119838 373492 119844 373556
rect 119908 373554 119914 373556
rect 122790 373554 122850 373630
rect 205449 373627 205515 373630
rect 217542 373628 217548 373692
rect 217612 373690 217618 373692
rect 266302 373690 266308 373692
rect 217612 373630 266308 373690
rect 217612 373628 217618 373630
rect 266302 373628 266308 373630
rect 266372 373628 266378 373692
rect 445845 373690 445892 373692
rect 445800 373688 445892 373690
rect 445800 373632 445850 373688
rect 445800 373630 445892 373632
rect 445845 373628 445892 373630
rect 445956 373628 445962 373692
rect 455413 373690 455460 373692
rect 455368 373688 455460 373690
rect 455368 373632 455418 373688
rect 455368 373630 455460 373632
rect 455413 373628 455460 373630
rect 455524 373628 455530 373692
rect 445845 373627 445911 373628
rect 455413 373627 455479 373628
rect 124121 373556 124187 373557
rect 124070 373554 124076 373556
rect 119908 373494 122850 373554
rect 124030 373494 124076 373554
rect 124140 373552 124187 373556
rect 125685 373556 125751 373557
rect 128905 373556 128971 373557
rect 125685 373554 125732 373556
rect 124182 373496 124187 373552
rect 119908 373492 119914 373494
rect 124070 373492 124076 373494
rect 124140 373492 124187 373496
rect 125640 373552 125732 373554
rect 125640 373496 125690 373552
rect 125640 373494 125732 373496
rect 110413 373491 110479 373492
rect 124121 373491 124187 373492
rect 125685 373492 125732 373494
rect 125796 373492 125802 373556
rect 128854 373554 128860 373556
rect 128814 373494 128860 373554
rect 128924 373552 128971 373556
rect 128966 373496 128971 373552
rect 128854 373492 128860 373494
rect 128924 373492 128971 373496
rect 125685 373491 125751 373492
rect 128905 373491 128971 373492
rect 131021 373556 131087 373557
rect 133689 373556 133755 373557
rect 136449 373556 136515 373557
rect 151721 373556 151787 373557
rect 154113 373556 154179 373557
rect 131021 373552 131068 373556
rect 131132 373554 131138 373556
rect 133638 373554 133644 373556
rect 131021 373496 131026 373552
rect 131021 373492 131068 373496
rect 131132 373494 131178 373554
rect 133598 373494 133644 373554
rect 133708 373552 133755 373556
rect 136398 373554 136404 373556
rect 133750 373496 133755 373552
rect 131132 373492 131138 373494
rect 133638 373492 133644 373494
rect 133708 373492 133755 373496
rect 136358 373494 136404 373554
rect 136468 373552 136515 373556
rect 151670 373554 151676 373556
rect 136510 373496 136515 373552
rect 136398 373492 136404 373494
rect 136468 373492 136515 373496
rect 151630 373494 151676 373554
rect 151740 373552 151787 373556
rect 154062 373554 154068 373556
rect 151782 373496 151787 373552
rect 151670 373492 151676 373494
rect 151740 373492 151787 373496
rect 154022 373494 154068 373554
rect 154132 373552 154179 373556
rect 263685 373556 263751 373557
rect 447685 373556 447751 373557
rect 458173 373556 458239 373557
rect 263685 373554 263732 373556
rect 154174 373496 154179 373552
rect 154062 373492 154068 373494
rect 154132 373492 154179 373496
rect 263640 373552 263732 373554
rect 263640 373496 263690 373552
rect 263640 373494 263732 373496
rect 131021 373491 131087 373492
rect 133689 373491 133755 373492
rect 136449 373491 136515 373492
rect 151721 373491 151787 373492
rect 154113 373491 154179 373492
rect 263685 373492 263732 373494
rect 263796 373492 263802 373556
rect 447685 373554 447732 373556
rect 447640 373552 447732 373554
rect 447640 373496 447690 373552
rect 447640 373494 447732 373496
rect 447685 373492 447732 373494
rect 447796 373492 447802 373556
rect 458173 373554 458220 373556
rect 458128 373552 458220 373554
rect 458128 373496 458178 373552
rect 458128 373494 458220 373496
rect 458173 373492 458220 373494
rect 458284 373492 458290 373556
rect 263685 373491 263751 373492
rect 447685 373491 447751 373492
rect 458173 373491 458239 373492
rect 93669 373420 93735 373421
rect 98269 373420 98335 373421
rect 269205 373420 269271 373421
rect 452837 373420 452903 373421
rect 485773 373420 485839 373421
rect 93669 373418 93716 373420
rect 93624 373416 93716 373418
rect 93624 373360 93674 373416
rect 93624 373358 93716 373360
rect 93669 373356 93716 373358
rect 93780 373356 93786 373420
rect 98269 373418 98316 373420
rect 98224 373416 98316 373418
rect 98224 373360 98274 373416
rect 98224 373358 98316 373360
rect 98269 373356 98316 373358
rect 98380 373356 98386 373420
rect 269205 373418 269252 373420
rect 269160 373416 269252 373418
rect 269160 373360 269210 373416
rect 269160 373358 269252 373360
rect 269205 373356 269252 373358
rect 269316 373356 269322 373420
rect 452837 373418 452884 373420
rect 452792 373416 452884 373418
rect 452792 373360 452842 373416
rect 452792 373358 452884 373360
rect 452837 373356 452884 373358
rect 452948 373356 452954 373420
rect 485773 373418 485820 373420
rect 485728 373416 485820 373418
rect 485728 373360 485778 373416
rect 485728 373358 485820 373360
rect 485773 373356 485820 373358
rect 485884 373356 485890 373420
rect 93669 373355 93735 373356
rect 98269 373355 98335 373356
rect 269205 373355 269271 373356
rect 452837 373355 452903 373356
rect 485773 373355 485839 373356
rect 88333 373284 88399 373285
rect 95969 373284 96035 373285
rect 88333 373282 88380 373284
rect 88288 373280 88380 373282
rect 88288 373224 88338 373280
rect 88288 373222 88380 373224
rect 88333 373220 88380 373222
rect 88444 373220 88450 373284
rect 95918 373282 95924 373284
rect 95878 373222 95924 373282
rect 95988 373280 96035 373284
rect 100845 373284 100911 373285
rect 242893 373284 242959 373285
rect 261293 373284 261359 373285
rect 100845 373282 100892 373284
rect 96030 373224 96035 373280
rect 95918 373220 95924 373222
rect 95988 373220 96035 373224
rect 100800 373280 100892 373282
rect 100800 373224 100850 373280
rect 100800 373222 100892 373224
rect 88333 373219 88399 373220
rect 95969 373219 96035 373220
rect 100845 373220 100892 373222
rect 100956 373220 100962 373284
rect 242893 373282 242940 373284
rect 242848 373280 242940 373282
rect 242848 373224 242898 373280
rect 242848 373222 242940 373224
rect 242893 373220 242940 373222
rect 243004 373220 243010 373284
rect 261293 373282 261340 373284
rect 261248 373280 261340 373282
rect 261248 373224 261298 373280
rect 261248 373222 261340 373224
rect 261293 373220 261340 373222
rect 261404 373220 261410 373284
rect 279182 373220 279188 373284
rect 279252 373282 279258 373284
rect 358813 373282 358879 373285
rect 279252 373280 358879 373282
rect 279252 373224 358818 373280
rect 358874 373224 358879 373280
rect 279252 373222 358879 373224
rect 279252 373220 279258 373222
rect 100845 373219 100911 373220
rect 242893 373219 242959 373220
rect 261293 373219 261359 373220
rect 358813 373219 358879 373222
rect 90173 373148 90239 373149
rect 92381 373148 92447 373149
rect 235993 373148 236059 373149
rect 90173 373146 90220 373148
rect 90128 373144 90220 373146
rect 90128 373088 90178 373144
rect 90128 373086 90220 373088
rect 90173 373084 90220 373086
rect 90284 373084 90290 373148
rect 92381 373144 92428 373148
rect 92492 373146 92498 373148
rect 92381 373088 92386 373144
rect 92381 373084 92428 373088
rect 92492 373086 92538 373146
rect 92492 373084 92498 373086
rect 235942 373084 235948 373148
rect 236012 373146 236059 373148
rect 253933 373148 253999 373149
rect 255405 373148 255471 373149
rect 271965 373148 272031 373149
rect 300853 373148 300919 373149
rect 253933 373146 253980 373148
rect 236012 373144 236104 373146
rect 236054 373088 236104 373144
rect 236012 373086 236104 373088
rect 253888 373144 253980 373146
rect 253888 373088 253938 373144
rect 253888 373086 253980 373088
rect 236012 373084 236059 373086
rect 90173 373083 90239 373084
rect 92381 373083 92447 373084
rect 235993 373083 236059 373084
rect 253933 373084 253980 373086
rect 254044 373084 254050 373148
rect 255405 373146 255452 373148
rect 255360 373144 255452 373146
rect 255360 373088 255410 373144
rect 255360 373086 255452 373088
rect 255405 373084 255452 373086
rect 255516 373084 255522 373148
rect 271965 373146 272012 373148
rect 271920 373144 272012 373146
rect 271920 373088 271970 373144
rect 271920 373086 272012 373088
rect 271965 373084 272012 373086
rect 272076 373084 272082 373148
rect 300853 373146 300900 373148
rect 300808 373144 300900 373146
rect 300808 373088 300858 373144
rect 300808 373086 300900 373088
rect 300853 373084 300900 373086
rect 300964 373084 300970 373148
rect 253933 373083 253999 373084
rect 255405 373083 255471 373084
rect 271965 373083 272031 373084
rect 300853 373083 300919 373084
rect 55581 373010 55647 373013
rect 59445 373010 59511 373013
rect 55581 373008 59511 373010
rect 55581 372952 55586 373008
rect 55642 372952 59450 373008
rect 59506 372952 59511 373008
rect 55581 372950 59511 372952
rect 55581 372947 55647 372950
rect 59445 372947 59511 372950
rect 56501 372874 56567 372877
rect 57094 372874 57100 372876
rect 56501 372872 57100 372874
rect 56501 372816 56506 372872
rect 56562 372816 57100 372872
rect 56501 372814 57100 372816
rect 56501 372811 56567 372814
rect 57094 372812 57100 372814
rect 57164 372812 57170 372876
rect 55673 372738 55739 372741
rect 57278 372738 57284 372740
rect 55673 372736 57284 372738
rect 55673 372680 55678 372736
rect 55734 372680 57284 372736
rect 55673 372678 57284 372680
rect 55673 372675 55739 372678
rect 57278 372676 57284 372678
rect 57348 372676 57354 372740
rect 58617 372738 58683 372741
rect 62113 372738 62179 372741
rect 58617 372736 62179 372738
rect 58617 372680 58622 372736
rect 58678 372680 62118 372736
rect 62174 372680 62179 372736
rect 58617 372678 62179 372680
rect 58617 372675 58683 372678
rect 62113 372675 62179 372678
rect 199142 372676 199148 372740
rect 199212 372738 199218 372740
rect 199469 372738 199535 372741
rect 199212 372736 199535 372738
rect 199212 372680 199474 372736
rect 199530 372680 199535 372736
rect 199212 372678 199535 372680
rect 199212 372676 199218 372678
rect 199469 372675 199535 372678
rect 209998 372676 210004 372740
rect 210068 372738 210074 372740
rect 210969 372738 211035 372741
rect 217041 372740 217107 372741
rect 216990 372738 216996 372740
rect 210068 372736 211035 372738
rect 210068 372680 210974 372736
rect 211030 372680 211035 372736
rect 210068 372678 211035 372680
rect 216950 372678 216996 372738
rect 217060 372736 217107 372740
rect 217102 372680 217107 372736
rect 210068 372676 210074 372678
rect 210969 372675 211035 372678
rect 216990 372676 216996 372678
rect 217060 372676 217107 372680
rect 217041 372675 217107 372676
rect 371601 372738 371667 372741
rect 376886 372738 376892 372740
rect 371601 372736 376892 372738
rect 371601 372680 371606 372736
rect 371662 372680 376892 372736
rect 371601 372678 376892 372680
rect 371601 372675 371667 372678
rect 77201 372604 77267 372605
rect 77150 372602 77156 372604
rect 77110 372542 77156 372602
rect 77220 372600 77267 372604
rect 77262 372544 77267 372600
rect 77150 372540 77156 372542
rect 77220 372540 77267 372544
rect 84510 372540 84516 372604
rect 84580 372602 84586 372604
rect 85481 372602 85547 372605
rect 86585 372604 86651 372605
rect 88057 372604 88123 372605
rect 89345 372604 89411 372605
rect 90081 372604 90147 372605
rect 86534 372602 86540 372604
rect 84580 372600 85547 372602
rect 84580 372544 85486 372600
rect 85542 372544 85547 372600
rect 84580 372542 85547 372544
rect 86494 372542 86540 372602
rect 86604 372600 86651 372604
rect 88006 372602 88012 372604
rect 86646 372544 86651 372600
rect 84580 372540 84586 372542
rect 77201 372539 77267 372540
rect 85481 372539 85547 372542
rect 86534 372540 86540 372542
rect 86604 372540 86651 372544
rect 87966 372542 88012 372602
rect 88076 372600 88123 372604
rect 89294 372602 89300 372604
rect 88118 372544 88123 372600
rect 88006 372540 88012 372542
rect 88076 372540 88123 372544
rect 89254 372542 89300 372602
rect 89364 372600 89411 372604
rect 90030 372602 90036 372604
rect 89406 372544 89411 372600
rect 89294 372540 89300 372542
rect 89364 372540 89411 372544
rect 89990 372542 90036 372602
rect 90100 372600 90147 372604
rect 90142 372544 90147 372600
rect 90030 372540 90036 372542
rect 90100 372540 90147 372544
rect 91502 372540 91508 372604
rect 91572 372602 91578 372604
rect 92197 372602 92263 372605
rect 91572 372600 92263 372602
rect 91572 372544 92202 372600
rect 92258 372544 92263 372600
rect 91572 372542 92263 372544
rect 91572 372540 91578 372542
rect 86585 372539 86651 372540
rect 88057 372539 88123 372540
rect 89345 372539 89411 372540
rect 90081 372539 90147 372540
rect 92197 372539 92263 372542
rect 93342 372540 93348 372604
rect 93412 372602 93418 372604
rect 93577 372602 93643 372605
rect 108849 372604 108915 372605
rect 108798 372602 108804 372604
rect 93412 372600 93643 372602
rect 93412 372544 93582 372600
rect 93638 372544 93643 372600
rect 93412 372542 93643 372544
rect 108758 372542 108804 372602
rect 108868 372600 108915 372604
rect 108910 372544 108915 372600
rect 93412 372540 93418 372542
rect 93577 372539 93643 372542
rect 108798 372540 108804 372542
rect 108868 372540 108915 372544
rect 113214 372540 113220 372604
rect 113284 372602 113290 372604
rect 114001 372602 114067 372605
rect 183185 372604 183251 372605
rect 183134 372602 183140 372604
rect 113284 372600 114067 372602
rect 113284 372544 114006 372600
rect 114062 372544 114067 372600
rect 113284 372542 114067 372544
rect 183094 372542 183140 372602
rect 183204 372600 183251 372604
rect 183246 372544 183251 372600
rect 113284 372540 113290 372542
rect 108849 372539 108915 372540
rect 114001 372539 114067 372542
rect 183134 372540 183140 372542
rect 183204 372540 183251 372544
rect 183185 372539 183251 372540
rect 236085 372602 236151 372605
rect 238109 372604 238175 372605
rect 239305 372604 239371 372605
rect 240409 372604 240475 372605
rect 241513 372604 241579 372605
rect 236494 372602 236500 372604
rect 236085 372600 236500 372602
rect 236085 372544 236090 372600
rect 236146 372544 236500 372600
rect 236085 372542 236500 372544
rect 236085 372539 236151 372542
rect 236494 372540 236500 372542
rect 236564 372540 236570 372604
rect 238109 372600 238156 372604
rect 238220 372602 238226 372604
rect 239254 372602 239260 372604
rect 238109 372544 238114 372600
rect 238109 372540 238156 372544
rect 238220 372542 238266 372602
rect 239214 372542 239260 372602
rect 239324 372600 239371 372604
rect 240358 372602 240364 372604
rect 239366 372544 239371 372600
rect 238220 372540 238226 372542
rect 239254 372540 239260 372542
rect 239324 372540 239371 372544
rect 240318 372542 240364 372602
rect 240428 372600 240475 372604
rect 241462 372602 241468 372604
rect 240470 372544 240475 372600
rect 240358 372540 240364 372542
rect 240428 372540 240475 372544
rect 241422 372542 241468 372602
rect 241532 372600 241579 372604
rect 241574 372544 241579 372600
rect 241462 372540 241468 372542
rect 241532 372540 241579 372544
rect 238109 372539 238175 372540
rect 239305 372539 239371 372540
rect 240409 372539 240475 372540
rect 241513 372539 241579 372540
rect 245653 372602 245719 372605
rect 248413 372604 248479 372605
rect 251173 372604 251239 372605
rect 256693 372604 256759 372605
rect 259453 372604 259519 372605
rect 245878 372602 245884 372604
rect 245653 372600 245884 372602
rect 245653 372544 245658 372600
rect 245714 372544 245884 372600
rect 245653 372542 245884 372544
rect 245653 372539 245719 372542
rect 245878 372540 245884 372542
rect 245948 372540 245954 372604
rect 248413 372600 248460 372604
rect 248524 372602 248530 372604
rect 251173 372602 251220 372604
rect 248413 372544 248418 372600
rect 248413 372540 248460 372544
rect 248524 372542 248570 372602
rect 251128 372600 251220 372602
rect 251128 372544 251178 372600
rect 251128 372542 251220 372544
rect 248524 372540 248530 372542
rect 251173 372540 251220 372542
rect 251284 372540 251290 372604
rect 256693 372602 256740 372604
rect 256648 372600 256740 372602
rect 256648 372544 256698 372600
rect 256648 372542 256740 372544
rect 256693 372540 256740 372542
rect 256804 372540 256810 372604
rect 259453 372602 259500 372604
rect 259408 372600 259500 372602
rect 259408 372544 259458 372600
rect 259408 372542 259500 372544
rect 259453 372540 259500 372542
rect 259564 372540 259570 372604
rect 259637 372602 259703 372605
rect 273253 372604 273319 372605
rect 260046 372602 260052 372604
rect 259637 372600 260052 372602
rect 259637 372544 259642 372600
rect 259698 372544 260052 372600
rect 259637 372542 260052 372544
rect 248413 372539 248479 372540
rect 251173 372539 251239 372540
rect 256693 372539 256759 372540
rect 259453 372539 259519 372540
rect 259637 372539 259703 372542
rect 260046 372540 260052 372542
rect 260116 372540 260122 372604
rect 273253 372602 273300 372604
rect 273208 372600 273300 372602
rect 273208 372544 273258 372600
rect 273208 372542 273300 372544
rect 273253 372540 273300 372542
rect 273364 372540 273370 372604
rect 310513 372602 310579 372605
rect 310646 372602 310652 372604
rect 310513 372600 310652 372602
rect 310513 372544 310518 372600
rect 310574 372544 310652 372600
rect 310513 372542 310652 372544
rect 273253 372539 273319 372540
rect 310513 372539 310579 372542
rect 310646 372540 310652 372542
rect 310716 372540 310722 372604
rect 313273 372602 313339 372605
rect 313406 372602 313412 372604
rect 313273 372600 313412 372602
rect 313273 372544 313278 372600
rect 313334 372544 313412 372600
rect 313273 372542 313412 372544
rect 313273 372539 313339 372542
rect 313406 372540 313412 372542
rect 313476 372540 313482 372604
rect 78489 372468 78555 372469
rect 79961 372468 80027 372469
rect 78438 372466 78444 372468
rect 78398 372406 78444 372466
rect 78508 372464 78555 372468
rect 79910 372466 79916 372468
rect 78550 372408 78555 372464
rect 78438 372404 78444 372406
rect 78508 372404 78555 372408
rect 79870 372406 79916 372466
rect 79980 372464 80027 372468
rect 80022 372408 80027 372464
rect 79910 372404 79916 372406
rect 79980 372404 80027 372408
rect 84694 372404 84700 372468
rect 84764 372466 84770 372468
rect 85113 372466 85179 372469
rect 102777 372468 102843 372469
rect 102726 372466 102732 372468
rect 84764 372464 85179 372466
rect 84764 372408 85118 372464
rect 85174 372408 85179 372464
rect 84764 372406 85179 372408
rect 102686 372406 102732 372466
rect 102796 372464 102843 372468
rect 102838 372408 102843 372464
rect 84764 372404 84770 372406
rect 78489 372403 78555 372404
rect 79961 372403 80027 372404
rect 85113 372403 85179 372406
rect 102726 372404 102732 372406
rect 102796 372404 102843 372408
rect 117078 372404 117084 372468
rect 117148 372466 117154 372468
rect 218605 372466 218671 372469
rect 276289 372466 276355 372469
rect 277158 372466 277164 372468
rect 117148 372464 277164 372466
rect 117148 372408 218610 372464
rect 218666 372408 276294 372464
rect 276350 372408 277164 372464
rect 117148 372406 277164 372408
rect 117148 372404 117154 372406
rect 102777 372403 102843 372404
rect 218605 372403 218671 372406
rect 276289 372403 276355 372406
rect 277158 372404 277164 372406
rect 277228 372404 277234 372468
rect 304993 372466 305059 372469
rect 305310 372466 305316 372468
rect 304993 372464 305316 372466
rect 304993 372408 304998 372464
rect 305054 372408 305316 372464
rect 304993 372406 305316 372408
rect 304993 372403 305059 372406
rect 305310 372404 305316 372406
rect 305380 372404 305386 372468
rect 376710 372466 376770 372678
rect 376886 372676 376892 372678
rect 376956 372676 376962 372740
rect 408493 372604 408559 372605
rect 426433 372604 426499 372605
rect 408493 372602 408540 372604
rect 408448 372600 408540 372602
rect 408448 372544 408498 372600
rect 408448 372542 408540 372544
rect 408493 372540 408540 372542
rect 408604 372540 408610 372604
rect 426382 372540 426388 372604
rect 426452 372602 426499 372604
rect 433333 372602 433399 372605
rect 433558 372602 433564 372604
rect 426452 372600 426544 372602
rect 426494 372544 426544 372600
rect 426452 372542 426544 372544
rect 433333 372600 433564 372602
rect 433333 372544 433338 372600
rect 433394 372544 433564 372600
rect 433333 372542 433564 372544
rect 426452 372540 426499 372542
rect 408493 372539 408559 372540
rect 426433 372539 426499 372540
rect 433333 372539 433399 372542
rect 433558 372540 433564 372542
rect 433628 372540 433634 372604
rect 437473 372602 437539 372605
rect 438342 372602 438348 372604
rect 437473 372600 438348 372602
rect 437473 372544 437478 372600
rect 437534 372544 438348 372600
rect 437473 372542 438348 372544
rect 437473 372539 437539 372542
rect 438342 372540 438348 372542
rect 438412 372540 438418 372604
rect 431166 372466 431172 372468
rect 376710 372406 431172 372466
rect 431166 372404 431172 372406
rect 431236 372404 431242 372468
rect 80513 372332 80579 372333
rect 80462 372330 80468 372332
rect 80422 372270 80468 372330
rect 80532 372328 80579 372332
rect 80574 372272 80579 372328
rect 80462 372268 80468 372270
rect 80532 372268 80579 372272
rect 80513 372267 80579 372268
rect 81893 372332 81959 372333
rect 102041 372332 102107 372333
rect 81893 372328 81940 372332
rect 82004 372330 82010 372332
rect 101990 372330 101996 372332
rect 81893 372272 81898 372328
rect 81893 372268 81940 372272
rect 82004 372270 82050 372330
rect 101950 372270 101996 372330
rect 102060 372328 102107 372332
rect 102102 372272 102107 372328
rect 82004 372268 82010 372270
rect 101990 372268 101996 372270
rect 102060 372268 102107 372272
rect 109534 372268 109540 372332
rect 109604 372330 109610 372332
rect 117957 372330 118023 372333
rect 109604 372328 118023 372330
rect 109604 372272 117962 372328
rect 118018 372272 118023 372328
rect 109604 372270 118023 372272
rect 109604 372268 109610 372270
rect 81893 372267 81959 372268
rect 102041 372267 102107 372268
rect 117957 372267 118023 372270
rect 118182 372268 118188 372332
rect 118252 372330 118258 372332
rect 215753 372330 215819 372333
rect 277526 372330 277532 372332
rect 118252 372328 277532 372330
rect 118252 372272 215758 372328
rect 215814 372272 277532 372328
rect 118252 372270 277532 372272
rect 118252 372268 118258 372270
rect 215753 372267 215819 372270
rect 277526 372268 277532 372270
rect 277596 372330 277602 372332
rect 278681 372330 278747 372333
rect 277596 372328 278747 372330
rect 277596 372272 278686 372328
rect 278742 372272 278747 372328
rect 277596 372270 278747 372272
rect 277596 372268 277602 372270
rect 278681 372267 278747 372270
rect 470593 372330 470659 372333
rect 470726 372330 470732 372332
rect 470593 372328 470732 372330
rect 470593 372272 470598 372328
rect 470654 372272 470732 372328
rect 470593 372270 470732 372272
rect 470593 372267 470659 372270
rect 470726 372268 470732 372270
rect 470796 372268 470802 372332
rect 76598 372132 76604 372196
rect 76668 372194 76674 372196
rect 77017 372194 77083 372197
rect 76668 372192 77083 372194
rect 76668 372136 77022 372192
rect 77078 372136 77083 372192
rect 76668 372134 77083 372136
rect 76668 372132 76674 372134
rect 77017 372131 77083 372134
rect 111742 372132 111748 372196
rect 111812 372194 111818 372196
rect 211613 372194 211679 372197
rect 222101 372194 222167 372197
rect 270217 372194 270283 372197
rect 111812 372192 270283 372194
rect 111812 372136 211618 372192
rect 211674 372136 222106 372192
rect 222162 372136 270222 372192
rect 270278 372136 270283 372192
rect 111812 372134 270283 372136
rect 111812 372132 111818 372134
rect 211613 372131 211679 372134
rect 222101 372131 222167 372134
rect 270217 372131 270283 372134
rect 404353 372194 404419 372197
rect 503161 372196 503227 372197
rect 503529 372196 503595 372197
rect 404854 372194 404860 372196
rect 404353 372192 404860 372194
rect 404353 372136 404358 372192
rect 404414 372136 404860 372192
rect 404353 372134 404860 372136
rect 404353 372131 404419 372134
rect 404854 372132 404860 372134
rect 404924 372132 404930 372196
rect 503110 372194 503116 372196
rect 503070 372134 503116 372194
rect 503180 372192 503227 372196
rect 503478 372194 503484 372196
rect 503222 372136 503227 372192
rect 503110 372132 503116 372134
rect 503180 372132 503227 372136
rect 503438 372134 503484 372194
rect 503548 372192 503595 372196
rect 503590 372136 503595 372192
rect 503478 372132 503484 372134
rect 503548 372132 503595 372136
rect 503161 372131 503227 372132
rect 503529 372131 503595 372132
rect 117957 372058 118023 372061
rect 222009 372058 222075 372061
rect 270309 372058 270375 372061
rect 117957 372056 210250 372058
rect 117957 372000 117962 372056
rect 118018 372000 210250 372056
rect 117957 371998 210250 372000
rect 117957 371995 118023 371998
rect 83825 371924 83891 371925
rect 104617 371924 104683 371925
rect 83774 371922 83780 371924
rect 83734 371862 83780 371922
rect 83844 371920 83891 371924
rect 104566 371922 104572 371924
rect 83886 371864 83891 371920
rect 83774 371860 83780 371862
rect 83844 371860 83891 371864
rect 104526 371862 104572 371922
rect 104636 371920 104683 371924
rect 104678 371864 104683 371920
rect 104566 371860 104572 371862
rect 104636 371860 104683 371864
rect 112846 371860 112852 371924
rect 112916 371922 112922 371924
rect 210049 371922 210115 371925
rect 112916 371920 210115 371922
rect 112916 371864 210054 371920
rect 210110 371864 210115 371920
rect 112916 371862 210115 371864
rect 210190 371922 210250 371998
rect 213870 372056 270375 372058
rect 213870 372000 222014 372056
rect 222070 372000 270314 372056
rect 270370 372000 270375 372056
rect 213870 371998 270375 372000
rect 210325 371922 210391 371925
rect 210190 371920 210391 371922
rect 210190 371864 210330 371920
rect 210386 371864 210391 371920
rect 210190 371862 210391 371864
rect 112916 371860 112922 371862
rect 83825 371859 83891 371860
rect 104617 371859 104683 371860
rect 210049 371859 210115 371862
rect 210325 371859 210391 371862
rect 105302 371724 105308 371788
rect 105372 371786 105378 371788
rect 105905 371786 105971 371789
rect 105372 371784 105971 371786
rect 105372 371728 105910 371784
rect 105966 371728 105971 371784
rect 105372 371726 105971 371728
rect 105372 371724 105378 371726
rect 105905 371723 105971 371726
rect 114502 371724 114508 371788
rect 114572 371786 114578 371788
rect 212257 371786 212323 371789
rect 213870 371786 213930 371998
rect 222009 371995 222075 371998
rect 270309 371995 270375 371998
rect 396073 372058 396139 372061
rect 397453 372060 397519 372061
rect 396206 372058 396212 372060
rect 396073 372056 396212 372058
rect 396073 372000 396078 372056
rect 396134 372000 396212 372056
rect 396073 371998 396212 372000
rect 396073 371995 396139 371998
rect 396206 371996 396212 371998
rect 396276 371996 396282 372060
rect 397453 372058 397500 372060
rect 397408 372056 397500 372058
rect 397408 372000 397458 372056
rect 397408 371998 397500 372000
rect 397453 371996 397500 371998
rect 397564 371996 397570 372060
rect 398833 372058 398899 372061
rect 400213 372060 400279 372061
rect 398966 372058 398972 372060
rect 398833 372056 398972 372058
rect 398833 372000 398838 372056
rect 398894 372000 398972 372056
rect 398833 371998 398972 372000
rect 397453 371995 397519 371996
rect 398833 371995 398899 371998
rect 398966 371996 398972 371998
rect 399036 371996 399042 372060
rect 400213 372058 400260 372060
rect 400168 372056 400260 372058
rect 400168 372000 400218 372056
rect 400168 371998 400260 372000
rect 400213 371996 400260 371998
rect 400324 371996 400330 372060
rect 409873 372058 409939 372061
rect 410006 372058 410012 372060
rect 409873 372056 410012 372058
rect 409873 372000 409878 372056
rect 409934 372000 410012 372056
rect 409873 371998 410012 372000
rect 400213 371995 400279 371996
rect 409873 371995 409939 371998
rect 410006 371996 410012 371998
rect 410076 371996 410082 372060
rect 271965 371922 272031 371925
rect 114572 371784 213930 371786
rect 114572 371728 212262 371784
rect 212318 371728 213930 371784
rect 114572 371726 213930 371728
rect 219390 371920 272031 371922
rect 219390 371864 271970 371920
rect 272026 371864 272031 371920
rect 219390 371862 272031 371864
rect 114572 371724 114578 371726
rect 212257 371723 212323 371726
rect 97574 371588 97580 371652
rect 97644 371650 97650 371652
rect 97717 371650 97783 371653
rect 97644 371648 97783 371650
rect 97644 371592 97722 371648
rect 97778 371592 97783 371648
rect 97644 371590 97783 371592
rect 97644 371588 97650 371590
rect 97717 371587 97783 371590
rect 98126 371588 98132 371652
rect 98196 371650 98202 371652
rect 99281 371650 99347 371653
rect 98196 371648 99347 371650
rect 98196 371592 99286 371648
rect 99342 371592 99347 371648
rect 98196 371590 99347 371592
rect 98196 371588 98202 371590
rect 99281 371587 99347 371590
rect 99966 371588 99972 371652
rect 100036 371650 100042 371652
rect 100109 371650 100175 371653
rect 100036 371648 100175 371650
rect 100036 371592 100114 371648
rect 100170 371592 100175 371648
rect 100036 371590 100175 371592
rect 100036 371588 100042 371590
rect 100109 371587 100175 371590
rect 210049 371650 210115 371653
rect 213637 371650 213703 371653
rect 218329 371650 218395 371653
rect 219390 371650 219450 371862
rect 271965 371859 272031 371862
rect 377438 371860 377444 371924
rect 377508 371922 377514 371924
rect 381077 371922 381143 371925
rect 433374 371922 433380 371924
rect 377508 371920 433380 371922
rect 377508 371864 381082 371920
rect 381138 371864 433380 371920
rect 377508 371862 433380 371864
rect 377508 371860 377514 371862
rect 381077 371859 381143 371862
rect 433374 371860 433380 371862
rect 433444 371860 433450 371924
rect 220721 371786 220787 371789
rect 275369 371788 275435 371789
rect 275318 371786 275324 371788
rect 220721 371784 275324 371786
rect 275388 371786 275435 371788
rect 317413 371786 317479 371789
rect 317822 371786 317828 371788
rect 275388 371784 275516 371786
rect 220721 371728 220726 371784
rect 220782 371728 275324 371784
rect 275430 371728 275516 371784
rect 220721 371726 275324 371728
rect 220721 371723 220787 371726
rect 275318 371724 275324 371726
rect 275388 371726 275516 371728
rect 317413 371784 317828 371786
rect 317413 371728 317418 371784
rect 317474 371728 317828 371784
rect 317413 371726 317828 371728
rect 275388 371724 275435 371726
rect 275369 371723 275435 371724
rect 317413 371723 317479 371726
rect 317822 371724 317828 371726
rect 317892 371724 317898 371788
rect 373809 371786 373875 371789
rect 439446 371786 439452 371788
rect 373809 371784 439452 371786
rect 373809 371728 373814 371784
rect 373870 371728 439452 371784
rect 373809 371726 439452 371728
rect 373809 371723 373875 371726
rect 439446 371724 439452 371726
rect 439516 371786 439522 371788
rect 439865 371786 439931 371789
rect 439516 371784 439931 371786
rect 439516 371728 439870 371784
rect 439926 371728 439931 371784
rect 439516 371726 439931 371728
rect 439516 371724 439522 371726
rect 439865 371723 439931 371726
rect 210049 371648 219450 371650
rect 210049 371592 210054 371648
rect 210110 371592 213642 371648
rect 213698 371592 218334 371648
rect 218390 371592 219450 371648
rect 210049 371590 219450 371592
rect 247033 371650 247099 371653
rect 247902 371650 247908 371652
rect 247033 371648 247908 371650
rect 247033 371592 247038 371648
rect 247094 371592 247908 371648
rect 247033 371590 247908 371592
rect 210049 371587 210115 371590
rect 213637 371587 213703 371590
rect 218329 371587 218395 371590
rect 247033 371587 247099 371590
rect 247902 371588 247908 371590
rect 247972 371588 247978 371652
rect 249885 371650 249951 371653
rect 250294 371650 250300 371652
rect 249885 371648 250300 371650
rect 249885 371592 249890 371648
rect 249946 371592 250300 371648
rect 249885 371590 250300 371592
rect 249885 371587 249951 371590
rect 250294 371588 250300 371590
rect 250364 371588 250370 371652
rect 251173 371650 251239 371653
rect 251950 371650 251956 371652
rect 251173 371648 251956 371650
rect 251173 371592 251178 371648
rect 251234 371592 251956 371648
rect 251173 371590 251956 371592
rect 251173 371587 251239 371590
rect 251950 371588 251956 371590
rect 252020 371588 252026 371652
rect 325877 371650 325943 371653
rect 326654 371650 326660 371652
rect 325877 371648 326660 371650
rect 325877 371592 325882 371648
rect 325938 371592 326660 371648
rect 325877 371590 326660 371592
rect 325877 371587 325943 371590
rect 326654 371588 326660 371590
rect 326724 371588 326730 371652
rect 401593 371650 401659 371653
rect 411253 371652 411319 371653
rect 402278 371650 402284 371652
rect 401593 371648 402284 371650
rect 401593 371592 401598 371648
rect 401654 371592 402284 371648
rect 401593 371590 402284 371592
rect 401593 371587 401659 371590
rect 402278 371588 402284 371590
rect 402348 371588 402354 371652
rect 411253 371650 411300 371652
rect 411208 371648 411300 371650
rect 411208 371592 411258 371648
rect 411208 371590 411300 371592
rect 411253 371588 411300 371590
rect 411364 371588 411370 371652
rect 418337 371650 418403 371653
rect 418838 371650 418844 371652
rect 418337 371648 418844 371650
rect 418337 371592 418342 371648
rect 418398 371592 418844 371648
rect 418337 371590 418844 371592
rect 411253 371587 411319 371588
rect 418337 371587 418403 371590
rect 418838 371588 418844 371590
rect 418908 371588 418914 371652
rect 423673 371650 423739 371653
rect 427813 371652 427879 371653
rect 423990 371650 423996 371652
rect 423673 371648 423996 371650
rect 423673 371592 423678 371648
rect 423734 371592 423996 371648
rect 423673 371590 423996 371592
rect 423673 371587 423739 371590
rect 423990 371588 423996 371590
rect 424060 371588 424066 371652
rect 427813 371650 427860 371652
rect 427768 371648 427860 371650
rect 427768 371592 427818 371648
rect 427768 371590 427860 371592
rect 427813 371588 427860 371590
rect 427924 371588 427930 371652
rect 462313 371650 462379 371653
rect 462630 371650 462636 371652
rect 462313 371648 462636 371650
rect 462313 371592 462318 371648
rect 462374 371592 462636 371648
rect 462313 371590 462636 371592
rect 427813 371587 427879 371588
rect 462313 371587 462379 371590
rect 462630 371588 462636 371590
rect 462700 371588 462706 371652
rect 465073 371650 465139 371653
rect 465390 371650 465396 371652
rect 465073 371648 465396 371650
rect 465073 371592 465078 371648
rect 465134 371592 465396 371648
rect 465073 371590 465396 371592
rect 465073 371587 465139 371590
rect 465390 371588 465396 371590
rect 465460 371588 465466 371652
rect 477493 371650 477559 371653
rect 478086 371650 478092 371652
rect 477493 371648 478092 371650
rect 477493 371592 477498 371648
rect 477554 371592 478092 371648
rect 477493 371590 478092 371592
rect 477493 371587 477559 371590
rect 478086 371588 478092 371590
rect 478156 371588 478162 371652
rect -960 371228 480 371468
rect 100702 371452 100708 371516
rect 100772 371514 100778 371516
rect 101029 371514 101095 371517
rect 100772 371512 101095 371514
rect 100772 371456 101034 371512
rect 101090 371456 101095 371512
rect 100772 371454 101095 371456
rect 100772 371452 100778 371454
rect 101029 371451 101095 371454
rect 182817 371514 182883 371517
rect 183318 371514 183324 371516
rect 182817 371512 183324 371514
rect 182817 371456 182822 371512
rect 182878 371456 183324 371512
rect 182817 371454 183324 371456
rect 182817 371451 182883 371454
rect 183318 371452 183324 371454
rect 183388 371452 183394 371516
rect 210325 371514 210391 371517
rect 218145 371514 218211 371517
rect 262765 371514 262831 371517
rect 210325 371512 262831 371514
rect 210325 371456 210330 371512
rect 210386 371456 218150 371512
rect 218206 371456 262770 371512
rect 262826 371456 262831 371512
rect 210325 371454 262831 371456
rect 210325 371451 210391 371454
rect 218145 371451 218211 371454
rect 262765 371451 262831 371454
rect 264973 371514 265039 371517
rect 265750 371514 265756 371516
rect 264973 371512 265756 371514
rect 264973 371456 264978 371512
rect 265034 371456 265756 371512
rect 264973 371454 265756 371456
rect 264973 371451 265039 371454
rect 265750 371452 265756 371454
rect 265820 371452 265826 371516
rect 273345 371514 273411 371517
rect 273662 371514 273668 371516
rect 273345 371512 273668 371514
rect 273345 371456 273350 371512
rect 273406 371456 273668 371512
rect 273345 371454 273668 371456
rect 273345 371451 273411 371454
rect 273662 371452 273668 371454
rect 273732 371452 273738 371516
rect 407113 371514 407179 371517
rect 407246 371514 407252 371516
rect 407113 371512 407252 371514
rect 407113 371456 407118 371512
rect 407174 371456 407252 371512
rect 407113 371454 407252 371456
rect 407113 371451 407179 371454
rect 407246 371452 407252 371454
rect 407316 371452 407322 371516
rect 411253 371514 411319 371517
rect 411846 371514 411852 371516
rect 411253 371512 411852 371514
rect 411253 371456 411258 371512
rect 411314 371456 411852 371512
rect 411253 371454 411852 371456
rect 411253 371451 411319 371454
rect 411846 371452 411852 371454
rect 411916 371452 411922 371516
rect 418102 371452 418108 371516
rect 418172 371514 418178 371516
rect 418245 371514 418311 371517
rect 418172 371512 418311 371514
rect 418172 371456 418250 371512
rect 418306 371456 418311 371512
rect 418172 371454 418311 371456
rect 418172 371452 418178 371454
rect 418245 371451 418311 371454
rect 420913 371514 420979 371517
rect 480253 371516 480319 371517
rect 421230 371514 421236 371516
rect 420913 371512 421236 371514
rect 420913 371456 420918 371512
rect 420974 371456 421236 371512
rect 420913 371454 421236 371456
rect 420913 371451 420979 371454
rect 421230 371452 421236 371454
rect 421300 371452 421306 371516
rect 480253 371512 480300 371516
rect 480364 371514 480370 371516
rect 480253 371456 480258 371512
rect 480253 371452 480300 371456
rect 480364 371454 480410 371514
rect 480364 371452 480370 371454
rect 480253 371451 480319 371452
rect 107561 371380 107627 371381
rect 106958 371316 106964 371380
rect 107028 371316 107034 371380
rect 107510 371378 107516 371380
rect 107470 371318 107516 371378
rect 107580 371376 107627 371380
rect 107622 371320 107627 371376
rect 107510 371316 107516 371318
rect 107580 371316 107627 371320
rect 115790 371316 115796 371380
rect 115860 371378 115866 371380
rect 219433 371378 219499 371381
rect 220721 371378 220787 371381
rect 115860 371376 220787 371378
rect 115860 371320 219438 371376
rect 219494 371320 220726 371376
rect 220782 371320 220787 371376
rect 115860 371318 220787 371320
rect 115860 371316 115866 371318
rect 106966 371242 107026 371316
rect 107561 371315 107627 371316
rect 219433 371315 219499 371318
rect 220721 371315 220787 371318
rect 249793 371378 249859 371381
rect 249926 371378 249932 371380
rect 249793 371376 249932 371378
rect 249793 371320 249798 371376
rect 249854 371320 249932 371376
rect 249793 371318 249932 371320
rect 249793 371315 249859 371318
rect 249926 371316 249932 371318
rect 249996 371316 250002 371380
rect 252553 371378 252619 371381
rect 253606 371378 253612 371380
rect 252553 371376 253612 371378
rect 252553 371320 252558 371376
rect 252614 371320 253612 371376
rect 252553 371318 253612 371320
rect 252553 371315 252619 371318
rect 253606 371316 253612 371318
rect 253676 371316 253682 371380
rect 255313 371378 255379 371381
rect 256182 371378 256188 371380
rect 255313 371376 256188 371378
rect 255313 371320 255318 371376
rect 255374 371320 256188 371376
rect 255313 371318 256188 371320
rect 255313 371315 255379 371318
rect 256182 371316 256188 371318
rect 256252 371316 256258 371380
rect 258165 371378 258231 371381
rect 258390 371378 258396 371380
rect 258165 371376 258396 371378
rect 258165 371320 258170 371376
rect 258226 371320 258396 371376
rect 258165 371318 258396 371320
rect 258165 371315 258231 371318
rect 258390 371316 258396 371318
rect 258460 371316 258466 371380
rect 260833 371378 260899 371381
rect 263593 371380 263659 371381
rect 260966 371378 260972 371380
rect 260833 371376 260972 371378
rect 260833 371320 260838 371376
rect 260894 371320 260972 371376
rect 260833 371318 260972 371320
rect 260833 371315 260899 371318
rect 260966 371316 260972 371318
rect 261036 371316 261042 371380
rect 263542 371316 263548 371380
rect 263612 371378 263659 371380
rect 266353 371378 266419 371381
rect 267733 371380 267799 371381
rect 267038 371378 267044 371380
rect 263612 371376 263704 371378
rect 263654 371320 263704 371376
rect 263612 371318 263704 371320
rect 266353 371376 267044 371378
rect 266353 371320 266358 371376
rect 266414 371320 267044 371376
rect 266353 371318 267044 371320
rect 263612 371316 263659 371318
rect 263593 371315 263659 371316
rect 266353 371315 266419 371318
rect 267038 371316 267044 371318
rect 267108 371316 267114 371380
rect 267733 371376 267780 371380
rect 267844 371378 267850 371380
rect 276013 371378 276079 371381
rect 276238 371378 276244 371380
rect 267733 371320 267738 371376
rect 267733 371316 267780 371320
rect 267844 371318 267890 371378
rect 276013 371376 276244 371378
rect 276013 371320 276018 371376
rect 276074 371320 276244 371376
rect 276013 371318 276244 371320
rect 267844 371316 267850 371318
rect 267733 371315 267799 371316
rect 276013 371315 276079 371318
rect 276238 371316 276244 371318
rect 276308 371316 276314 371380
rect 277761 371378 277827 371381
rect 278262 371378 278268 371380
rect 277761 371376 278268 371378
rect 277761 371320 277766 371376
rect 277822 371320 278268 371376
rect 277761 371318 278268 371320
rect 277761 371315 277827 371318
rect 278262 371316 278268 371318
rect 278332 371316 278338 371380
rect 280153 371378 280219 371381
rect 280286 371378 280292 371380
rect 280153 371376 280292 371378
rect 280153 371320 280158 371376
rect 280214 371320 280292 371376
rect 280153 371318 280292 371320
rect 280153 371315 280219 371318
rect 280286 371316 280292 371318
rect 280356 371316 280362 371380
rect 285673 371378 285739 371381
rect 285806 371378 285812 371380
rect 285673 371376 285812 371378
rect 285673 371320 285678 371376
rect 285734 371320 285812 371376
rect 285673 371318 285812 371320
rect 285673 371315 285739 371318
rect 285806 371316 285812 371318
rect 285876 371316 285882 371380
rect 287237 371378 287303 371381
rect 287646 371378 287652 371380
rect 287237 371376 287652 371378
rect 287237 371320 287242 371376
rect 287298 371320 287652 371376
rect 287237 371318 287652 371320
rect 287237 371315 287303 371318
rect 287646 371316 287652 371318
rect 287716 371316 287722 371380
rect 289813 371378 289879 371381
rect 290590 371378 290596 371380
rect 289813 371376 290596 371378
rect 289813 371320 289818 371376
rect 289874 371320 290596 371376
rect 289813 371318 290596 371320
rect 289813 371315 289879 371318
rect 290590 371316 290596 371318
rect 290660 371316 290666 371380
rect 292573 371378 292639 371381
rect 295333 371380 295399 371381
rect 298093 371380 298159 371381
rect 292798 371378 292804 371380
rect 292573 371376 292804 371378
rect 292573 371320 292578 371376
rect 292634 371320 292804 371376
rect 292573 371318 292804 371320
rect 292573 371315 292639 371318
rect 292798 371316 292804 371318
rect 292868 371316 292874 371380
rect 295333 371378 295380 371380
rect 295288 371376 295380 371378
rect 295288 371320 295338 371376
rect 295288 371318 295380 371320
rect 295333 371316 295380 371318
rect 295444 371316 295450 371380
rect 298093 371378 298140 371380
rect 298048 371376 298140 371378
rect 298048 371320 298098 371376
rect 298048 371318 298140 371320
rect 298093 371316 298140 371318
rect 298204 371316 298210 371380
rect 302233 371378 302299 371381
rect 302918 371378 302924 371380
rect 302233 371376 302924 371378
rect 302233 371320 302238 371376
rect 302294 371320 302924 371376
rect 302233 371318 302924 371320
rect 295333 371315 295399 371316
rect 298093 371315 298159 371316
rect 302233 371315 302299 371318
rect 302918 371316 302924 371318
rect 302988 371316 302994 371380
rect 307753 371378 307819 371381
rect 322933 371380 322999 371381
rect 308622 371378 308628 371380
rect 307753 371376 308628 371378
rect 307753 371320 307758 371376
rect 307814 371320 308628 371376
rect 307753 371318 308628 371320
rect 307753 371315 307819 371318
rect 308622 371316 308628 371318
rect 308692 371316 308698 371380
rect 322933 371378 322980 371380
rect 322888 371376 322980 371378
rect 322888 371320 322938 371376
rect 322888 371318 322980 371320
rect 322933 371316 322980 371318
rect 323044 371316 323050 371380
rect 343081 371378 343147 371381
rect 343449 371380 343515 371381
rect 343214 371378 343220 371380
rect 343081 371376 343220 371378
rect 343081 371320 343086 371376
rect 343142 371320 343220 371376
rect 343081 371318 343220 371320
rect 322933 371315 322999 371316
rect 343081 371315 343147 371318
rect 343214 371316 343220 371318
rect 343284 371316 343290 371380
rect 343398 371316 343404 371380
rect 343468 371378 343515 371380
rect 396073 371378 396139 371381
rect 402973 371380 403039 371381
rect 396574 371378 396580 371380
rect 343468 371376 343560 371378
rect 343510 371320 343560 371376
rect 343468 371318 343560 371320
rect 396073 371376 396580 371378
rect 396073 371320 396078 371376
rect 396134 371320 396580 371376
rect 396073 371318 396580 371320
rect 343468 371316 343515 371318
rect 343449 371315 343515 371316
rect 396073 371315 396139 371318
rect 396574 371316 396580 371318
rect 396644 371316 396650 371380
rect 402973 371376 403020 371380
rect 403084 371378 403090 371380
rect 405733 371378 405799 371381
rect 406142 371378 406148 371380
rect 402973 371320 402978 371376
rect 402973 371316 403020 371320
rect 403084 371318 403130 371378
rect 405733 371376 406148 371378
rect 405733 371320 405738 371376
rect 405794 371320 406148 371376
rect 405733 371318 406148 371320
rect 403084 371316 403090 371318
rect 402973 371315 403039 371316
rect 405733 371315 405799 371318
rect 406142 371316 406148 371318
rect 406212 371316 406218 371380
rect 412633 371378 412699 371381
rect 412766 371378 412772 371380
rect 412633 371376 412772 371378
rect 412633 371320 412638 371376
rect 412694 371320 412772 371376
rect 412633 371318 412772 371320
rect 412633 371315 412699 371318
rect 412766 371316 412772 371318
rect 412836 371316 412842 371380
rect 413185 371378 413251 371381
rect 414013 371380 414079 371381
rect 413686 371378 413692 371380
rect 413185 371376 413692 371378
rect 413185 371320 413190 371376
rect 413246 371320 413692 371376
rect 413185 371318 413692 371320
rect 413185 371315 413251 371318
rect 413686 371316 413692 371318
rect 413756 371316 413762 371380
rect 414013 371378 414060 371380
rect 413968 371376 414060 371378
rect 413968 371320 414018 371376
rect 413968 371318 414060 371320
rect 414013 371316 414060 371318
rect 414124 371316 414130 371380
rect 415393 371378 415459 371381
rect 416773 371380 416839 371381
rect 415526 371378 415532 371380
rect 415393 371376 415532 371378
rect 415393 371320 415398 371376
rect 415454 371320 415532 371376
rect 415393 371318 415532 371320
rect 414013 371315 414079 371316
rect 415393 371315 415459 371318
rect 415526 371316 415532 371318
rect 415596 371316 415602 371380
rect 416773 371378 416820 371380
rect 416728 371376 416820 371378
rect 416728 371320 416778 371376
rect 416728 371318 416820 371320
rect 416773 371316 416820 371318
rect 416884 371316 416890 371380
rect 418153 371378 418219 371381
rect 418286 371378 418292 371380
rect 418153 371376 418292 371378
rect 418153 371320 418158 371376
rect 418214 371320 418292 371376
rect 418153 371318 418292 371320
rect 416773 371315 416839 371316
rect 418153 371315 418219 371318
rect 418286 371316 418292 371318
rect 418356 371316 418362 371380
rect 419533 371378 419599 371381
rect 422293 371380 422359 371381
rect 420310 371378 420316 371380
rect 419533 371376 420316 371378
rect 419533 371320 419538 371376
rect 419594 371320 420316 371376
rect 419533 371318 420316 371320
rect 419533 371315 419599 371318
rect 420310 371316 420316 371318
rect 420380 371316 420386 371380
rect 422293 371376 422340 371380
rect 422404 371378 422410 371380
rect 425053 371378 425119 371381
rect 425646 371378 425652 371380
rect 422293 371320 422298 371376
rect 422293 371316 422340 371320
rect 422404 371318 422450 371378
rect 425053 371376 425652 371378
rect 425053 371320 425058 371376
rect 425114 371320 425652 371376
rect 425053 371318 425652 371320
rect 422404 371316 422410 371318
rect 422293 371315 422359 371316
rect 425053 371315 425119 371318
rect 425646 371316 425652 371318
rect 425716 371316 425722 371380
rect 427905 371378 427971 371381
rect 428590 371378 428596 371380
rect 427905 371376 428596 371378
rect 427905 371320 427910 371376
rect 427966 371320 428596 371376
rect 427905 371318 428596 371320
rect 427905 371315 427971 371318
rect 428590 371316 428596 371318
rect 428660 371316 428666 371380
rect 431953 371378 432019 371381
rect 432086 371378 432092 371380
rect 431953 371376 432092 371378
rect 431953 371320 431958 371376
rect 432014 371320 432092 371376
rect 431953 371318 432092 371320
rect 431953 371315 432019 371318
rect 432086 371316 432092 371318
rect 432156 371316 432162 371380
rect 434713 371378 434779 371381
rect 434846 371378 434852 371380
rect 434713 371376 434852 371378
rect 434713 371320 434718 371376
rect 434774 371320 434852 371376
rect 434713 371318 434852 371320
rect 434713 371315 434779 371318
rect 434846 371316 434852 371318
rect 434916 371316 434922 371380
rect 436093 371378 436159 371381
rect 460933 371380 460999 371381
rect 436318 371378 436324 371380
rect 436093 371376 436324 371378
rect 436093 371320 436098 371376
rect 436154 371320 436324 371376
rect 436093 371318 436324 371320
rect 436093 371315 436159 371318
rect 436318 371316 436324 371318
rect 436388 371316 436394 371380
rect 460933 371376 460980 371380
rect 461044 371378 461050 371380
rect 467833 371378 467899 371381
rect 473353 371380 473419 371381
rect 467966 371378 467972 371380
rect 460933 371320 460938 371376
rect 460933 371316 460980 371320
rect 461044 371318 461090 371378
rect 467833 371376 467972 371378
rect 467833 371320 467838 371376
rect 467894 371320 467972 371376
rect 467833 371318 467972 371320
rect 461044 371316 461050 371318
rect 460933 371315 460999 371316
rect 467833 371315 467899 371318
rect 467966 371316 467972 371318
rect 468036 371316 468042 371380
rect 473302 371316 473308 371380
rect 473372 371378 473419 371380
rect 483013 371378 483079 371381
rect 483238 371378 483244 371380
rect 473372 371376 473464 371378
rect 473414 371320 473464 371376
rect 473372 371318 473464 371320
rect 483013 371376 483244 371378
rect 483013 371320 483018 371376
rect 483074 371320 483244 371376
rect 483013 371318 483244 371320
rect 473372 371316 473419 371318
rect 473353 371315 473419 371316
rect 483013 371315 483079 371318
rect 483238 371316 483244 371318
rect 483308 371316 483314 371380
rect 106966 371182 200130 371242
rect 200070 370970 200130 371182
rect 216990 370970 216996 370972
rect 200070 370910 216996 370970
rect 216990 370908 216996 370910
rect 217060 370970 217066 370972
rect 217542 370970 217548 370972
rect 217060 370910 217548 370970
rect 217060 370908 217066 370910
rect 217542 370908 217548 370910
rect 217612 370908 217618 370972
rect 214782 369820 214788 369884
rect 214852 369882 214858 369884
rect 215201 369882 215267 369885
rect 214852 369880 215267 369882
rect 214852 369824 215206 369880
rect 215262 369824 215267 369880
rect 214852 369822 215267 369824
rect 214852 369820 214858 369822
rect 215201 369819 215267 369822
rect 104617 369746 104683 369749
rect 215661 369746 215727 369749
rect 104617 369744 215727 369746
rect 104617 369688 104622 369744
rect 104678 369688 215666 369744
rect 215722 369688 215727 369744
rect 104617 369686 215727 369688
rect 104617 369683 104683 369686
rect 215661 369683 215727 369686
rect 105905 369610 105971 369613
rect 215385 369610 215451 369613
rect 105905 369608 215451 369610
rect 105905 369552 105910 369608
rect 105966 369552 215390 369608
rect 215446 369552 215451 369608
rect 105905 369550 215451 369552
rect 105905 369547 105971 369550
rect 215385 369547 215451 369550
rect 208945 369202 209011 369205
rect 209262 369202 209268 369204
rect 208945 369200 209268 369202
rect 208945 369144 208950 369200
rect 209006 369144 209268 369200
rect 208945 369142 209268 369144
rect 208945 369139 209011 369142
rect 209262 369140 209268 369142
rect 209332 369140 209338 369204
rect 212574 369140 212580 369204
rect 212644 369202 212650 369204
rect 213821 369202 213887 369205
rect 212644 369200 213887 369202
rect 212644 369144 213826 369200
rect 213882 369144 213887 369200
rect 212644 369142 213887 369144
rect 212644 369140 212650 369142
rect 213821 369139 213887 369142
rect 376937 368524 377003 368525
rect 376886 368522 376892 368524
rect 376846 368462 376892 368522
rect 376956 368520 377003 368524
rect 376998 368464 377003 368520
rect 376886 368460 376892 368462
rect 376956 368460 377003 368464
rect 376937 368459 377003 368460
rect 583520 364972 584960 365212
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 179638 355268 179644 355332
rect 179708 355330 179714 355332
rect 179781 355330 179847 355333
rect 179708 355328 179847 355330
rect 179708 355272 179786 355328
rect 179842 355272 179847 355328
rect 179708 355270 179847 355272
rect 179708 355268 179714 355270
rect 179781 355267 179847 355270
rect 190862 355268 190868 355332
rect 190932 355330 190938 355332
rect 191373 355330 191439 355333
rect 190932 355328 191439 355330
rect 190932 355272 191378 355328
rect 191434 355272 191439 355328
rect 190932 355270 191439 355272
rect 190932 355268 190938 355270
rect 191373 355267 191439 355270
rect 339718 354996 339724 355060
rect 339788 355058 339794 355060
rect 340045 355058 340111 355061
rect 339788 355056 340111 355058
rect 339788 355000 340050 355056
rect 340106 355000 340111 355056
rect 339788 354998 340111 355000
rect 339788 354996 339794 354998
rect 340045 354995 340111 354998
rect 350942 354996 350948 355060
rect 351012 355058 351018 355060
rect 351729 355058 351795 355061
rect 351012 355056 351795 355058
rect 351012 355000 351734 355056
rect 351790 355000 351795 355056
rect 351012 354998 351795 355000
rect 351012 354996 351018 354998
rect 351729 354995 351795 354998
rect 498510 354996 498516 355060
rect 498580 355058 498586 355060
rect 498837 355058 498903 355061
rect 498580 355056 498903 355058
rect 498580 355000 498842 355056
rect 498898 355000 498903 355056
rect 498580 354998 498903 355000
rect 498580 354996 498586 354998
rect 498837 354995 498903 354998
rect 499798 354860 499804 354924
rect 499868 354922 499874 354924
rect 500861 354922 500927 354925
rect 499868 354920 500927 354922
rect 499868 354864 500866 354920
rect 500922 354864 500927 354920
rect 499868 354862 500927 354864
rect 499868 354860 499874 354862
rect 500861 354859 500927 354862
rect 178585 354788 178651 354789
rect 338113 354788 338179 354789
rect 510889 354788 510955 354789
rect 178534 354786 178540 354788
rect 178494 354726 178540 354786
rect 178604 354784 178651 354788
rect 338062 354786 338068 354788
rect 178646 354728 178651 354784
rect 178534 354724 178540 354726
rect 178604 354724 178651 354728
rect 338022 354726 338068 354786
rect 338132 354784 338179 354788
rect 510838 354786 510844 354788
rect 338174 354728 338179 354784
rect 338062 354724 338068 354726
rect 338132 354724 338179 354728
rect 510798 354726 510844 354786
rect 510908 354784 510955 354788
rect 510950 354728 510955 354784
rect 510838 354724 510844 354726
rect 510908 354724 510955 354728
rect 178585 354723 178651 354724
rect 338113 354723 338179 354724
rect 510889 354723 510955 354724
rect 580349 351930 580415 351933
rect 583520 351930 584960 352020
rect 580349 351928 584960 351930
rect 580349 351872 580354 351928
rect 580410 351872 584960 351928
rect 580349 351870 584960 351872
rect 580349 351867 580415 351870
rect 583520 351780 584960 351870
rect 198733 349618 198799 349621
rect 199009 349618 199075 349621
rect 358905 349618 358971 349621
rect 196558 349616 199075 349618
rect 196558 349560 198738 349616
rect 198794 349560 199014 349616
rect 199070 349560 199075 349616
rect 196558 349558 199075 349560
rect 196558 349190 196618 349558
rect 198733 349555 198799 349558
rect 199009 349555 199075 349558
rect 356562 349616 358971 349618
rect 356562 349560 358910 349616
rect 358966 349560 358971 349616
rect 356562 349558 358971 349560
rect 356562 349190 356622 349558
rect 358905 349555 358971 349558
rect 518893 349210 518959 349213
rect 516558 349208 518959 349210
rect 516558 349152 518898 349208
rect 518954 349152 518959 349208
rect 516558 349150 518959 349152
rect 518893 349147 518959 349150
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580257 325274 580323 325277
rect 583520 325274 584960 325364
rect 580257 325272 584960 325274
rect 580257 325216 580262 325272
rect 580318 325216 584960 325272
rect 580257 325214 584960 325216
rect 580257 325211 580323 325214
rect 583520 325124 584960 325214
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect 217777 307730 217843 307733
rect 217961 307730 218027 307733
rect 217777 307728 218027 307730
rect 217777 307672 217782 307728
rect 217838 307672 217966 307728
rect 218022 307672 218027 307728
rect 217777 307670 218027 307672
rect 217777 307667 217843 307670
rect 217961 307667 218027 307670
rect 57421 306914 57487 306917
rect 217777 306914 217843 306917
rect 219390 306914 220064 306924
rect 57421 306912 60062 306914
rect 57421 306856 57426 306912
rect 57482 306856 60062 306912
rect 57421 306854 60062 306856
rect 217777 306912 220064 306914
rect 217777 306856 217782 306912
rect 217838 306864 220064 306912
rect 377029 306914 377095 306917
rect 379470 306914 380052 306924
rect 377029 306912 380052 306914
rect 217838 306856 219450 306864
rect 217777 306854 219450 306856
rect 377029 306856 377034 306912
rect 377090 306864 380052 306912
rect 377090 306856 379530 306864
rect 377029 306854 379530 306856
rect 57421 306851 57487 306854
rect 217777 306851 217843 306854
rect 377029 306851 377095 306854
rect -960 306234 480 306324
rect -960 306174 674 306234
rect -960 306098 480 306174
rect 614 306098 674 306174
rect -960 306084 674 306098
rect 246 306038 674 306084
rect 246 305554 306 306038
rect 57881 305962 57947 305965
rect 217685 305962 217751 305965
rect 219390 305962 220064 305972
rect 57881 305960 60062 305962
rect 57881 305904 57886 305960
rect 57942 305904 60062 305960
rect 57881 305902 60062 305904
rect 217685 305960 220064 305962
rect 217685 305904 217690 305960
rect 217746 305912 220064 305960
rect 377765 305962 377831 305965
rect 379470 305962 380052 305972
rect 377765 305960 380052 305962
rect 217746 305904 219450 305912
rect 217685 305902 219450 305904
rect 377765 305904 377770 305960
rect 377826 305912 380052 305960
rect 377826 305904 379530 305912
rect 377765 305902 379530 305904
rect 57881 305899 57947 305902
rect 217685 305899 217751 305902
rect 377765 305899 377831 305902
rect 246 305494 6930 305554
rect 6870 305010 6930 305494
rect 54334 305010 54340 305012
rect 6870 304950 54340 305010
rect 54334 304948 54340 304950
rect 54404 304948 54410 305012
rect 57145 305010 57211 305013
rect 57881 305010 57947 305013
rect 57145 305008 57947 305010
rect 57145 304952 57150 305008
rect 57206 304952 57886 305008
rect 57942 304952 57947 305008
rect 57145 304950 57947 304952
rect 57145 304947 57211 304950
rect 57881 304947 57947 304950
rect 377305 305010 377371 305013
rect 377765 305010 377831 305013
rect 377305 305008 377831 305010
rect 377305 304952 377310 305008
rect 377366 304952 377770 305008
rect 377826 304952 377831 305008
rect 377305 304950 377831 304952
rect 377305 304947 377371 304950
rect 377765 304947 377831 304950
rect 216949 303786 217015 303789
rect 217409 303786 217475 303789
rect 219390 303786 220064 303796
rect 216949 303784 220064 303786
rect 56685 303650 56751 303653
rect 57789 303650 57855 303653
rect 60002 303650 60062 303766
rect 216949 303728 216954 303784
rect 217010 303728 217414 303784
rect 217470 303736 220064 303784
rect 379470 303736 380052 303796
rect 217470 303728 219450 303736
rect 216949 303726 219450 303728
rect 216949 303723 217015 303726
rect 217409 303723 217475 303726
rect 56685 303648 60062 303650
rect 56685 303592 56690 303648
rect 56746 303592 57794 303648
rect 57850 303592 60062 303648
rect 56685 303590 60062 303592
rect 377029 303650 377095 303653
rect 377857 303650 377923 303653
rect 379470 303650 379530 303736
rect 377029 303648 379530 303650
rect 377029 303592 377034 303648
rect 377090 303592 377862 303648
rect 377918 303592 379530 303648
rect 377029 303590 379530 303592
rect 56685 303587 56751 303590
rect 57789 303587 57855 303590
rect 377029 303587 377095 303590
rect 377857 303587 377923 303590
rect 216857 302834 216923 302837
rect 217501 302834 217567 302837
rect 219390 302834 220064 302844
rect 216857 302832 220064 302834
rect 56777 302290 56843 302293
rect 57605 302290 57671 302293
rect 60002 302290 60062 302814
rect 216857 302776 216862 302832
rect 216918 302776 217506 302832
rect 217562 302784 220064 302832
rect 377489 302834 377555 302837
rect 379470 302834 380052 302844
rect 377489 302832 380052 302834
rect 217562 302776 219450 302784
rect 216857 302774 219450 302776
rect 377489 302776 377494 302832
rect 377550 302784 380052 302832
rect 377550 302776 379530 302784
rect 377489 302774 379530 302776
rect 216857 302771 216923 302774
rect 217501 302771 217567 302774
rect 377489 302771 377555 302774
rect 56777 302288 60062 302290
rect 56777 302232 56782 302288
rect 56838 302232 57610 302288
rect 57666 302232 60062 302288
rect 56777 302230 60062 302232
rect 56777 302227 56843 302230
rect 57605 302227 57671 302230
rect 57513 301338 57579 301341
rect 57513 301336 60062 301338
rect 57513 301280 57518 301336
rect 57574 301280 60062 301336
rect 57513 301278 60062 301280
rect 57513 301275 57579 301278
rect 60002 301046 60062 301278
rect 217041 301066 217107 301069
rect 217317 301066 217383 301069
rect 219390 301066 220064 301076
rect 217041 301064 220064 301066
rect 217041 301008 217046 301064
rect 217102 301008 217322 301064
rect 217378 301016 220064 301064
rect 377213 301066 377279 301069
rect 379470 301066 380052 301076
rect 377213 301064 380052 301066
rect 217378 301008 219450 301016
rect 217041 301006 219450 301008
rect 377213 301008 377218 301064
rect 377274 301016 380052 301064
rect 377274 301008 379530 301016
rect 377213 301006 379530 301008
rect 217041 301003 217107 301006
rect 217317 301003 217383 301006
rect 377213 301003 377279 301006
rect 57053 300522 57119 300525
rect 57697 300522 57763 300525
rect 57053 300520 60062 300522
rect 57053 300464 57058 300520
rect 57114 300464 57702 300520
rect 57758 300464 60062 300520
rect 57053 300462 60062 300464
rect 57053 300459 57119 300462
rect 57697 300459 57763 300462
rect 60002 299958 60062 300462
rect 217225 299978 217291 299981
rect 219390 299978 220064 299988
rect 217225 299976 220064 299978
rect 217225 299920 217230 299976
rect 217286 299928 220064 299976
rect 377581 299978 377647 299981
rect 377765 299978 377831 299981
rect 379470 299978 380052 299988
rect 377581 299976 380052 299978
rect 217286 299920 219450 299928
rect 217225 299918 219450 299920
rect 377581 299920 377586 299976
rect 377642 299920 377770 299976
rect 377826 299928 380052 299976
rect 377826 299920 379530 299928
rect 377581 299918 379530 299920
rect 217225 299915 217291 299918
rect 377581 299915 377647 299918
rect 377765 299915 377831 299918
rect 216765 299434 216831 299437
rect 217593 299434 217659 299437
rect 216765 299432 217659 299434
rect 216765 299376 216770 299432
rect 216826 299376 217598 299432
rect 217654 299376 217659 299432
rect 216765 299374 217659 299376
rect 216765 299371 216831 299374
rect 217593 299371 217659 299374
rect 583520 298604 584960 298844
rect 57513 298210 57579 298213
rect 217593 298210 217659 298213
rect 219390 298210 220064 298220
rect 57513 298208 60062 298210
rect 57513 298152 57518 298208
rect 57574 298152 60062 298208
rect 57513 298150 60062 298152
rect 217593 298208 220064 298210
rect 217593 298152 217598 298208
rect 217654 298160 220064 298208
rect 377857 298210 377923 298213
rect 379470 298210 380052 298220
rect 377857 298208 380052 298210
rect 217654 298152 219450 298160
rect 217593 298150 219450 298152
rect 377857 298152 377862 298208
rect 377918 298160 380052 298208
rect 377918 298152 379530 298160
rect 377857 298150 379530 298152
rect 57513 298147 57579 298150
rect 217593 298147 217659 298150
rect 377857 298147 377923 298150
rect -960 293028 480 293268
rect 199009 289778 199075 289781
rect 199745 289778 199811 289781
rect 196558 289776 199811 289778
rect 196558 289720 199014 289776
rect 199070 289720 199750 289776
rect 199806 289720 199811 289776
rect 196558 289718 199811 289720
rect 196558 289350 196618 289718
rect 199009 289715 199075 289718
rect 199745 289715 199811 289718
rect 359089 289370 359155 289373
rect 518985 289370 519051 289373
rect 519537 289370 519603 289373
rect 356562 289368 359155 289370
rect 356562 289312 359094 289368
rect 359150 289312 359155 289368
rect 356562 289310 359155 289312
rect 516558 289368 519603 289370
rect 516558 289312 518990 289368
rect 519046 289312 519542 289368
rect 519598 289312 519603 289368
rect 516558 289310 519603 289312
rect 359089 289307 359155 289310
rect 518985 289307 519051 289310
rect 519537 289307 519603 289310
rect 198825 288418 198891 288421
rect 199377 288418 199443 288421
rect 358997 288418 359063 288421
rect 359549 288418 359615 288421
rect 198825 288416 199443 288418
rect 198825 288360 198830 288416
rect 198886 288360 199382 288416
rect 199438 288360 199443 288416
rect 198825 288358 199443 288360
rect 198825 288355 198891 288358
rect 199377 288355 199443 288358
rect 356562 288416 359615 288418
rect 356562 288360 359002 288416
rect 359058 288360 359554 288416
rect 359610 288360 359615 288416
rect 356562 288358 359615 288360
rect 198825 287738 198891 287741
rect 196558 287736 198891 287738
rect 196558 287680 198830 287736
rect 198886 287680 198891 287736
rect 356562 287718 356622 288358
rect 358997 288355 359063 288358
rect 359549 288355 359615 288358
rect 518985 288418 519051 288421
rect 519169 288418 519235 288421
rect 518985 288416 519235 288418
rect 518985 288360 518990 288416
rect 519046 288360 519174 288416
rect 519230 288360 519235 288416
rect 518985 288358 519235 288360
rect 518985 288355 519051 288358
rect 519169 288355 519235 288358
rect 196558 287678 198891 287680
rect 198825 287675 198891 287678
rect 516558 287194 516618 287718
rect 518985 287194 519051 287197
rect 516558 287192 519051 287194
rect 516558 287136 518990 287192
rect 519046 287136 519051 287192
rect 516558 287134 519051 287136
rect 518985 287131 519051 287134
rect 199561 286378 199627 286381
rect 359273 286378 359339 286381
rect 196558 286376 199627 286378
rect 196558 286320 199566 286376
rect 199622 286320 199627 286376
rect 196558 286318 199627 286320
rect 356562 286376 359339 286378
rect 356562 286320 359278 286376
rect 359334 286320 359339 286376
rect 356562 286318 359339 286320
rect 199561 286315 199627 286318
rect 359273 286315 359339 286318
rect 516558 285834 516618 286358
rect 519261 285834 519327 285837
rect 519629 285834 519695 285837
rect 516558 285832 519695 285834
rect 516558 285776 519266 285832
rect 519322 285776 519634 285832
rect 519690 285776 519695 285832
rect 516558 285774 519695 285776
rect 519261 285771 519327 285774
rect 519629 285771 519695 285774
rect 583520 285276 584960 285516
rect 199101 284882 199167 284885
rect 359457 284882 359523 284885
rect 519353 284882 519419 284885
rect 520181 284882 520247 284885
rect 196558 284880 199167 284882
rect 196558 284824 199106 284880
rect 199162 284824 199167 284880
rect 196558 284822 199167 284824
rect 356562 284880 359523 284882
rect 356562 284824 359462 284880
rect 359518 284824 359523 284880
rect 356562 284822 359523 284824
rect 516558 284880 520247 284882
rect 516558 284824 519358 284880
rect 519414 284824 520186 284880
rect 520242 284824 520247 284880
rect 516558 284822 520247 284824
rect 199101 284819 199167 284822
rect 359457 284819 359523 284822
rect 519353 284819 519419 284822
rect 520181 284819 520247 284822
rect 519077 284202 519143 284205
rect 516558 284200 519143 284202
rect 516558 284144 519082 284200
rect 519138 284144 519143 284200
rect 516558 284142 519143 284144
rect 516558 283638 516618 284142
rect 519077 284139 519143 284142
rect 196558 283114 196618 283638
rect 198917 283114 198983 283117
rect 199653 283114 199719 283117
rect 196558 283112 199719 283114
rect 196558 283056 198922 283112
rect 198978 283056 199658 283112
rect 199714 283056 199719 283112
rect 196558 283054 199719 283056
rect 356562 283114 356622 283638
rect 358997 283114 359063 283117
rect 359181 283114 359247 283117
rect 356562 283112 359247 283114
rect 356562 283056 359002 283112
rect 359058 283056 359186 283112
rect 359242 283056 359247 283112
rect 356562 283054 359247 283056
rect 198917 283051 198983 283054
rect 199653 283051 199719 283054
rect 358997 283051 359063 283054
rect 359181 283051 359247 283054
rect -960 279972 480 280212
rect 58709 279986 58775 279989
rect 216673 279986 216739 279989
rect 219390 279986 220064 279996
rect 58709 279984 60062 279986
rect 58709 279928 58714 279984
rect 58770 279928 60062 279984
rect 58709 279926 60062 279928
rect 216673 279984 220064 279986
rect 216673 279928 216678 279984
rect 216734 279936 220064 279984
rect 216734 279928 219450 279936
rect 216673 279926 219450 279928
rect 58709 279923 58775 279926
rect 216673 279923 216739 279926
rect 359774 279924 359780 279988
rect 359844 279986 359850 279988
rect 379470 279986 380052 279996
rect 359844 279936 380052 279986
rect 359844 279926 379530 279936
rect 359844 279924 359850 279926
rect 57237 278762 57303 278765
rect 57881 278762 57947 278765
rect 57237 278760 60062 278762
rect 57237 278704 57242 278760
rect 57298 278704 57886 278760
rect 57942 278704 60062 278760
rect 57237 278702 60062 278704
rect 57237 278699 57303 278702
rect 57881 278699 57947 278702
rect 60002 278334 60062 278702
rect 216949 278354 217015 278357
rect 219390 278354 220064 278364
rect 216949 278352 220064 278354
rect 216949 278296 216954 278352
rect 217010 278304 220064 278352
rect 376845 278354 376911 278357
rect 379470 278354 380052 278364
rect 376845 278352 380052 278354
rect 217010 278296 219450 278304
rect 216949 278294 219450 278296
rect 376845 278296 376850 278352
rect 376906 278304 380052 278352
rect 376906 278296 379530 278304
rect 376845 278294 379530 278296
rect 216949 278291 217015 278294
rect 376845 278291 376911 278294
rect 58801 278082 58867 278085
rect 216673 278082 216739 278085
rect 219390 278082 220064 278092
rect 58801 278080 60062 278082
rect 58801 278024 58806 278080
rect 58862 278024 60062 278080
rect 58801 278022 60062 278024
rect 216673 278080 220064 278082
rect 216673 278024 216678 278080
rect 216734 278032 220064 278080
rect 376753 278082 376819 278085
rect 379470 278082 380052 278092
rect 376753 278080 380052 278082
rect 216734 278024 219450 278032
rect 216673 278022 219450 278024
rect 376753 278024 376758 278080
rect 376814 278032 380052 278080
rect 376814 278024 379530 278032
rect 376753 278022 379530 278024
rect 58801 278019 58867 278022
rect 216673 278019 216739 278022
rect 376753 278019 376819 278022
rect 580349 272234 580415 272237
rect 583520 272234 584960 272324
rect 580349 272232 584960 272234
rect 580349 272176 580354 272232
rect 580410 272176 584960 272232
rect 580349 272174 584960 272176
rect 580349 272171 580415 272174
rect 583520 272084 584960 272174
rect 110965 269924 111031 269925
rect 148501 269924 148567 269925
rect 110965 269920 111006 269924
rect 111070 269922 111076 269924
rect 110965 269864 110970 269920
rect 110965 269860 111006 269864
rect 111070 269862 111122 269922
rect 148501 269920 148542 269924
rect 148606 269922 148612 269924
rect 148501 269864 148506 269920
rect 111070 269860 111076 269862
rect 148501 269860 148542 269864
rect 148606 269862 148658 269922
rect 148606 269860 148612 269862
rect 110965 269859 111031 269860
rect 148501 269859 148567 269860
rect 133413 269788 133479 269789
rect 135897 269788 135963 269789
rect 138473 269788 138539 269789
rect 140865 269788 140931 269789
rect 250713 269788 250779 269789
rect 416037 269788 416103 269789
rect 425237 269788 425303 269789
rect 433333 269788 433399 269789
rect 133413 269784 133446 269788
rect 133510 269786 133516 269788
rect 135888 269786 135894 269788
rect 133413 269728 133418 269784
rect 133413 269724 133446 269728
rect 133510 269726 133570 269786
rect 135806 269726 135894 269786
rect 133510 269724 133516 269726
rect 135888 269724 135894 269726
rect 135958 269724 135964 269788
rect 138472 269724 138478 269788
rect 138542 269786 138548 269788
rect 138542 269726 138630 269786
rect 140865 269784 140926 269788
rect 140865 269728 140870 269784
rect 138542 269724 138548 269726
rect 140865 269724 140926 269728
rect 140990 269786 140996 269788
rect 140990 269726 141022 269786
rect 250713 269784 250742 269788
rect 250806 269786 250812 269788
rect 250713 269728 250718 269784
rect 140990 269724 140996 269726
rect 250713 269724 250742 269728
rect 250806 269726 250870 269786
rect 416037 269784 416046 269788
rect 416110 269786 416116 269788
rect 416037 269728 416042 269784
rect 250806 269724 250812 269726
rect 416037 269724 416046 269728
rect 416110 269726 416194 269786
rect 425237 269784 425294 269788
rect 425358 269786 425364 269788
rect 433312 269786 433318 269788
rect 425237 269728 425242 269784
rect 416110 269724 416116 269726
rect 425237 269724 425294 269728
rect 425358 269726 425394 269786
rect 433242 269726 433318 269786
rect 433382 269784 433399 269788
rect 433394 269728 433399 269784
rect 425358 269724 425364 269726
rect 433312 269724 433318 269726
rect 433382 269724 433399 269728
rect 133413 269723 133479 269724
rect 135897 269723 135963 269724
rect 138473 269723 138539 269724
rect 140865 269723 140931 269724
rect 250713 269723 250779 269724
rect 416037 269723 416103 269724
rect 425237 269723 425303 269724
rect 433333 269723 433399 269724
rect 434345 269788 434411 269789
rect 434345 269784 434406 269788
rect 434345 269728 434350 269784
rect 434345 269724 434406 269728
rect 434470 269786 434476 269788
rect 434470 269726 434502 269786
rect 434470 269724 434476 269726
rect 434345 269723 434411 269724
rect 83089 269652 83155 269653
rect 91277 269652 91343 269653
rect 93577 269652 93643 269653
rect 94497 269652 94563 269653
rect 143533 269652 143599 269653
rect 83089 269648 83126 269652
rect 83190 269650 83196 269652
rect 83089 269592 83094 269648
rect 83089 269588 83126 269592
rect 83190 269590 83246 269650
rect 91277 269648 91286 269652
rect 91350 269650 91356 269652
rect 91277 269592 91282 269648
rect 83190 269588 83196 269590
rect 91277 269588 91286 269592
rect 91350 269590 91434 269650
rect 93577 269648 93598 269652
rect 93662 269650 93668 269652
rect 93577 269592 93582 269648
rect 91350 269588 91356 269590
rect 93577 269588 93598 269592
rect 93662 269590 93734 269650
rect 94497 269648 94550 269652
rect 94614 269650 94620 269652
rect 143504 269650 143510 269652
rect 94497 269592 94502 269648
rect 93662 269588 93668 269590
rect 94497 269588 94550 269592
rect 94614 269590 94654 269650
rect 143442 269590 143510 269650
rect 143574 269648 143599 269652
rect 143594 269592 143599 269648
rect 94614 269588 94620 269590
rect 143504 269588 143510 269590
rect 143574 269588 143599 269592
rect 83089 269587 83155 269588
rect 91277 269587 91343 269588
rect 93577 269587 93643 269588
rect 94497 269587 94563 269588
rect 143533 269587 143599 269588
rect 145925 269652 145991 269653
rect 283465 269652 283531 269653
rect 288249 269652 288315 269653
rect 291009 269652 291075 269653
rect 145925 269648 145958 269652
rect 146022 269650 146028 269652
rect 145925 269592 145930 269648
rect 145925 269588 145958 269592
rect 146022 269590 146082 269650
rect 283465 269648 283518 269652
rect 283582 269650 283588 269652
rect 283465 269592 283470 269648
rect 146022 269588 146028 269590
rect 283465 269588 283518 269592
rect 283582 269590 283622 269650
rect 288249 269648 288278 269652
rect 288342 269650 288348 269652
rect 290992 269650 290998 269652
rect 288249 269592 288254 269648
rect 283582 269588 283588 269590
rect 288249 269588 288278 269592
rect 288342 269590 288406 269650
rect 290918 269590 290998 269650
rect 291062 269648 291075 269652
rect 291070 269592 291075 269648
rect 288342 269588 288348 269590
rect 290992 269588 290998 269590
rect 291062 269588 291075 269592
rect 145925 269587 145991 269588
rect 283465 269587 283531 269588
rect 288249 269587 288315 269588
rect 291009 269587 291075 269588
rect 293401 269652 293467 269653
rect 305913 269652 305979 269653
rect 318425 269652 318491 269653
rect 429745 269652 429811 269653
rect 436001 269652 436067 269653
rect 468477 269652 468543 269653
rect 470961 269652 471027 269653
rect 480897 269652 480963 269653
rect 293401 269648 293446 269652
rect 293510 269650 293516 269652
rect 293401 269592 293406 269648
rect 293401 269588 293446 269592
rect 293510 269590 293558 269650
rect 305913 269648 305958 269652
rect 306022 269650 306028 269652
rect 305913 269592 305918 269648
rect 293510 269588 293516 269590
rect 305913 269588 305958 269592
rect 306022 269590 306070 269650
rect 318425 269648 318470 269652
rect 318534 269650 318540 269652
rect 318425 269592 318430 269648
rect 306022 269588 306028 269590
rect 318425 269588 318470 269592
rect 318534 269590 318582 269650
rect 429745 269648 429782 269652
rect 429846 269650 429852 269652
rect 429745 269592 429750 269648
rect 318534 269588 318540 269590
rect 429745 269588 429782 269592
rect 429846 269590 429902 269650
rect 436001 269648 436038 269652
rect 436102 269650 436108 269652
rect 436001 269592 436006 269648
rect 429846 269588 429852 269590
rect 436001 269588 436038 269592
rect 436102 269590 436158 269650
rect 468477 269648 468542 269652
rect 468477 269592 468482 269648
rect 468538 269592 468542 269648
rect 436102 269588 436108 269590
rect 468477 269588 468542 269592
rect 468606 269650 468612 269652
rect 468606 269590 468634 269650
rect 470961 269648 470990 269652
rect 471054 269650 471060 269652
rect 470961 269592 470966 269648
rect 468606 269588 468612 269590
rect 470961 269588 470990 269592
rect 471054 269590 471118 269650
rect 480897 269648 480918 269652
rect 480982 269650 480988 269652
rect 480897 269592 480902 269648
rect 471054 269588 471060 269590
rect 480897 269588 480918 269592
rect 480982 269590 481054 269650
rect 480982 269588 480988 269590
rect 293401 269587 293467 269588
rect 305913 269587 305979 269588
rect 318425 269587 318491 269588
rect 429745 269587 429811 269588
rect 436001 269587 436067 269588
rect 468477 269587 468543 269588
rect 470961 269587 471027 269588
rect 480897 269587 480963 269588
rect 370313 269378 370379 269381
rect 376886 269378 376892 269380
rect 370313 269376 376892 269378
rect 370313 269320 370318 269376
rect 370374 269320 376892 269376
rect 370313 269318 376892 269320
rect 370313 269315 370379 269318
rect 376886 269316 376892 269318
rect 376956 269378 376962 269380
rect 377990 269378 377996 269380
rect 376956 269318 377996 269378
rect 376956 269316 376962 269318
rect 377990 269316 377996 269318
rect 378060 269316 378066 269380
rect 359590 269180 359596 269244
rect 359660 269242 359666 269244
rect 473486 269242 473492 269244
rect 359660 269182 473492 269242
rect 359660 269180 359666 269182
rect 473486 269180 473492 269182
rect 473556 269180 473562 269244
rect 54385 269106 54451 269109
rect 323301 269108 323367 269109
rect 115790 269106 115796 269108
rect 54385 269104 115796 269106
rect 54385 269048 54390 269104
rect 54446 269048 115796 269104
rect 54385 269046 115796 269048
rect 54385 269043 54451 269046
rect 115790 269044 115796 269046
rect 115860 269044 115866 269108
rect 196750 269044 196756 269108
rect 196820 269106 196826 269108
rect 311014 269106 311020 269108
rect 196820 269046 311020 269106
rect 196820 269044 196826 269046
rect 311014 269044 311020 269046
rect 311084 269044 311090 269108
rect 323301 269104 323348 269108
rect 323412 269106 323418 269108
rect 358537 269106 358603 269109
rect 485998 269106 486004 269108
rect 323301 269048 323306 269104
rect 323301 269044 323348 269048
rect 323412 269046 323458 269106
rect 358537 269104 486004 269106
rect 358537 269048 358542 269104
rect 358598 269048 486004 269104
rect 358537 269046 486004 269048
rect 323412 269044 323418 269046
rect 323301 269043 323367 269044
rect 358537 269043 358603 269046
rect 485998 269044 486004 269046
rect 486068 269044 486074 269108
rect 56961 268970 57027 268973
rect 422845 268972 422911 268973
rect 425973 268972 426039 268973
rect 430941 268972 431007 268973
rect 432229 268972 432295 268973
rect 475837 268972 475903 268973
rect 478413 268972 478479 268973
rect 483381 268972 483447 268973
rect 116894 268970 116900 268972
rect 56961 268968 116900 268970
rect 56961 268912 56966 268968
rect 57022 268912 116900 268968
rect 56961 268910 116900 268912
rect 56961 268907 57027 268910
rect 116894 268908 116900 268910
rect 116964 268908 116970 268972
rect 217358 268908 217364 268972
rect 217428 268970 217434 268972
rect 320950 268970 320956 268972
rect 217428 268910 320956 268970
rect 217428 268908 217434 268910
rect 320950 268908 320956 268910
rect 321020 268908 321026 268972
rect 359406 268908 359412 268972
rect 359476 268970 359482 268972
rect 359476 268910 422310 268970
rect 359476 268908 359482 268910
rect 76005 268836 76071 268837
rect 77109 268836 77175 268837
rect 90725 268836 90791 268837
rect 95877 268836 95943 268837
rect 96061 268836 96127 268837
rect 98453 268836 98519 268837
rect 99373 268836 99439 268837
rect 100753 268836 100819 268837
rect 76005 268832 76052 268836
rect 76116 268834 76122 268836
rect 76005 268776 76010 268832
rect 76005 268772 76052 268776
rect 76116 268774 76162 268834
rect 77109 268832 77156 268836
rect 77220 268834 77226 268836
rect 77109 268776 77114 268832
rect 76116 268772 76122 268774
rect 77109 268772 77156 268776
rect 77220 268774 77266 268834
rect 90725 268832 90772 268836
rect 90836 268834 90842 268836
rect 95877 268834 95924 268836
rect 90725 268776 90730 268832
rect 77220 268772 77226 268774
rect 90725 268772 90772 268776
rect 90836 268774 90882 268834
rect 95832 268832 95924 268834
rect 95832 268776 95882 268832
rect 95832 268774 95924 268776
rect 90836 268772 90842 268774
rect 95877 268772 95924 268774
rect 95988 268772 95994 268836
rect 96061 268832 96108 268836
rect 96172 268834 96178 268836
rect 96061 268776 96066 268832
rect 96061 268772 96108 268776
rect 96172 268774 96218 268834
rect 98453 268832 98500 268836
rect 98564 268834 98570 268836
rect 98453 268776 98458 268832
rect 96172 268772 96178 268774
rect 98453 268772 98500 268776
rect 98564 268774 98610 268834
rect 99373 268832 99420 268836
rect 99484 268834 99490 268836
rect 100702 268834 100708 268836
rect 99373 268776 99378 268832
rect 98564 268772 98570 268774
rect 99373 268772 99420 268776
rect 99484 268774 99530 268834
rect 100662 268774 100708 268834
rect 100772 268832 100819 268836
rect 100814 268776 100819 268832
rect 99484 268772 99490 268774
rect 100702 268772 100708 268774
rect 100772 268772 100819 268776
rect 76005 268771 76071 268772
rect 77109 268771 77175 268772
rect 90725 268771 90791 268772
rect 95877 268771 95943 268772
rect 96061 268771 96127 268772
rect 98453 268771 98519 268772
rect 99373 268771 99439 268772
rect 100753 268771 100819 268772
rect 106365 268836 106431 268837
rect 106365 268832 106412 268836
rect 106476 268834 106482 268836
rect 216949 268834 217015 268837
rect 243077 268836 243143 268837
rect 217542 268834 217548 268836
rect 106365 268776 106370 268832
rect 106365 268772 106412 268776
rect 106476 268774 106522 268834
rect 216949 268832 217548 268834
rect 216949 268776 216954 268832
rect 217010 268776 217548 268832
rect 216949 268774 217548 268776
rect 106476 268772 106482 268774
rect 106365 268771 106431 268772
rect 216949 268771 217015 268774
rect 217542 268772 217548 268774
rect 217612 268772 217618 268836
rect 243077 268832 243124 268836
rect 243188 268834 243194 268836
rect 243077 268776 243082 268832
rect 243077 268772 243124 268776
rect 243188 268774 243234 268834
rect 243188 268772 243194 268774
rect 257838 268772 257844 268836
rect 257908 268834 257914 268836
rect 258073 268834 258139 268837
rect 257908 268832 258139 268834
rect 257908 268776 258078 268832
rect 258134 268776 258139 268832
rect 257908 268774 258139 268776
rect 257908 268772 257914 268774
rect 243077 268771 243143 268772
rect 258073 268771 258139 268774
rect 261661 268836 261727 268837
rect 295885 268836 295951 268837
rect 298461 268836 298527 268837
rect 300853 268836 300919 268837
rect 303429 268836 303495 268837
rect 416957 268836 417023 268837
rect 421005 268836 421071 268837
rect 261661 268832 261708 268836
rect 261772 268834 261778 268836
rect 261661 268776 261666 268832
rect 261661 268772 261708 268776
rect 261772 268774 261818 268834
rect 295885 268832 295932 268836
rect 295996 268834 296002 268836
rect 295885 268776 295890 268832
rect 261772 268772 261778 268774
rect 295885 268772 295932 268776
rect 295996 268774 296042 268834
rect 298461 268832 298508 268836
rect 298572 268834 298578 268836
rect 298461 268776 298466 268832
rect 295996 268772 296002 268774
rect 298461 268772 298508 268776
rect 298572 268774 298618 268834
rect 300853 268832 300900 268836
rect 300964 268834 300970 268836
rect 300853 268776 300858 268832
rect 298572 268772 298578 268774
rect 300853 268772 300900 268776
rect 300964 268774 301010 268834
rect 303429 268832 303476 268836
rect 303540 268834 303546 268836
rect 303429 268776 303434 268832
rect 300964 268772 300970 268774
rect 303429 268772 303476 268776
rect 303540 268774 303586 268834
rect 303540 268772 303546 268774
rect 377990 268772 377996 268836
rect 378060 268834 378066 268836
rect 378060 268774 412650 268834
rect 378060 268772 378066 268774
rect 261661 268771 261727 268772
rect 295885 268771 295951 268772
rect 298461 268771 298527 268772
rect 300853 268771 300919 268772
rect 303429 268771 303495 268772
rect 412590 268698 412650 268774
rect 416957 268832 417004 268836
rect 417068 268834 417074 268836
rect 416957 268776 416962 268832
rect 416957 268772 417004 268776
rect 417068 268774 417114 268834
rect 421005 268832 421052 268836
rect 421116 268834 421122 268836
rect 422250 268834 422310 268910
rect 422845 268968 422892 268972
rect 422956 268970 422962 268972
rect 422845 268912 422850 268968
rect 422845 268908 422892 268912
rect 422956 268910 423002 268970
rect 425973 268968 426020 268972
rect 426084 268970 426090 268972
rect 425973 268912 425978 268968
rect 422956 268908 422962 268910
rect 425973 268908 426020 268912
rect 426084 268910 426130 268970
rect 430941 268968 430988 268972
rect 431052 268970 431058 268972
rect 430941 268912 430946 268968
rect 426084 268908 426090 268910
rect 430941 268908 430988 268912
rect 431052 268910 431098 268970
rect 432229 268968 432276 268972
rect 432340 268970 432346 268972
rect 432229 268912 432234 268968
rect 431052 268908 431058 268910
rect 432229 268908 432276 268912
rect 432340 268910 432386 268970
rect 475837 268968 475884 268972
rect 475948 268970 475954 268972
rect 475837 268912 475842 268968
rect 432340 268908 432346 268910
rect 475837 268908 475884 268912
rect 475948 268910 475994 268970
rect 478413 268968 478460 268972
rect 478524 268970 478530 268972
rect 478413 268912 478418 268968
rect 475948 268908 475954 268910
rect 478413 268908 478460 268912
rect 478524 268910 478570 268970
rect 483381 268968 483428 268972
rect 483492 268970 483498 268972
rect 483381 268912 483386 268968
rect 478524 268908 478530 268910
rect 483381 268908 483428 268912
rect 483492 268910 483538 268970
rect 483492 268908 483498 268910
rect 422845 268907 422911 268908
rect 425973 268907 426039 268908
rect 430941 268907 431007 268908
rect 432229 268907 432295 268908
rect 475837 268907 475903 268908
rect 478413 268907 478479 268908
rect 483381 268907 483447 268908
rect 423438 268834 423444 268836
rect 421005 268776 421010 268832
rect 417068 268772 417074 268774
rect 421005 268772 421052 268776
rect 421116 268774 421162 268834
rect 422250 268774 423444 268834
rect 421116 268772 421122 268774
rect 423438 268772 423444 268774
rect 423508 268772 423514 268836
rect 416957 268771 417023 268772
rect 421005 268771 421071 268772
rect 423990 268698 423996 268700
rect 412590 268638 423996 268698
rect 423990 268636 423996 268638
rect 424060 268636 424066 268700
rect 53741 268562 53807 268565
rect 101806 268562 101812 268564
rect 53741 268560 101812 268562
rect 53741 268504 53746 268560
rect 53802 268504 101812 268560
rect 53741 268502 101812 268504
rect 53741 268499 53807 268502
rect 101806 268500 101812 268502
rect 101876 268500 101882 268564
rect 50981 268426 51047 268429
rect 103830 268426 103836 268428
rect 50981 268424 103836 268426
rect 50981 268368 50986 268424
rect 51042 268368 103836 268424
rect 50981 268366 103836 268368
rect 50981 268363 51047 268366
rect 103830 268364 103836 268366
rect 103900 268364 103906 268428
rect 85389 268156 85455 268157
rect 92381 268156 92447 268157
rect 85389 268152 85436 268156
rect 85500 268154 85506 268156
rect 85389 268096 85394 268152
rect 85389 268092 85436 268096
rect 85500 268094 85546 268154
rect 92381 268152 92428 268156
rect 92492 268154 92498 268156
rect 92381 268096 92386 268152
rect 85500 268092 85506 268094
rect 92381 268092 92428 268096
rect 92492 268094 92538 268154
rect 92492 268092 92498 268094
rect 103278 268092 103284 268156
rect 103348 268154 103354 268156
rect 103513 268154 103579 268157
rect 103348 268152 103579 268154
rect 103348 268096 103518 268152
rect 103574 268096 103579 268152
rect 103348 268094 103579 268096
rect 103348 268092 103354 268094
rect 85389 268091 85455 268092
rect 92381 268091 92447 268092
rect 103513 268091 103579 268094
rect 113541 268156 113607 268157
rect 128353 268156 128419 268157
rect 113541 268152 113588 268156
rect 113652 268154 113658 268156
rect 128302 268154 128308 268156
rect 113541 268096 113546 268152
rect 113541 268092 113588 268096
rect 113652 268094 113698 268154
rect 128262 268094 128308 268154
rect 128372 268152 128419 268156
rect 128414 268096 128419 268152
rect 113652 268092 113658 268094
rect 128302 268092 128308 268094
rect 128372 268092 128419 268096
rect 113541 268091 113607 268092
rect 128353 268091 128419 268092
rect 265157 268156 265223 268157
rect 275921 268156 275987 268157
rect 265157 268152 265204 268156
rect 265268 268154 265274 268156
rect 275870 268154 275876 268156
rect 265157 268096 265162 268152
rect 265157 268092 265204 268096
rect 265268 268094 265314 268154
rect 275830 268094 275876 268154
rect 275940 268152 275987 268156
rect 275982 268096 275987 268152
rect 265268 268092 265274 268094
rect 275870 268092 275876 268094
rect 275940 268092 275987 268096
rect 265157 268091 265223 268092
rect 275921 268091 275987 268092
rect 398189 268156 398255 268157
rect 401685 268156 401751 268157
rect 455781 268156 455847 268157
rect 398189 268152 398236 268156
rect 398300 268154 398306 268156
rect 398189 268096 398194 268152
rect 398189 268092 398236 268096
rect 398300 268094 398346 268154
rect 401685 268152 401732 268156
rect 401796 268154 401802 268156
rect 401685 268096 401690 268152
rect 398300 268092 398306 268094
rect 401685 268092 401732 268096
rect 401796 268094 401842 268154
rect 455781 268152 455828 268156
rect 455892 268154 455898 268156
rect 455781 268096 455786 268152
rect 401796 268092 401802 268094
rect 455781 268092 455828 268096
rect 455892 268094 455938 268154
rect 455892 268092 455898 268094
rect 463550 268092 463556 268156
rect 463620 268092 463626 268156
rect 398189 268091 398255 268092
rect 401685 268091 401751 268092
rect 455781 268091 455847 268092
rect 217542 267956 217548 268020
rect 217612 268018 217618 268020
rect 217961 268018 218027 268021
rect 217612 268016 218027 268018
rect 217612 267960 217966 268016
rect 218022 267960 218027 268016
rect 217612 267958 218027 267960
rect 217612 267956 217618 267958
rect 217961 267955 218027 267958
rect 216990 267820 216996 267884
rect 217060 267882 217066 267884
rect 220813 267882 220879 267885
rect 217060 267880 220879 267882
rect 217060 267824 220818 267880
rect 220874 267824 220879 267880
rect 217060 267822 220879 267824
rect 217060 267820 217066 267822
rect 220813 267819 220879 267822
rect 83958 267684 83964 267748
rect 84028 267746 84034 267748
rect 84193 267746 84259 267749
rect 96981 267748 97047 267749
rect 96981 267746 97028 267748
rect 84028 267744 84259 267746
rect 84028 267688 84198 267744
rect 84254 267688 84259 267744
rect 84028 267686 84259 267688
rect 96936 267744 97028 267746
rect 96936 267688 96986 267744
rect 96936 267686 97028 267688
rect 84028 267684 84034 267686
rect 84193 267683 84259 267686
rect 96981 267684 97028 267686
rect 97092 267684 97098 267748
rect 97993 267746 98059 267749
rect 102685 267748 102751 267749
rect 111241 267748 111307 267749
rect 112345 267748 112411 267749
rect 98126 267746 98132 267748
rect 97993 267744 98132 267746
rect 97993 267688 97998 267744
rect 98054 267688 98132 267744
rect 97993 267686 98132 267688
rect 96981 267683 97047 267684
rect 97993 267683 98059 267686
rect 98126 267684 98132 267686
rect 98196 267684 98202 267748
rect 102685 267746 102732 267748
rect 102640 267744 102732 267746
rect 102640 267688 102690 267744
rect 102640 267686 102732 267688
rect 102685 267684 102732 267686
rect 102796 267684 102802 267748
rect 111190 267746 111196 267748
rect 111150 267686 111196 267746
rect 111260 267744 111307 267748
rect 112294 267746 112300 267748
rect 111302 267688 111307 267744
rect 111190 267684 111196 267686
rect 111260 267684 111307 267688
rect 112254 267686 112300 267746
rect 112364 267744 112411 267748
rect 119061 267748 119127 267749
rect 119061 267746 119108 267748
rect 112406 267688 112411 267744
rect 112294 267684 112300 267686
rect 112364 267684 112411 267688
rect 119016 267744 119108 267746
rect 119016 267688 119066 267744
rect 119016 267686 119108 267688
rect 102685 267683 102751 267684
rect 111241 267683 111307 267684
rect 112345 267683 112411 267684
rect 119061 267684 119108 267686
rect 119172 267684 119178 267748
rect 120073 267746 120139 267749
rect 120758 267746 120764 267748
rect 120073 267744 120764 267746
rect 120073 267688 120078 267744
rect 120134 267688 120764 267744
rect 120073 267686 120764 267688
rect 119061 267683 119127 267684
rect 120073 267683 120139 267686
rect 120758 267684 120764 267686
rect 120828 267684 120834 267748
rect 125593 267746 125659 267749
rect 150985 267748 151051 267749
rect 158529 267748 158595 267749
rect 163497 267748 163563 267749
rect 125910 267746 125916 267748
rect 125593 267744 125916 267746
rect 125593 267688 125598 267744
rect 125654 267688 125916 267744
rect 125593 267686 125916 267688
rect 125593 267683 125659 267686
rect 125910 267684 125916 267686
rect 125980 267684 125986 267748
rect 150934 267746 150940 267748
rect 150894 267686 150940 267746
rect 151004 267744 151051 267748
rect 158478 267746 158484 267748
rect 151046 267688 151051 267744
rect 150934 267684 150940 267686
rect 151004 267684 151051 267688
rect 158438 267686 158484 267746
rect 158548 267744 158595 267748
rect 163446 267746 163452 267748
rect 158590 267688 158595 267744
rect 158478 267684 158484 267686
rect 158548 267684 158595 267688
rect 163406 267686 163452 267746
rect 163516 267744 163563 267748
rect 163558 267688 163563 267744
rect 163446 267684 163452 267686
rect 163516 267684 163563 267688
rect 150985 267683 151051 267684
rect 158529 267683 158595 267684
rect 163497 267683 163563 267684
rect 255313 267746 255379 267749
rect 255814 267746 255820 267748
rect 255313 267744 255820 267746
rect 255313 267688 255318 267744
rect 255374 267688 255820 267744
rect 255313 267686 255820 267688
rect 255313 267683 255379 267686
rect 255814 267684 255820 267686
rect 255884 267684 255890 267748
rect 258257 267746 258323 267749
rect 258390 267746 258396 267748
rect 258257 267744 258396 267746
rect 258257 267688 258262 267744
rect 258318 267688 258396 267744
rect 258257 267686 258396 267688
rect 258257 267683 258323 267686
rect 258390 267684 258396 267686
rect 258460 267684 258466 267748
rect 260833 267746 260899 267749
rect 263593 267748 263659 267749
rect 260966 267746 260972 267748
rect 260833 267744 260972 267746
rect 260833 267688 260838 267744
rect 260894 267688 260972 267744
rect 260833 267686 260972 267688
rect 260833 267683 260899 267686
rect 260966 267684 260972 267686
rect 261036 267684 261042 267748
rect 263542 267684 263548 267748
rect 263612 267746 263659 267748
rect 264973 267746 265039 267749
rect 265934 267746 265940 267748
rect 263612 267744 263704 267746
rect 263654 267688 263704 267744
rect 263612 267686 263704 267688
rect 264973 267744 265940 267746
rect 264973 267688 264978 267744
rect 265034 267688 265940 267744
rect 264973 267686 265940 267688
rect 263612 267684 263659 267686
rect 263593 267683 263659 267684
rect 264973 267683 265039 267686
rect 265934 267684 265940 267686
rect 266004 267684 266010 267748
rect 267825 267746 267891 267749
rect 268326 267746 268332 267748
rect 267825 267744 268332 267746
rect 267825 267688 267830 267744
rect 267886 267688 268332 267744
rect 267825 267686 268332 267688
rect 267825 267683 267891 267686
rect 268326 267684 268332 267686
rect 268396 267684 268402 267748
rect 270493 267746 270559 267749
rect 270902 267746 270908 267748
rect 270493 267744 270908 267746
rect 270493 267688 270498 267744
rect 270554 267688 270908 267744
rect 270493 267686 270908 267688
rect 270493 267683 270559 267686
rect 270902 267684 270908 267686
rect 270972 267684 270978 267748
rect 273253 267746 273319 267749
rect 273478 267746 273484 267748
rect 273253 267744 273484 267746
rect 273253 267688 273258 267744
rect 273314 267688 273484 267744
rect 273253 267686 273484 267688
rect 273253 267683 273319 267686
rect 273478 267684 273484 267686
rect 273548 267684 273554 267748
rect 276013 267746 276079 267749
rect 277025 267748 277091 267749
rect 278129 267748 278195 267749
rect 276238 267746 276244 267748
rect 276013 267744 276244 267746
rect 276013 267688 276018 267744
rect 276074 267688 276244 267744
rect 276013 267686 276244 267688
rect 276013 267683 276079 267686
rect 276238 267684 276244 267686
rect 276308 267684 276314 267748
rect 276974 267746 276980 267748
rect 276934 267686 276980 267746
rect 277044 267744 277091 267748
rect 278078 267746 278084 267748
rect 277086 267688 277091 267744
rect 276974 267684 276980 267686
rect 277044 267684 277091 267688
rect 278038 267686 278084 267746
rect 278148 267744 278195 267748
rect 278190 267688 278195 267744
rect 278078 267684 278084 267686
rect 278148 267684 278195 267688
rect 277025 267683 277091 267684
rect 278129 267683 278195 267684
rect 280153 267746 280219 267749
rect 402973 267748 403039 267749
rect 414381 267748 414447 267749
rect 280838 267746 280844 267748
rect 280153 267744 280844 267746
rect 280153 267688 280158 267744
rect 280214 267688 280844 267744
rect 280153 267686 280844 267688
rect 280153 267683 280219 267686
rect 280838 267684 280844 267686
rect 280908 267684 280914 267748
rect 402973 267744 403020 267748
rect 403084 267746 403090 267748
rect 414381 267746 414428 267748
rect 402973 267688 402978 267744
rect 402973 267684 403020 267688
rect 403084 267686 403130 267746
rect 414336 267744 414428 267746
rect 414336 267688 414386 267744
rect 414336 267686 414428 267688
rect 403084 267684 403090 267686
rect 414381 267684 414428 267686
rect 414492 267684 414498 267748
rect 415393 267746 415459 267749
rect 428641 267748 428707 267749
rect 415526 267746 415532 267748
rect 415393 267744 415532 267746
rect 415393 267688 415398 267744
rect 415454 267688 415532 267744
rect 415393 267686 415532 267688
rect 402973 267683 403039 267684
rect 414381 267683 414447 267684
rect 415393 267683 415459 267686
rect 415526 267684 415532 267686
rect 415596 267684 415602 267748
rect 428590 267684 428596 267748
rect 428660 267746 428707 267748
rect 434713 267746 434779 267749
rect 435582 267746 435588 267748
rect 428660 267744 428752 267746
rect 428702 267688 428752 267744
rect 428660 267686 428752 267688
rect 434713 267744 435588 267746
rect 434713 267688 434718 267744
rect 434774 267688 435588 267744
rect 434713 267686 435588 267688
rect 428660 267684 428707 267686
rect 428641 267683 428707 267684
rect 434713 267683 434779 267686
rect 435582 267684 435588 267686
rect 435652 267684 435658 267748
rect 449893 267746 449959 267749
rect 451038 267746 451044 267748
rect 449893 267744 451044 267746
rect 449893 267688 449898 267744
rect 449954 267688 451044 267744
rect 449893 267686 451044 267688
rect 449893 267683 449959 267686
rect 451038 267684 451044 267686
rect 451108 267684 451114 267748
rect 452653 267746 452719 267749
rect 453430 267746 453436 267748
rect 452653 267744 453436 267746
rect 452653 267688 452658 267744
rect 452714 267688 453436 267744
rect 452653 267686 453436 267688
rect 452653 267683 452719 267686
rect 453430 267684 453436 267686
rect 453500 267684 453506 267748
rect 458173 267746 458239 267749
rect 460933 267748 460999 267749
rect 458398 267746 458404 267748
rect 458173 267744 458404 267746
rect 458173 267688 458178 267744
rect 458234 267688 458404 267744
rect 458173 267686 458404 267688
rect 458173 267683 458239 267686
rect 458398 267684 458404 267686
rect 458468 267684 458474 267748
rect 460933 267744 460980 267748
rect 461044 267746 461050 267748
rect 460933 267688 460938 267744
rect 460933 267684 460980 267688
rect 461044 267686 461090 267746
rect 461044 267684 461050 267686
rect 460933 267683 460999 267684
rect 57830 267548 57836 267612
rect 57900 267610 57906 267612
rect 123518 267610 123524 267612
rect 57900 267550 123524 267610
rect 57900 267548 57906 267550
rect 123518 267548 123524 267550
rect 123588 267548 123594 267612
rect 129733 267610 129799 267613
rect 155953 267612 156019 267613
rect 160921 267612 160987 267613
rect 130878 267610 130884 267612
rect 129733 267608 130884 267610
rect 129733 267552 129738 267608
rect 129794 267552 130884 267608
rect 129733 267550 130884 267552
rect 129733 267547 129799 267550
rect 130878 267548 130884 267550
rect 130948 267548 130954 267612
rect 155902 267610 155908 267612
rect 155862 267550 155908 267610
rect 155972 267608 156019 267612
rect 160870 267610 160876 267612
rect 156014 267552 156019 267608
rect 155902 267548 155908 267550
rect 155972 267548 156019 267552
rect 160830 267550 160876 267610
rect 160940 267608 160987 267612
rect 198774 267610 198780 267612
rect 160982 267552 160987 267608
rect 160870 267548 160876 267550
rect 160940 267548 160987 267552
rect 155953 267547 156019 267548
rect 160921 267547 160987 267548
rect 161430 267550 198780 267610
rect 46289 267474 46355 267477
rect 115933 267476 115999 267477
rect 80462 267474 80468 267476
rect 46289 267472 80468 267474
rect 46289 267416 46294 267472
rect 46350 267416 80468 267472
rect 46289 267414 80468 267416
rect 46289 267411 46355 267414
rect 80462 267412 80468 267414
rect 80532 267412 80538 267476
rect 115933 267474 115980 267476
rect 115888 267472 115980 267474
rect 115888 267416 115938 267472
rect 115888 267414 115980 267416
rect 115933 267412 115980 267414
rect 116044 267412 116050 267476
rect 117313 267474 117379 267477
rect 118366 267474 118372 267476
rect 117313 267472 118372 267474
rect 117313 267416 117318 267472
rect 117374 267416 118372 267472
rect 117313 267414 118372 267416
rect 115933 267411 115999 267412
rect 117313 267411 117379 267414
rect 118366 267412 118372 267414
rect 118436 267412 118442 267476
rect 154062 267412 154068 267476
rect 154132 267474 154138 267476
rect 161430 267474 161490 267550
rect 198774 267548 198780 267550
rect 198844 267548 198850 267612
rect 203701 267610 203767 267613
rect 315982 267610 315988 267612
rect 203701 267608 315988 267610
rect 203701 267552 203706 267608
rect 203762 267552 315988 267608
rect 203701 267550 315988 267552
rect 203701 267547 203767 267550
rect 315982 267548 315988 267550
rect 316052 267548 316058 267612
rect 378961 267610 379027 267613
rect 463558 267610 463618 268092
rect 378961 267608 463618 267610
rect 378961 267552 378966 267608
rect 379022 267552 463618 267608
rect 378961 267550 463618 267552
rect 378961 267547 379027 267550
rect 154132 267414 161490 267474
rect 212073 267474 212139 267477
rect 313406 267474 313412 267476
rect 212073 267472 313412 267474
rect 212073 267416 212078 267472
rect 212134 267416 313412 267472
rect 212073 267414 313412 267416
rect 154132 267412 154138 267414
rect 212073 267411 212139 267414
rect 313406 267412 313412 267414
rect 313476 267412 313482 267476
rect 343214 267412 343220 267476
rect 343284 267474 343290 267476
rect 343449 267474 343515 267477
rect 343284 267472 343515 267474
rect 343284 267416 343454 267472
rect 343510 267416 343515 267472
rect 343284 267414 343515 267416
rect 343284 267412 343290 267414
rect 343449 267411 343515 267414
rect 379462 267412 379468 267476
rect 379532 267474 379538 267476
rect 428222 267474 428228 267476
rect 379532 267414 428228 267474
rect 379532 267412 379538 267414
rect 428222 267412 428228 267414
rect 428292 267412 428298 267476
rect 442993 267474 443059 267477
rect 503161 267476 503227 267477
rect 503529 267476 503595 267477
rect 443494 267474 443500 267476
rect 442993 267472 443500 267474
rect 442993 267416 442998 267472
rect 443054 267416 443500 267472
rect 442993 267414 443500 267416
rect 442993 267411 443059 267414
rect 443494 267412 443500 267414
rect 443564 267412 443570 267476
rect 503110 267474 503116 267476
rect 503070 267414 503116 267474
rect 503180 267472 503227 267476
rect 503478 267474 503484 267476
rect 503222 267416 503227 267472
rect 503110 267412 503116 267414
rect 503180 267412 503227 267416
rect 503438 267414 503484 267474
rect 503548 267472 503595 267476
rect 503590 267416 503595 267472
rect 503478 267412 503484 267414
rect 503548 267412 503595 267416
rect 503161 267411 503227 267412
rect 503529 267411 503595 267412
rect 48865 267338 48931 267341
rect 81934 267338 81940 267340
rect 48865 267336 81940 267338
rect -960 267052 480 267292
rect 48865 267280 48870 267336
rect 48926 267280 81940 267336
rect 48865 267278 81940 267280
rect 48865 267275 48931 267278
rect 81934 267276 81940 267278
rect 82004 267276 82010 267340
rect 107653 267338 107719 267341
rect 108246 267338 108252 267340
rect 107653 267336 108252 267338
rect 107653 267280 107658 267336
rect 107714 267280 108252 267336
rect 107653 267278 108252 267280
rect 107653 267275 107719 267278
rect 108246 267276 108252 267278
rect 108316 267276 108322 267340
rect 183134 267276 183140 267340
rect 183204 267338 183210 267340
rect 183277 267338 183343 267341
rect 183204 267336 183343 267338
rect 183204 267280 183282 267336
rect 183338 267280 183343 267336
rect 183204 267278 183343 267280
rect 183204 267276 183210 267278
rect 183277 267275 183343 267278
rect 213269 267338 213335 267341
rect 308622 267338 308628 267340
rect 213269 267336 308628 267338
rect 213269 267280 213274 267336
rect 213330 267280 308628 267336
rect 213269 267278 308628 267280
rect 213269 267275 213335 267278
rect 308622 267276 308628 267278
rect 308692 267276 308698 267340
rect 377254 267276 377260 267340
rect 377324 267338 377330 267340
rect 408166 267338 408172 267340
rect 377324 267278 408172 267338
rect 377324 267276 377330 267278
rect 408166 267276 408172 267278
rect 408236 267276 408242 267340
rect 439262 267276 439268 267340
rect 439332 267338 439338 267340
rect 440049 267338 440115 267341
rect 439332 267336 440115 267338
rect 439332 267280 440054 267336
rect 440110 267280 440115 267336
rect 439332 267278 440115 267280
rect 439332 267276 439338 267278
rect 440049 267275 440115 267278
rect 440233 267338 440299 267341
rect 440918 267338 440924 267340
rect 440233 267336 440924 267338
rect 440233 267280 440238 267336
rect 440294 267280 440924 267336
rect 440233 267278 440924 267280
rect 440233 267275 440299 267278
rect 440918 267276 440924 267278
rect 440988 267276 440994 267340
rect 447133 267338 447199 267341
rect 448278 267338 448284 267340
rect 447133 267336 448284 267338
rect 447133 267280 447138 267336
rect 447194 267280 448284 267336
rect 447133 267278 448284 267280
rect 447133 267275 447199 267278
rect 448278 267276 448284 267278
rect 448348 267276 448354 267340
rect 104893 267202 104959 267205
rect 105854 267202 105860 267204
rect 104893 267200 105860 267202
rect 104893 267144 104898 267200
rect 104954 267144 105860 267200
rect 104893 267142 105860 267144
rect 104893 267139 104959 267142
rect 105854 267140 105860 267142
rect 105924 267140 105930 267204
rect 217174 267140 217180 267204
rect 217244 267202 217250 267204
rect 278446 267202 278452 267204
rect 217244 267142 278452 267202
rect 217244 267140 217250 267142
rect 278446 267140 278452 267142
rect 278516 267140 278522 267204
rect 278998 267140 279004 267204
rect 279068 267202 279074 267204
rect 279141 267202 279207 267205
rect 279068 267200 279207 267202
rect 279068 267144 279146 267200
rect 279202 267144 279207 267200
rect 279068 267142 279207 267144
rect 279068 267140 279074 267142
rect 279141 267139 279207 267142
rect 376569 267202 376635 267205
rect 397126 267202 397132 267204
rect 376569 267200 397132 267202
rect 376569 267144 376574 267200
rect 376630 267144 397132 267200
rect 376569 267142 397132 267144
rect 376569 267139 376635 267142
rect 397126 267140 397132 267142
rect 397196 267140 397202 267204
rect 418153 267202 418219 267205
rect 418470 267202 418476 267204
rect 418153 267200 418476 267202
rect 418153 267144 418158 267200
rect 418214 267144 418476 267200
rect 418153 267142 418476 267144
rect 418153 267139 418219 267142
rect 418470 267140 418476 267142
rect 418540 267140 418546 267204
rect 437473 267202 437539 267205
rect 438526 267202 438532 267204
rect 437473 267200 438532 267202
rect 437473 267144 437478 267200
rect 437534 267144 438532 267200
rect 437473 267142 438532 267144
rect 437473 267139 437539 267142
rect 438526 267140 438532 267142
rect 438596 267140 438602 267204
rect 445753 267202 445819 267205
rect 445886 267202 445892 267204
rect 445753 267200 445892 267202
rect 445753 267144 445758 267200
rect 445814 267144 445892 267200
rect 445753 267142 445892 267144
rect 445753 267139 445819 267142
rect 445886 267140 445892 267142
rect 445956 267140 445962 267204
rect 52913 267066 52979 267069
rect 66253 267066 66319 267069
rect 52913 267064 66319 267066
rect 52913 267008 52918 267064
rect 52974 267008 66258 267064
rect 66314 267008 66319 267064
rect 52913 267006 66319 267008
rect 52913 267003 52979 267006
rect 66253 267003 66319 267006
rect 77293 267066 77359 267069
rect 78254 267066 78260 267068
rect 77293 267064 78260 267066
rect 77293 267008 77298 267064
rect 77354 267008 78260 267064
rect 77293 267006 78260 267008
rect 77293 267003 77359 267006
rect 78254 267004 78260 267006
rect 78324 267004 78330 267068
rect 78673 267066 78739 267069
rect 88333 267068 88399 267069
rect 79542 267066 79548 267068
rect 78673 267064 79548 267066
rect 78673 267008 78678 267064
rect 78734 267008 79548 267064
rect 78673 267006 79548 267008
rect 78673 267003 78739 267006
rect 79542 267004 79548 267006
rect 79612 267004 79618 267068
rect 88333 267066 88380 267068
rect 88288 267064 88380 267066
rect 88288 267008 88338 267064
rect 88288 267006 88380 267008
rect 88333 267004 88380 267006
rect 88444 267004 88450 267068
rect 100753 267066 100819 267069
rect 101070 267066 101076 267068
rect 100753 267064 101076 267066
rect 100753 267008 100758 267064
rect 100814 267008 101076 267064
rect 100753 267006 101076 267008
rect 88333 267003 88399 267004
rect 100753 267003 100819 267006
rect 101070 267004 101076 267006
rect 101140 267004 101146 267068
rect 109534 267004 109540 267068
rect 109604 267066 109610 267068
rect 109953 267066 110019 267069
rect 109604 267064 110019 267066
rect 109604 267008 109958 267064
rect 110014 267008 110019 267064
rect 109604 267006 110019 267008
rect 109604 267004 109610 267006
rect 109953 267003 110019 267006
rect 183461 267068 183527 267069
rect 183461 267064 183508 267068
rect 183572 267066 183578 267068
rect 216305 267066 216371 267069
rect 236494 267066 236500 267068
rect 183461 267008 183466 267064
rect 183461 267004 183508 267008
rect 183572 267006 183618 267066
rect 216305 267064 236500 267066
rect 216305 267008 216310 267064
rect 216366 267008 236500 267064
rect 216305 267006 236500 267008
rect 183572 267004 183578 267006
rect 183461 267003 183527 267004
rect 216305 267003 216371 267006
rect 236494 267004 236500 267006
rect 236564 267004 236570 267068
rect 255313 267066 255379 267069
rect 273253 267068 273319 267069
rect 343449 267068 343515 267069
rect 256182 267066 256188 267068
rect 255313 267064 256188 267066
rect 255313 267008 255318 267064
rect 255374 267008 256188 267064
rect 255313 267006 256188 267008
rect 255313 267003 255379 267006
rect 256182 267004 256188 267006
rect 256252 267004 256258 267068
rect 273253 267066 273300 267068
rect 273208 267064 273300 267066
rect 273208 267008 273258 267064
rect 273208 267006 273300 267008
rect 273253 267004 273300 267006
rect 273364 267004 273370 267068
rect 343398 267066 343404 267068
rect 343358 267006 343404 267066
rect 343468 267064 343515 267068
rect 343510 267008 343515 267064
rect 343398 267004 343404 267006
rect 343468 267004 343515 267008
rect 273253 267003 273319 267004
rect 343449 267003 343515 267004
rect 409873 267066 409939 267069
rect 410742 267066 410748 267068
rect 409873 267064 410748 267066
rect 409873 267008 409878 267064
rect 409934 267008 410748 267064
rect 409873 267006 410748 267008
rect 409873 267003 409939 267006
rect 410742 267004 410748 267006
rect 410812 267004 410818 267068
rect 412909 267066 412975 267069
rect 413686 267066 413692 267068
rect 412909 267064 413692 267066
rect 412909 267008 412914 267064
rect 412970 267008 413692 267064
rect 412909 267006 413692 267008
rect 412909 267003 412975 267006
rect 413686 267004 413692 267006
rect 413756 267004 413762 267068
rect 433333 267066 433399 267069
rect 433558 267066 433564 267068
rect 433333 267064 433564 267066
rect 433333 267008 433338 267064
rect 433394 267008 433564 267064
rect 433333 267006 433564 267008
rect 433333 267003 433399 267006
rect 433558 267004 433564 267006
rect 433628 267004 433634 267068
rect 47945 266930 48011 266933
rect 165838 266930 165844 266932
rect 47945 266928 165844 266930
rect 47945 266872 47950 266928
rect 48006 266872 165844 266928
rect 47945 266870 165844 266872
rect 47945 266867 48011 266870
rect 165838 266868 165844 266870
rect 165908 266868 165914 266932
rect 218421 266930 218487 266933
rect 219249 266930 219315 266933
rect 237046 266930 237052 266932
rect 218421 266928 237052 266930
rect 218421 266872 218426 266928
rect 218482 266872 219254 266928
rect 219310 266872 237052 266928
rect 218421 266870 237052 266872
rect 218421 266867 218487 266870
rect 219249 266867 219315 266870
rect 237046 266868 237052 266870
rect 237116 266868 237122 266932
rect 247033 266930 247099 266933
rect 248270 266930 248276 266932
rect 247033 266928 248276 266930
rect 247033 266872 247038 266928
rect 247094 266872 248276 266928
rect 247033 266870 248276 266872
rect 247033 266867 247099 266870
rect 248270 266868 248276 266870
rect 248340 266868 248346 266932
rect 252553 266930 252619 266933
rect 253606 266930 253612 266932
rect 252553 266928 253612 266930
rect 252553 266872 252558 266928
rect 252614 266872 253612 266928
rect 252553 266870 253612 266872
rect 252553 266867 252619 266870
rect 253606 266868 253612 266870
rect 253676 266868 253682 266932
rect 285673 266930 285739 266933
rect 285990 266930 285996 266932
rect 285673 266928 285996 266930
rect 285673 266872 285678 266928
rect 285734 266872 285996 266928
rect 285673 266870 285996 266872
rect 285673 266867 285739 266870
rect 285990 266868 285996 266870
rect 286060 266868 286066 266932
rect 361113 266930 361179 266933
rect 465942 266930 465948 266932
rect 361113 266928 465948 266930
rect 361113 266872 361118 266928
rect 361174 266872 465948 266928
rect 361113 266870 465948 266872
rect 361113 266867 361179 266870
rect 465942 266868 465948 266870
rect 466012 266868 466018 266932
rect 209405 266794 209471 266797
rect 326654 266794 326660 266796
rect 209405 266792 326660 266794
rect 209405 266736 209410 266792
rect 209466 266736 326660 266792
rect 209405 266734 326660 266736
rect 209405 266731 209471 266734
rect 326654 266732 326660 266734
rect 326724 266732 326730 266796
rect 113214 266596 113220 266660
rect 113284 266658 113290 266660
rect 114369 266658 114435 266661
rect 113284 266656 114435 266658
rect 113284 266600 114374 266656
rect 114430 266600 114435 266656
rect 113284 266598 114435 266600
rect 113284 266596 113290 266598
rect 114369 266595 114435 266598
rect 117313 266658 117379 266661
rect 117998 266658 118004 266660
rect 117313 266656 118004 266658
rect 117313 266600 117318 266656
rect 117374 266600 118004 266656
rect 117313 266598 118004 266600
rect 117313 266595 117379 266598
rect 117998 266596 118004 266598
rect 118068 266596 118074 266660
rect 249793 266658 249859 266661
rect 250110 266658 250116 266660
rect 249793 266656 250116 266658
rect 249793 266600 249798 266656
rect 249854 266600 250116 266656
rect 249793 266598 250116 266600
rect 249793 266595 249859 266598
rect 250110 266596 250116 266598
rect 250180 266596 250186 266660
rect 408493 266658 408559 266661
rect 408718 266658 408724 266660
rect 408493 266656 408724 266658
rect 408493 266600 408498 266656
rect 408554 266600 408724 266656
rect 408493 266598 408724 266600
rect 408493 266595 408559 266598
rect 408718 266596 408724 266598
rect 408788 266596 408794 266660
rect 437473 266658 437539 266661
rect 438342 266658 438348 266660
rect 437473 266656 438348 266658
rect 437473 266600 437478 266656
rect 437534 266600 438348 266656
rect 437473 266598 438348 266600
rect 437473 266595 437539 266598
rect 438342 266596 438348 266598
rect 438412 266596 438418 266660
rect 104893 266522 104959 266525
rect 105302 266522 105308 266524
rect 104893 266520 105308 266522
rect 104893 266464 104898 266520
rect 104954 266464 105308 266520
rect 104893 266462 105308 266464
rect 104893 266459 104959 266462
rect 105302 266460 105308 266462
rect 105372 266460 105378 266524
rect 215334 266460 215340 266524
rect 215404 266522 215410 266524
rect 216489 266522 216555 266525
rect 215404 266520 216555 266522
rect 215404 266464 216494 266520
rect 216550 266464 216555 266520
rect 215404 266462 216555 266464
rect 215404 266460 215410 266462
rect 216489 266459 216555 266462
rect 244222 266460 244228 266524
rect 244292 266522 244298 266524
rect 244365 266522 244431 266525
rect 244292 266520 244431 266522
rect 244292 266464 244370 266520
rect 244426 266464 244431 266520
rect 244292 266462 244431 266464
rect 244292 266460 244298 266462
rect 244365 266459 244431 266462
rect 251265 266522 251331 266525
rect 252318 266522 252324 266524
rect 251265 266520 252324 266522
rect 251265 266464 251270 266520
rect 251326 266464 252324 266520
rect 251265 266462 252324 266464
rect 251265 266459 251331 266462
rect 252318 266460 252324 266462
rect 252388 266460 252394 266524
rect 259545 266522 259611 266525
rect 260598 266522 260604 266524
rect 259545 266520 260604 266522
rect 259545 266464 259550 266520
rect 259606 266464 260604 266520
rect 259545 266462 260604 266464
rect 259545 266459 259611 266462
rect 260598 266460 260604 266462
rect 260668 266460 260674 266524
rect 266353 266522 266419 266525
rect 267590 266522 267596 266524
rect 266353 266520 267596 266522
rect 266353 266464 266358 266520
rect 266414 266464 267596 266520
rect 266353 266462 267596 266464
rect 266353 266459 266419 266462
rect 267590 266460 267596 266462
rect 267660 266460 267666 266524
rect 411345 266522 411411 266525
rect 412398 266522 412404 266524
rect 411345 266520 412404 266522
rect 411345 266464 411350 266520
rect 411406 266464 412404 266520
rect 411345 266462 412404 266464
rect 411345 266459 411411 266462
rect 412398 266460 412404 266462
rect 412468 266460 412474 266524
rect 418245 266522 418311 266525
rect 419206 266522 419212 266524
rect 418245 266520 419212 266522
rect 418245 266464 418250 266520
rect 418306 266464 419212 266520
rect 418245 266462 419212 266464
rect 418245 266459 418311 266462
rect 419206 266460 419212 266462
rect 419276 266460 419282 266524
rect 46289 266386 46355 266389
rect 46473 266386 46539 266389
rect 46289 266384 46539 266386
rect 46289 266328 46294 266384
rect 46350 266328 46478 266384
rect 46534 266328 46539 266384
rect 46289 266326 46539 266328
rect 46289 266323 46355 266326
rect 46473 266323 46539 266326
rect 48865 266386 48931 266389
rect 49141 266386 49207 266389
rect 48865 266384 49207 266386
rect 48865 266328 48870 266384
rect 48926 266328 49146 266384
rect 49202 266328 49207 266384
rect 48865 266326 49207 266328
rect 48865 266323 48931 266326
rect 49141 266323 49207 266326
rect 85573 266386 85639 266389
rect 86534 266386 86540 266388
rect 85573 266384 86540 266386
rect 85573 266328 85578 266384
rect 85634 266328 86540 266384
rect 85573 266326 86540 266328
rect 85573 266323 85639 266326
rect 86534 266324 86540 266326
rect 86604 266324 86610 266388
rect 86953 266386 87019 266389
rect 87454 266386 87460 266388
rect 86953 266384 87460 266386
rect 86953 266328 86958 266384
rect 87014 266328 87460 266384
rect 86953 266326 87460 266328
rect 86953 266323 87019 266326
rect 87454 266324 87460 266326
rect 87524 266324 87530 266388
rect 88333 266386 88399 266389
rect 88742 266386 88748 266388
rect 88333 266384 88748 266386
rect 88333 266328 88338 266384
rect 88394 266328 88748 266384
rect 88333 266326 88748 266328
rect 88333 266323 88399 266326
rect 88742 266324 88748 266326
rect 88812 266324 88818 266388
rect 89713 266386 89779 266389
rect 90030 266386 90036 266388
rect 89713 266384 90036 266386
rect 89713 266328 89718 266384
rect 89774 266328 90036 266384
rect 89713 266326 90036 266328
rect 89713 266323 89779 266326
rect 90030 266324 90036 266326
rect 90100 266324 90106 266388
rect 92473 266386 92539 266389
rect 93342 266386 93348 266388
rect 92473 266384 93348 266386
rect 92473 266328 92478 266384
rect 92534 266328 93348 266384
rect 92473 266326 93348 266328
rect 92473 266323 92539 266326
rect 93342 266324 93348 266326
rect 93412 266324 93418 266388
rect 106273 266386 106339 266389
rect 107510 266386 107516 266388
rect 106273 266384 107516 266386
rect 106273 266328 106278 266384
rect 106334 266328 107516 266384
rect 106273 266326 107516 266328
rect 106273 266323 106339 266326
rect 107510 266324 107516 266326
rect 107580 266324 107586 266388
rect 107653 266386 107719 266389
rect 108614 266386 108620 266388
rect 107653 266384 108620 266386
rect 107653 266328 107658 266384
rect 107714 266328 108620 266384
rect 107653 266326 108620 266328
rect 107653 266323 107719 266326
rect 108614 266324 108620 266326
rect 108684 266324 108690 266388
rect 113725 266386 113791 266389
rect 114318 266386 114324 266388
rect 113725 266384 114324 266386
rect 113725 266328 113730 266384
rect 113786 266328 114324 266384
rect 113725 266326 114324 266328
rect 113725 266323 113791 266326
rect 114318 266324 114324 266326
rect 114388 266324 114394 266388
rect 215293 266386 215359 266389
rect 215518 266386 215524 266388
rect 215293 266384 215524 266386
rect 215293 266328 215298 266384
rect 215354 266328 215524 266384
rect 215293 266326 215524 266328
rect 215293 266323 215359 266326
rect 215518 266324 215524 266326
rect 215588 266324 215594 266388
rect 244273 266386 244339 266389
rect 245326 266386 245332 266388
rect 244273 266384 245332 266386
rect 244273 266328 244278 266384
rect 244334 266328 245332 266384
rect 244273 266326 245332 266328
rect 244273 266323 244339 266326
rect 245326 266324 245332 266326
rect 245396 266324 245402 266388
rect 245653 266386 245719 266389
rect 246430 266386 246436 266388
rect 245653 266384 246436 266386
rect 245653 266328 245658 266384
rect 245714 266328 246436 266384
rect 245653 266326 246436 266328
rect 245653 266323 245719 266326
rect 246430 266324 246436 266326
rect 246500 266324 246506 266388
rect 247033 266386 247099 266389
rect 247718 266386 247724 266388
rect 247033 266384 247724 266386
rect 247033 266328 247038 266384
rect 247094 266328 247724 266384
rect 247033 266326 247724 266328
rect 247033 266323 247099 266326
rect 247718 266324 247724 266326
rect 247788 266324 247794 266388
rect 248505 266386 248571 266389
rect 251173 266388 251239 266389
rect 248638 266386 248644 266388
rect 248505 266384 248644 266386
rect 248505 266328 248510 266384
rect 248566 266328 248644 266384
rect 248505 266326 248644 266328
rect 248505 266323 248571 266326
rect 248638 266324 248644 266326
rect 248708 266324 248714 266388
rect 251173 266386 251220 266388
rect 251128 266384 251220 266386
rect 251128 266328 251178 266384
rect 251128 266326 251220 266328
rect 251173 266324 251220 266326
rect 251284 266324 251290 266388
rect 252553 266386 252619 266389
rect 253422 266386 253428 266388
rect 252553 266384 253428 266386
rect 252553 266328 252558 266384
rect 252614 266328 253428 266384
rect 252553 266326 253428 266328
rect 251173 266323 251239 266324
rect 252553 266323 252619 266326
rect 253422 266324 253428 266326
rect 253492 266324 253498 266388
rect 253933 266386 253999 266389
rect 254526 266386 254532 266388
rect 253933 266384 254532 266386
rect 253933 266328 253938 266384
rect 253994 266328 254532 266384
rect 253933 266326 254532 266328
rect 253933 266323 253999 266326
rect 254526 266324 254532 266326
rect 254596 266324 254602 266388
rect 256693 266386 256759 266389
rect 259453 266388 259519 266389
rect 256918 266386 256924 266388
rect 256693 266384 256924 266386
rect 256693 266328 256698 266384
rect 256754 266328 256924 266384
rect 256693 266326 256924 266328
rect 256693 266323 256759 266326
rect 256918 266324 256924 266326
rect 256988 266324 256994 266388
rect 259453 266386 259500 266388
rect 259408 266384 259500 266386
rect 259408 266328 259458 266384
rect 259408 266326 259500 266328
rect 259453 266324 259500 266326
rect 259564 266324 259570 266388
rect 262213 266386 262279 266389
rect 262806 266386 262812 266388
rect 262213 266384 262812 266386
rect 262213 266328 262218 266384
rect 262274 266328 262812 266384
rect 262213 266326 262812 266328
rect 259453 266323 259519 266324
rect 262213 266323 262279 266326
rect 262806 266324 262812 266326
rect 262876 266324 262882 266388
rect 263593 266386 263659 266389
rect 263910 266386 263916 266388
rect 263593 266384 263916 266386
rect 263593 266328 263598 266384
rect 263654 266328 263916 266384
rect 263593 266326 263916 266328
rect 263593 266323 263659 266326
rect 263910 266324 263916 266326
rect 263980 266324 263986 266388
rect 266302 266324 266308 266388
rect 266372 266386 266378 266388
rect 266445 266386 266511 266389
rect 266372 266384 266511 266386
rect 266372 266328 266450 266384
rect 266506 266328 266511 266384
rect 266372 266326 266511 266328
rect 266372 266324 266378 266326
rect 266445 266323 266511 266326
rect 267733 266386 267799 266389
rect 268694 266386 268700 266388
rect 267733 266384 268700 266386
rect 267733 266328 267738 266384
rect 267794 266328 268700 266384
rect 267733 266326 268700 266328
rect 267733 266323 267799 266326
rect 268694 266324 268700 266326
rect 268764 266324 268770 266388
rect 269113 266386 269179 266389
rect 269798 266386 269804 266388
rect 269113 266384 269804 266386
rect 269113 266328 269118 266384
rect 269174 266328 269804 266384
rect 269113 266326 269804 266328
rect 269113 266323 269179 266326
rect 269798 266324 269804 266326
rect 269868 266324 269874 266388
rect 270493 266386 270559 266389
rect 271270 266386 271276 266388
rect 270493 266384 271276 266386
rect 270493 266328 270498 266384
rect 270554 266328 271276 266384
rect 270493 266326 271276 266328
rect 270493 266323 270559 266326
rect 271270 266324 271276 266326
rect 271340 266324 271346 266388
rect 273161 266386 273227 266389
rect 274398 266386 274404 266388
rect 273161 266384 274404 266386
rect 273161 266328 273166 266384
rect 273222 266328 274404 266384
rect 273161 266326 274404 266328
rect 273161 266323 273227 266326
rect 274398 266324 274404 266326
rect 274468 266324 274474 266388
rect 375833 266386 375899 266389
rect 376569 266386 376635 266389
rect 396073 266388 396139 266389
rect 375833 266384 376635 266386
rect 375833 266328 375838 266384
rect 375894 266328 376574 266384
rect 376630 266328 376635 266384
rect 375833 266326 376635 266328
rect 375833 266323 375899 266326
rect 376569 266323 376635 266326
rect 396022 266324 396028 266388
rect 396092 266386 396139 266388
rect 398833 266386 398899 266389
rect 399518 266386 399524 266388
rect 396092 266384 396184 266386
rect 396134 266328 396184 266384
rect 396092 266326 396184 266328
rect 398833 266384 399524 266386
rect 398833 266328 398838 266384
rect 398894 266328 399524 266384
rect 398833 266326 399524 266328
rect 396092 266324 396139 266326
rect 396073 266323 396139 266324
rect 398833 266323 398899 266326
rect 399518 266324 399524 266326
rect 399588 266324 399594 266388
rect 400213 266386 400279 266389
rect 400438 266386 400444 266388
rect 400213 266384 400444 266386
rect 400213 266328 400218 266384
rect 400274 266328 400444 266384
rect 400213 266326 400444 266328
rect 400213 266323 400279 266326
rect 400438 266324 400444 266326
rect 400508 266324 400514 266388
rect 403157 266386 403223 266389
rect 404118 266386 404124 266388
rect 403157 266384 404124 266386
rect 403157 266328 403162 266384
rect 403218 266328 404124 266384
rect 403157 266326 404124 266328
rect 403157 266323 403223 266326
rect 404118 266324 404124 266326
rect 404188 266324 404194 266388
rect 404353 266386 404419 266389
rect 405038 266386 405044 266388
rect 404353 266384 405044 266386
rect 404353 266328 404358 266384
rect 404414 266328 405044 266384
rect 404353 266326 405044 266328
rect 404353 266323 404419 266326
rect 405038 266324 405044 266326
rect 405108 266324 405114 266388
rect 405733 266386 405799 266389
rect 406510 266386 406516 266388
rect 405733 266384 406516 266386
rect 405733 266328 405738 266384
rect 405794 266328 406516 266384
rect 405733 266326 406516 266328
rect 405733 266323 405799 266326
rect 406510 266324 406516 266326
rect 406580 266324 406586 266388
rect 407113 266386 407179 266389
rect 407614 266386 407620 266388
rect 407113 266384 407620 266386
rect 407113 266328 407118 266384
rect 407174 266328 407620 266384
rect 407113 266326 407620 266328
rect 407113 266323 407179 266326
rect 407614 266324 407620 266326
rect 407684 266324 407690 266388
rect 409873 266386 409939 266389
rect 411253 266388 411319 266389
rect 410006 266386 410012 266388
rect 409873 266384 410012 266386
rect 409873 266328 409878 266384
rect 409934 266328 410012 266384
rect 409873 266326 410012 266328
rect 409873 266323 409939 266326
rect 410006 266324 410012 266326
rect 410076 266324 410082 266388
rect 411253 266386 411300 266388
rect 411208 266384 411300 266386
rect 411208 266328 411258 266384
rect 411208 266326 411300 266328
rect 411253 266324 411300 266326
rect 411364 266324 411370 266388
rect 413001 266386 413067 266389
rect 418153 266388 418219 266389
rect 413318 266386 413324 266388
rect 413001 266384 413324 266386
rect 413001 266328 413006 266384
rect 413062 266328 413324 266384
rect 413001 266326 413324 266328
rect 411253 266323 411319 266324
rect 413001 266323 413067 266326
rect 413318 266324 413324 266326
rect 413388 266324 413394 266388
rect 418102 266324 418108 266388
rect 418172 266386 418219 266388
rect 419533 266386 419599 266389
rect 420678 266386 420684 266388
rect 418172 266384 418264 266386
rect 418214 266328 418264 266384
rect 418172 266326 418264 266328
rect 419533 266384 420684 266386
rect 419533 266328 419538 266384
rect 419594 266328 420684 266384
rect 419533 266326 420684 266328
rect 418172 266324 418219 266326
rect 418153 266323 418219 266324
rect 419533 266323 419599 266326
rect 420678 266324 420684 266326
rect 420748 266324 420754 266388
rect 420913 266386 420979 266389
rect 421782 266386 421788 266388
rect 420913 266384 421788 266386
rect 420913 266328 420918 266384
rect 420974 266328 421788 266384
rect 420913 266326 421788 266328
rect 420913 266323 420979 266326
rect 421782 266324 421788 266326
rect 421852 266324 421858 266388
rect 426433 266386 426499 266389
rect 427670 266386 427676 266388
rect 426433 266384 427676 266386
rect 426433 266328 426438 266384
rect 426494 266328 427676 266384
rect 426433 266326 427676 266328
rect 426433 266323 426499 266326
rect 427670 266324 427676 266326
rect 427740 266324 427746 266388
rect 436093 266386 436159 266389
rect 436870 266386 436876 266388
rect 436093 266384 436876 266386
rect 436093 266328 436098 266384
rect 436154 266328 436876 266384
rect 436093 266326 436876 266328
rect 436093 266323 436159 266326
rect 436870 266324 436876 266326
rect 436940 266324 436946 266388
rect 213453 266250 213519 266253
rect 272558 266250 272564 266252
rect 213453 266248 272564 266250
rect 213453 266192 213458 266248
rect 213514 266192 272564 266248
rect 213453 266190 272564 266192
rect 213453 266187 213519 266190
rect 272558 266188 272564 266190
rect 272628 266188 272634 266252
rect 215569 266114 215635 266117
rect 240542 266114 240548 266116
rect 215569 266112 240548 266114
rect 215569 266056 215574 266112
rect 215630 266056 240548 266112
rect 215569 266054 240548 266056
rect 215569 266051 215635 266054
rect 240542 266052 240548 266054
rect 240612 266052 240618 266116
rect 241646 265978 241652 265980
rect 219390 265918 241652 265978
rect 217869 265842 217935 265845
rect 219390 265842 219450 265918
rect 241646 265916 241652 265918
rect 241716 265916 241722 265980
rect 217869 265840 219450 265842
rect 217869 265784 217874 265840
rect 217930 265784 219450 265840
rect 217869 265782 219450 265784
rect 217869 265779 217935 265782
rect 209589 265706 209655 265709
rect 215845 265706 215911 265709
rect 239254 265706 239260 265708
rect 209589 265704 239260 265706
rect 209589 265648 209594 265704
rect 209650 265648 215850 265704
rect 215906 265648 239260 265704
rect 209589 265646 239260 265648
rect 209589 265643 209655 265646
rect 215845 265643 215911 265646
rect 239254 265644 239260 265646
rect 239324 265644 239330 265708
rect 379421 265706 379487 265709
rect 426382 265706 426388 265708
rect 379421 265704 426388 265706
rect 379421 265648 379426 265704
rect 379482 265648 426388 265704
rect 379421 265646 426388 265648
rect 379421 265643 379487 265646
rect 426382 265644 426388 265646
rect 426452 265644 426458 265708
rect 208209 265570 208275 265573
rect 209589 265570 209655 265573
rect 238150 265570 238156 265572
rect 208209 265568 238156 265570
rect 208209 265512 208214 265568
rect 208270 265512 209594 265568
rect 209650 265512 238156 265568
rect 208209 265510 238156 265512
rect 208209 265507 208275 265510
rect 209589 265507 209655 265510
rect 238150 265508 238156 265510
rect 238220 265508 238226 265572
rect 371601 265570 371667 265573
rect 373809 265570 373875 265573
rect 431166 265570 431172 265572
rect 371601 265568 431172 265570
rect 371601 265512 371606 265568
rect 371662 265512 373814 265568
rect 373870 265512 431172 265568
rect 371601 265510 431172 265512
rect 371601 265507 371667 265510
rect 373809 265507 373875 265510
rect 431166 265508 431172 265510
rect 431236 265508 431242 265572
rect 213361 265162 213427 265165
rect 215569 265162 215635 265165
rect 213361 265160 215635 265162
rect 213361 265104 213366 265160
rect 213422 265104 215574 265160
rect 215630 265104 215635 265160
rect 213361 265102 215635 265104
rect 213361 265099 213427 265102
rect 215569 265099 215635 265102
rect 371785 265162 371851 265165
rect 376201 265162 376267 265165
rect 388437 265162 388503 265165
rect 371785 265160 388503 265162
rect 371785 265104 371790 265160
rect 371846 265104 376206 265160
rect 376262 265104 388442 265160
rect 388498 265104 388503 265160
rect 371785 265102 388503 265104
rect 371785 265099 371851 265102
rect 376201 265099 376267 265102
rect 388437 265099 388503 265102
rect 214925 265026 214991 265029
rect 217869 265026 217935 265029
rect 214925 265024 217935 265026
rect 214925 264968 214930 265024
rect 214986 264968 217874 265024
rect 217930 264968 217935 265024
rect 214925 264966 217935 264968
rect 214925 264963 214991 264966
rect 217869 264963 217935 264966
rect 377121 265026 377187 265029
rect 377673 265026 377739 265029
rect 379421 265026 379487 265029
rect 379973 265026 380039 265029
rect 389173 265026 389239 265029
rect 377121 265024 379346 265026
rect 377121 264968 377126 265024
rect 377182 264968 377678 265024
rect 377734 264968 379346 265024
rect 377121 264966 379346 264968
rect 377121 264963 377187 264966
rect 377673 264963 377739 264966
rect 379286 264890 379346 264966
rect 379421 265024 380039 265026
rect 379421 264968 379426 265024
rect 379482 264968 379978 265024
rect 380034 264968 380039 265024
rect 379421 264966 380039 264968
rect 379421 264963 379487 264966
rect 379973 264963 380039 264966
rect 380206 265024 389239 265026
rect 380206 264968 389178 265024
rect 389234 264968 389239 265024
rect 380206 264966 389239 264968
rect 380206 264890 380266 264966
rect 389173 264963 389239 264966
rect 379286 264830 380266 264890
rect 57094 262244 57100 262308
rect 57164 262306 57170 262308
rect 57237 262306 57303 262309
rect 57164 262304 57303 262306
rect 57164 262248 57242 262304
rect 57298 262248 57303 262304
rect 57164 262246 57303 262248
rect 57164 262244 57170 262246
rect 57237 262243 57303 262246
rect 583520 258756 584960 258996
rect -960 254146 480 254236
rect -960 254086 6930 254146
rect -960 253996 480 254086
rect 6870 254010 6930 254086
rect 53046 254010 53052 254012
rect 6870 253950 53052 254010
rect 53046 253948 53052 253950
rect 53116 253948 53122 254012
rect 377990 250956 377996 251020
rect 378060 251018 378066 251020
rect 379421 251018 379487 251021
rect 378060 251016 379487 251018
rect 378060 250960 379426 251016
rect 379482 250960 379487 251016
rect 378060 250958 379487 250960
rect 378060 250956 378066 250958
rect 379421 250955 379487 250958
rect 178534 249868 178540 249932
rect 178604 249930 178610 249932
rect 179321 249930 179387 249933
rect 178604 249928 179387 249930
rect 178604 249872 179326 249928
rect 179382 249872 179387 249928
rect 178604 249870 179387 249872
rect 178604 249868 178610 249870
rect 179321 249867 179387 249870
rect 179638 249868 179644 249932
rect 179708 249930 179714 249932
rect 179781 249930 179847 249933
rect 190913 249932 190979 249933
rect 338481 249932 338547 249933
rect 190862 249930 190868 249932
rect 179708 249928 179847 249930
rect 179708 249872 179786 249928
rect 179842 249872 179847 249928
rect 179708 249870 179847 249872
rect 190822 249870 190868 249930
rect 190932 249928 190979 249932
rect 338430 249930 338436 249932
rect 190974 249872 190979 249928
rect 179708 249868 179714 249870
rect 179781 249867 179847 249870
rect 190862 249868 190868 249870
rect 190932 249868 190979 249872
rect 338390 249870 338436 249930
rect 338500 249928 338547 249932
rect 338542 249872 338547 249928
rect 338430 249868 338436 249870
rect 338500 249868 338547 249872
rect 339718 249868 339724 249932
rect 339788 249930 339794 249932
rect 340045 249930 340111 249933
rect 339788 249928 340111 249930
rect 339788 249872 340050 249928
rect 340106 249872 340111 249928
rect 339788 249870 340111 249872
rect 339788 249868 339794 249870
rect 190913 249867 190979 249868
rect 338481 249867 338547 249868
rect 340045 249867 340111 249870
rect 350942 249868 350948 249932
rect 351012 249930 351018 249932
rect 351729 249930 351795 249933
rect 351012 249928 351795 249930
rect 351012 249872 351734 249928
rect 351790 249872 351795 249928
rect 351012 249870 351795 249872
rect 351012 249868 351018 249870
rect 351729 249867 351795 249870
rect 498510 249868 498516 249932
rect 498580 249930 498586 249932
rect 499021 249930 499087 249933
rect 498580 249928 499087 249930
rect 498580 249872 499026 249928
rect 499082 249872 499087 249928
rect 498580 249870 499087 249872
rect 498580 249868 498586 249870
rect 499021 249867 499087 249870
rect 499798 249868 499804 249932
rect 499868 249930 499874 249932
rect 500033 249930 500099 249933
rect 510889 249932 510955 249933
rect 510838 249930 510844 249932
rect 499868 249928 500099 249930
rect 499868 249872 500038 249928
rect 500094 249872 500099 249928
rect 499868 249870 500099 249872
rect 510798 249870 510844 249930
rect 510908 249928 510955 249932
rect 510950 249872 510955 249928
rect 499868 249868 499874 249870
rect 500033 249867 500099 249870
rect 510838 249868 510844 249870
rect 510908 249868 510955 249872
rect 510889 249867 510955 249868
rect 44766 249732 44772 249796
rect 44836 249794 44842 249796
rect 58617 249794 58683 249797
rect 44836 249792 58683 249794
rect 44836 249736 58622 249792
rect 58678 249736 58683 249792
rect 44836 249734 58683 249736
rect 44836 249732 44842 249734
rect 58617 249731 58683 249734
rect 44950 249052 44956 249116
rect 45020 249114 45026 249116
rect 47853 249114 47919 249117
rect 85849 249114 85915 249117
rect 45020 249112 85915 249114
rect 45020 249056 47858 249112
rect 47914 249056 85854 249112
rect 85910 249056 85915 249112
rect 45020 249054 85915 249056
rect 45020 249052 45026 249054
rect 47853 249051 47919 249054
rect 85849 249051 85915 249054
rect 583520 245428 584960 245668
rect 196604 244218 197186 244220
rect 198733 244218 198799 244221
rect 199193 244218 199259 244221
rect 518893 244218 518959 244221
rect 519353 244218 519419 244221
rect 196604 244216 199259 244218
rect 196604 244160 198738 244216
rect 198794 244160 199198 244216
rect 199254 244160 199259 244216
rect 516558 244216 519419 244218
rect 197126 244158 199259 244160
rect 198733 244155 198799 244158
rect 199193 244155 199259 244158
rect 356562 243810 356622 244190
rect 516558 244160 518898 244216
rect 518954 244160 519358 244216
rect 519414 244160 519419 244216
rect 516558 244158 519419 244160
rect 518893 244155 518959 244158
rect 519353 244155 519419 244158
rect 358905 243810 358971 243813
rect 359365 243810 359431 243813
rect 356562 243808 359431 243810
rect 356562 243752 358910 243808
rect 358966 243752 359370 243808
rect 359426 243752 359431 243808
rect 356562 243750 359431 243752
rect 358905 243747 358971 243750
rect 359365 243747 359431 243750
rect -960 240940 480 241180
rect 580257 232386 580323 232389
rect 583520 232386 584960 232476
rect 580257 232384 584960 232386
rect 580257 232328 580262 232384
rect 580318 232328 584960 232384
rect 580257 232326 584960 232328
rect 580257 232323 580323 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect 376937 202874 377003 202877
rect 377581 202874 377647 202877
rect 376937 202872 377647 202874
rect 376937 202816 376942 202872
rect 376998 202816 377586 202872
rect 377642 202816 377647 202872
rect 376937 202814 377647 202816
rect 376937 202811 377003 202814
rect 377581 202811 377647 202814
rect -960 201922 480 202012
rect 3049 201922 3115 201925
rect -960 201920 3115 201922
rect -960 201864 3054 201920
rect 3110 201864 3115 201920
rect -960 201862 3115 201864
rect -960 201772 480 201862
rect 3049 201859 3115 201862
rect 57329 201922 57395 201925
rect 216673 201922 216739 201925
rect 217777 201922 217843 201925
rect 219390 201922 220064 201924
rect 57329 201920 60062 201922
rect 57329 201864 57334 201920
rect 57390 201864 60062 201920
rect 57329 201862 60062 201864
rect 216673 201920 220064 201922
rect 216673 201864 216678 201920
rect 216734 201864 217782 201920
rect 217838 201864 220064 201920
rect 377581 201922 377647 201925
rect 379470 201922 380052 201924
rect 377581 201920 380052 201922
rect 377581 201864 377586 201920
rect 377642 201864 380052 201920
rect 216673 201862 219450 201864
rect 377581 201862 379530 201864
rect 57329 201859 57395 201862
rect 216673 201859 216739 201862
rect 217777 201859 217843 201862
rect 377581 201859 377647 201862
rect 216765 201378 216831 201381
rect 217685 201378 217751 201381
rect 216765 201376 217751 201378
rect 216765 201320 216770 201376
rect 216826 201320 217690 201376
rect 217746 201320 217751 201376
rect 216765 201318 217751 201320
rect 216765 201315 216831 201318
rect 217685 201315 217751 201318
rect 57145 200970 57211 200973
rect 217685 200970 217751 200973
rect 219390 200970 220064 200972
rect 57145 200968 60062 200970
rect 57145 200912 57150 200968
rect 57206 200912 60062 200968
rect 57145 200910 60062 200912
rect 217685 200968 220064 200970
rect 217685 200912 217690 200968
rect 217746 200912 220064 200968
rect 377305 200970 377371 200973
rect 379470 200970 380052 200972
rect 377305 200968 380052 200970
rect 377305 200912 377310 200968
rect 377366 200912 380052 200968
rect 217685 200910 219450 200912
rect 377305 200910 379530 200912
rect 57145 200907 57211 200910
rect 217685 200907 217751 200910
rect 377305 200907 377371 200910
rect 56685 198794 56751 198797
rect 57605 198794 57671 198797
rect 217409 198794 217475 198797
rect 217777 198794 217843 198797
rect 219390 198794 220064 198796
rect 56685 198792 60062 198794
rect 56685 198736 56690 198792
rect 56746 198736 57610 198792
rect 57666 198736 60062 198792
rect 56685 198734 60062 198736
rect 217409 198792 220064 198794
rect 217409 198736 217414 198792
rect 217470 198736 217782 198792
rect 217838 198736 220064 198792
rect 376937 198794 377003 198797
rect 379470 198794 380052 198796
rect 376937 198792 380052 198794
rect 376937 198736 376942 198792
rect 376998 198736 380052 198792
rect 217409 198734 219450 198736
rect 376937 198734 379530 198736
rect 56685 198731 56751 198734
rect 57605 198731 57671 198734
rect 217409 198731 217475 198734
rect 217777 198731 217843 198734
rect 376937 198731 377003 198734
rect 217501 197842 217567 197845
rect 219390 197842 220064 197844
rect 217501 197840 220064 197842
rect 56777 197434 56843 197437
rect 57329 197434 57395 197437
rect 60002 197434 60062 197814
rect 217501 197784 217506 197840
rect 217562 197784 220064 197840
rect 377489 197842 377555 197845
rect 379470 197842 380052 197844
rect 377489 197840 380052 197842
rect 377489 197784 377494 197840
rect 377550 197784 380052 197840
rect 217501 197782 219450 197784
rect 377489 197782 379530 197784
rect 217501 197779 217567 197782
rect 377489 197779 377555 197782
rect 56777 197432 60062 197434
rect 56777 197376 56782 197432
rect 56838 197376 57334 197432
rect 57390 197376 60062 197432
rect 56777 197374 60062 197376
rect 216857 197434 216923 197437
rect 217501 197434 217567 197437
rect 216857 197432 217567 197434
rect 216857 197376 216862 197432
rect 216918 197376 217506 197432
rect 217562 197376 217567 197432
rect 216857 197374 217567 197376
rect 56777 197371 56843 197374
rect 57329 197371 57395 197374
rect 216857 197371 216923 197374
rect 217501 197371 217567 197374
rect 57421 196074 57487 196077
rect 57697 196074 57763 196077
rect 217041 196074 217107 196077
rect 217685 196074 217751 196077
rect 219390 196074 220064 196076
rect 57421 196072 60062 196074
rect 57421 196016 57426 196072
rect 57482 196016 57702 196072
rect 57758 196016 60062 196072
rect 57421 196014 60062 196016
rect 217041 196072 220064 196074
rect 217041 196016 217046 196072
rect 217102 196016 217690 196072
rect 217746 196016 220064 196072
rect 377029 196074 377095 196077
rect 377213 196074 377279 196077
rect 379470 196074 380052 196076
rect 377029 196072 380052 196074
rect 377029 196016 377034 196072
rect 377090 196016 377218 196072
rect 377274 196016 380052 196072
rect 217041 196014 219450 196016
rect 377029 196014 379530 196016
rect 57421 196011 57487 196014
rect 57697 196011 57763 196014
rect 217041 196011 217107 196014
rect 217685 196011 217751 196014
rect 377029 196011 377095 196014
rect 377213 196011 377279 196014
rect 57053 195258 57119 195261
rect 57421 195258 57487 195261
rect 57053 195256 60062 195258
rect 57053 195200 57058 195256
rect 57114 195200 57426 195256
rect 57482 195200 60062 195256
rect 57053 195198 60062 195200
rect 57053 195195 57119 195198
rect 57421 195195 57487 195198
rect 60002 194958 60062 195198
rect 217225 194986 217291 194989
rect 219390 194986 220064 194988
rect 217225 194984 220064 194986
rect 217225 194928 217230 194984
rect 217286 194928 220064 194984
rect 377765 194986 377831 194989
rect 379470 194986 380052 194988
rect 377765 194984 380052 194986
rect 377765 194928 377770 194984
rect 377826 194928 380052 194984
rect 217225 194926 219450 194928
rect 377765 194926 379530 194928
rect 217225 194923 217291 194926
rect 377765 194923 377831 194926
rect 57513 193218 57579 193221
rect 217593 193218 217659 193221
rect 219390 193218 220064 193220
rect 57513 193216 60062 193218
rect 57513 193160 57518 193216
rect 57574 193160 60062 193216
rect 57513 193158 60062 193160
rect 217593 193216 220064 193218
rect 217593 193160 217598 193216
rect 217654 193160 220064 193216
rect 377213 193218 377279 193221
rect 377857 193218 377923 193221
rect 379470 193218 380052 193220
rect 377213 193216 380052 193218
rect 377213 193160 377218 193216
rect 377274 193160 377862 193216
rect 377918 193160 380052 193216
rect 217593 193158 219450 193160
rect 377213 193158 379530 193160
rect 57513 193155 57579 193158
rect 217593 193155 217659 193158
rect 377213 193155 377279 193158
rect 377857 193155 377923 193158
rect 580349 192538 580415 192541
rect 583520 192538 584960 192628
rect 580349 192536 584960 192538
rect 580349 192480 580354 192536
rect 580410 192480 584960 192536
rect 580349 192478 584960 192480
rect 580349 192475 580415 192478
rect 583520 192388 584960 192478
rect -960 188716 480 188956
rect 359089 184922 359155 184925
rect 519261 184922 519327 184925
rect 519537 184922 519603 184925
rect 356562 184920 359155 184922
rect 356562 184864 359094 184920
rect 359150 184864 359155 184920
rect 356562 184862 359155 184864
rect 196604 184378 197186 184380
rect 199009 184378 199075 184381
rect 196604 184376 199075 184378
rect 196604 184320 199014 184376
rect 199070 184320 199075 184376
rect 356562 184350 356622 184862
rect 359089 184859 359155 184862
rect 516558 184920 519603 184922
rect 516558 184864 519266 184920
rect 519322 184864 519542 184920
rect 519598 184864 519603 184920
rect 516558 184862 519603 184864
rect 516558 184350 516618 184862
rect 519261 184859 519327 184862
rect 519537 184859 519603 184862
rect 197126 184318 199075 184320
rect 199009 184315 199075 184318
rect 198825 183562 198891 183565
rect 199377 183562 199443 183565
rect 198825 183560 199443 183562
rect 198825 183504 198830 183560
rect 198886 183504 199382 183560
rect 199438 183504 199443 183560
rect 198825 183502 199443 183504
rect 198825 183499 198891 183502
rect 199377 183499 199443 183502
rect 358905 183562 358971 183565
rect 359549 183562 359615 183565
rect 358905 183560 359615 183562
rect 358905 183504 358910 183560
rect 358966 183504 359554 183560
rect 359610 183504 359615 183560
rect 358905 183502 359615 183504
rect 358905 183499 358971 183502
rect 359549 183499 359615 183502
rect 196604 182746 197186 182748
rect 199377 182746 199443 182749
rect 358905 182746 358971 182749
rect 518985 182746 519051 182749
rect 519169 182746 519235 182749
rect 520181 182746 520247 182749
rect 196604 182744 199443 182746
rect 196604 182688 199382 182744
rect 199438 182688 199443 182744
rect 197126 182686 199443 182688
rect 356562 182744 358971 182746
rect 356562 182688 358910 182744
rect 358966 182688 358971 182744
rect 356562 182686 358971 182688
rect 516558 182744 520247 182746
rect 516558 182688 518990 182744
rect 519046 182688 519174 182744
rect 519230 182688 520186 182744
rect 520242 182688 520247 182744
rect 516558 182686 520247 182688
rect 199377 182683 199443 182686
rect 358905 182683 358971 182686
rect 518985 182683 519051 182686
rect 519169 182683 519235 182686
rect 520181 182683 520247 182686
rect 198825 182066 198891 182069
rect 199285 182066 199351 182069
rect 198825 182064 199351 182066
rect 198825 182008 198830 182064
rect 198886 182008 199290 182064
rect 199346 182008 199351 182064
rect 198825 182006 199351 182008
rect 198825 182003 198891 182006
rect 199285 182003 199351 182006
rect 196604 181386 197186 181388
rect 198825 181386 198891 181389
rect 359273 181386 359339 181389
rect 519537 181386 519603 181389
rect 196604 181384 198891 181386
rect 196604 181328 198830 181384
rect 198886 181328 198891 181384
rect 197126 181326 198891 181328
rect 356562 181384 359339 181386
rect 356562 181328 359278 181384
rect 359334 181328 359339 181384
rect 356562 181326 359339 181328
rect 516558 181384 519603 181386
rect 516558 181328 519542 181384
rect 519598 181328 519603 181384
rect 516558 181326 519603 181328
rect 198825 181323 198891 181326
rect 359273 181323 359339 181326
rect 519537 181323 519603 181326
rect 196558 179482 196618 179862
rect 198733 179482 198799 179485
rect 199101 179482 199167 179485
rect 196558 179480 199167 179482
rect 196558 179424 198738 179480
rect 198794 179424 199106 179480
rect 199162 179424 199167 179480
rect 196558 179422 199167 179424
rect 356562 179482 356622 179862
rect 359273 179482 359339 179485
rect 359457 179482 359523 179485
rect 356562 179480 359523 179482
rect 356562 179424 359278 179480
rect 359334 179424 359462 179480
rect 359518 179424 359523 179480
rect 356562 179422 359523 179424
rect 516558 179482 516618 179862
rect 518985 179482 519051 179485
rect 519445 179482 519511 179485
rect 516558 179480 519511 179482
rect 516558 179424 518990 179480
rect 519046 179424 519450 179480
rect 519506 179424 519511 179480
rect 516558 179422 519511 179424
rect 198733 179419 198799 179422
rect 199101 179419 199167 179422
rect 359273 179419 359339 179422
rect 359457 179419 359523 179422
rect 518985 179419 519051 179422
rect 519445 179419 519511 179422
rect 583520 179060 584960 179300
rect 518893 178802 518959 178805
rect 516558 178800 518959 178802
rect 516558 178744 518898 178800
rect 518954 178744 518959 178800
rect 516558 178742 518959 178744
rect 196604 178666 197186 178668
rect 198917 178666 198983 178669
rect 358997 178666 359063 178669
rect 196604 178664 198983 178666
rect 196604 178608 198922 178664
rect 198978 178608 198983 178664
rect 197126 178606 198983 178608
rect 356562 178664 359063 178666
rect 356562 178608 359002 178664
rect 359058 178608 359063 178664
rect 516558 178638 516618 178742
rect 518893 178739 518959 178742
rect 356562 178606 359063 178608
rect 198917 178603 198983 178606
rect 358997 178603 359063 178606
rect -960 175796 480 176036
rect 58985 175266 59051 175269
rect 58985 175264 60062 175266
rect 58985 175208 58990 175264
rect 59046 175208 60062 175264
rect 58985 175206 60062 175208
rect 58985 175203 59051 175206
rect 60002 174966 60062 175206
rect 200798 174932 200804 174996
rect 200868 174994 200874 174996
rect 219390 174994 220064 174996
rect 200868 174936 220064 174994
rect 376845 174994 376911 174997
rect 379470 174994 380052 174996
rect 376845 174992 380052 174994
rect 376845 174936 376850 174992
rect 376906 174936 380052 174992
rect 200868 174934 219450 174936
rect 376845 174934 379530 174936
rect 200868 174932 200874 174934
rect 376845 174931 376911 174934
rect 57881 173362 57947 173365
rect 59494 173362 60032 173364
rect 57881 173360 60032 173362
rect 57881 173304 57886 173360
rect 57942 173304 60032 173360
rect 216673 173362 216739 173365
rect 219390 173362 220064 173364
rect 216673 173360 220064 173362
rect 216673 173304 216678 173360
rect 216734 173304 220064 173360
rect 376845 173362 376911 173365
rect 379470 173362 380052 173364
rect 376845 173360 380052 173362
rect 376845 173304 376850 173360
rect 376906 173304 380052 173360
rect 57881 173302 59554 173304
rect 216673 173302 219450 173304
rect 376845 173302 379530 173304
rect 57881 173299 57947 173302
rect 216673 173299 216739 173302
rect 376845 173299 376911 173302
rect 57789 173090 57855 173093
rect 217041 173090 217107 173093
rect 219390 173090 220064 173092
rect 57789 173088 60062 173090
rect 57789 173032 57794 173088
rect 57850 173032 60062 173088
rect 57789 173030 60062 173032
rect 217041 173088 220064 173090
rect 217041 173032 217046 173088
rect 217102 173032 220064 173088
rect 377121 173090 377187 173093
rect 379470 173090 380052 173092
rect 377121 173088 380052 173090
rect 377121 173032 377126 173088
rect 377182 173032 380052 173088
rect 217041 173030 219450 173032
rect 377121 173030 379530 173032
rect 57789 173027 57855 173030
rect 217041 173027 217107 173030
rect 377121 173027 377187 173030
rect 583520 165732 584960 165972
rect 96061 164932 96127 164933
rect 115749 164932 115815 164933
rect 96061 164928 96108 164932
rect 96172 164930 96178 164932
rect 96061 164872 96066 164928
rect 96061 164868 96108 164872
rect 96172 164870 96218 164930
rect 115749 164928 115766 164932
rect 115830 164930 115836 164932
rect 412541 164930 412607 164933
rect 413456 164930 413462 164932
rect 115749 164872 115754 164928
rect 96172 164868 96178 164870
rect 115749 164868 115766 164872
rect 115830 164870 115906 164930
rect 412496 164928 413462 164930
rect 412496 164872 412546 164928
rect 412602 164872 413462 164928
rect 412496 164870 413462 164872
rect 115830 164868 115836 164870
rect 96061 164867 96127 164868
rect 115749 164867 115815 164868
rect 412541 164867 412607 164870
rect 413456 164868 413462 164870
rect 413526 164868 413532 164932
rect 138473 164796 138539 164797
rect 140865 164796 140931 164797
rect 143533 164796 143599 164797
rect 138472 164732 138478 164796
rect 138542 164794 138548 164796
rect 138542 164734 138630 164794
rect 140865 164792 140926 164796
rect 140865 164736 140870 164792
rect 138542 164732 138548 164734
rect 140865 164732 140926 164736
rect 140990 164794 140996 164796
rect 143504 164794 143510 164796
rect 140990 164734 141022 164794
rect 143442 164734 143510 164794
rect 143574 164792 143599 164796
rect 143594 164736 143599 164792
rect 140990 164732 140996 164734
rect 143504 164732 143510 164734
rect 143574 164732 143599 164736
rect 138473 164731 138539 164732
rect 140865 164731 140931 164732
rect 143533 164731 143599 164732
rect 163313 164796 163379 164797
rect 261017 164796 261083 164797
rect 425973 164796 426039 164797
rect 450997 164796 451063 164797
rect 163313 164792 163366 164796
rect 163430 164794 163436 164796
rect 163313 164736 163318 164792
rect 163313 164732 163366 164736
rect 163430 164734 163470 164794
rect 261017 164792 261078 164796
rect 261017 164736 261022 164792
rect 163430 164732 163436 164734
rect 261017 164732 261078 164736
rect 261142 164794 261148 164796
rect 425968 164794 425974 164796
rect 261142 164734 261174 164794
rect 425882 164734 425974 164794
rect 261142 164732 261148 164734
rect 425968 164732 425974 164734
rect 426038 164732 426044 164796
rect 450992 164794 450998 164796
rect 450906 164734 450998 164794
rect 450992 164732 450998 164734
rect 451062 164732 451068 164796
rect 163313 164731 163379 164732
rect 261017 164731 261083 164732
rect 425973 164731 426039 164732
rect 450997 164731 451063 164732
rect 84101 164658 84167 164661
rect 103513 164660 103579 164661
rect 105905 164660 105971 164661
rect 114369 164660 114435 164661
rect 118049 164660 118115 164661
rect 153377 164660 153443 164661
rect 165889 164660 165955 164661
rect 288249 164660 288315 164661
rect 305913 164660 305979 164661
rect 423489 164660 423555 164661
rect 429745 164660 429811 164661
rect 436921 164660 436987 164661
rect 470961 164660 471027 164661
rect 480897 164660 480963 164661
rect 85432 164658 85438 164660
rect 84101 164656 85438 164658
rect 84101 164600 84106 164656
rect 84162 164600 85438 164656
rect 84101 164598 85438 164600
rect 84101 164595 84167 164598
rect 85432 164596 85438 164598
rect 85502 164596 85508 164660
rect 103513 164656 103526 164660
rect 103590 164658 103596 164660
rect 103513 164600 103518 164656
rect 103513 164596 103526 164600
rect 103590 164598 103670 164658
rect 105905 164656 105974 164660
rect 105905 164600 105910 164656
rect 105966 164600 105974 164656
rect 103590 164596 103596 164598
rect 105905 164596 105974 164600
rect 106038 164658 106044 164660
rect 106038 164598 106062 164658
rect 114369 164656 114406 164660
rect 114470 164658 114476 164660
rect 114369 164600 114374 164656
rect 106038 164596 106044 164598
rect 114369 164596 114406 164600
rect 114470 164598 114526 164658
rect 118049 164656 118078 164660
rect 118142 164658 118148 164660
rect 118049 164600 118054 164656
rect 114470 164596 114476 164598
rect 118049 164596 118078 164600
rect 118142 164598 118206 164658
rect 153377 164656 153438 164660
rect 153377 164600 153382 164656
rect 118142 164596 118148 164598
rect 153377 164596 153438 164600
rect 153502 164658 153508 164660
rect 153502 164598 153534 164658
rect 165889 164656 165950 164660
rect 165889 164600 165894 164656
rect 153502 164596 153508 164598
rect 165889 164596 165950 164600
rect 166014 164658 166020 164660
rect 166014 164598 166046 164658
rect 288249 164656 288278 164660
rect 288342 164658 288348 164660
rect 288249 164600 288254 164656
rect 166014 164596 166020 164598
rect 288249 164596 288278 164600
rect 288342 164598 288406 164658
rect 305913 164656 305958 164660
rect 306022 164658 306028 164660
rect 305913 164600 305918 164656
rect 288342 164596 288348 164598
rect 305913 164596 305958 164600
rect 306022 164598 306070 164658
rect 306022 164596 306028 164598
rect 318464 164596 318470 164660
rect 318534 164596 318540 164660
rect 423489 164656 423526 164660
rect 423590 164658 423596 164660
rect 423489 164600 423494 164656
rect 423489 164596 423526 164600
rect 423590 164598 423646 164658
rect 429745 164656 429782 164660
rect 429846 164658 429852 164660
rect 429745 164600 429750 164656
rect 423590 164596 423596 164598
rect 429745 164596 429782 164600
rect 429846 164598 429902 164658
rect 436921 164656 436990 164660
rect 436921 164600 436926 164656
rect 436982 164600 436990 164656
rect 429846 164596 429852 164598
rect 436921 164596 436990 164600
rect 437054 164658 437060 164660
rect 437054 164598 437078 164658
rect 470961 164656 470990 164660
rect 471054 164658 471060 164660
rect 470961 164600 470966 164656
rect 437054 164596 437060 164598
rect 470961 164596 470990 164600
rect 471054 164598 471118 164658
rect 480897 164656 480918 164660
rect 480982 164658 480988 164660
rect 480897 164600 480902 164656
rect 471054 164596 471060 164598
rect 480897 164596 480918 164600
rect 480982 164598 481054 164658
rect 480982 164596 480988 164598
rect 103513 164595 103579 164596
rect 105905 164595 105971 164596
rect 114369 164595 114435 164596
rect 118049 164595 118115 164596
rect 153377 164595 153443 164596
rect 165889 164595 165955 164596
rect 288249 164595 288315 164596
rect 305913 164595 305979 164596
rect 265893 164524 265959 164525
rect 265893 164520 265940 164524
rect 266004 164522 266010 164524
rect 265893 164464 265898 164520
rect 265893 164460 265940 164464
rect 266004 164462 266050 164522
rect 266004 164460 266010 164462
rect 265893 164459 265959 164460
rect 205214 164324 205220 164388
rect 205284 164386 205290 164388
rect 290958 164386 290964 164388
rect 205284 164326 290964 164386
rect 205284 164324 205290 164326
rect 290958 164324 290964 164326
rect 291028 164324 291034 164388
rect 318472 164386 318532 164596
rect 423489 164595 423555 164596
rect 429745 164595 429811 164596
rect 436921 164595 436987 164596
rect 470961 164595 471027 164596
rect 480897 164595 480963 164596
rect 296670 164326 318532 164386
rect 98453 164252 98519 164253
rect 101029 164252 101095 164253
rect 108205 164252 108271 164253
rect 98453 164248 98500 164252
rect 98564 164250 98570 164252
rect 98453 164192 98458 164248
rect 98453 164188 98500 164192
rect 98564 164190 98610 164250
rect 101029 164248 101076 164252
rect 101140 164250 101146 164252
rect 101029 164192 101034 164248
rect 98564 164188 98570 164190
rect 101029 164188 101076 164192
rect 101140 164190 101186 164250
rect 108205 164248 108252 164252
rect 108316 164250 108322 164252
rect 122741 164250 122807 164253
rect 145925 164252 145991 164253
rect 148501 164252 148567 164253
rect 150893 164252 150959 164253
rect 123518 164250 123524 164252
rect 108205 164192 108210 164248
rect 101140 164188 101146 164190
rect 108205 164188 108252 164192
rect 108316 164190 108362 164250
rect 122696 164248 123524 164250
rect 122696 164192 122746 164248
rect 122802 164192 123524 164248
rect 122696 164190 123524 164192
rect 108316 164188 108322 164190
rect 98453 164187 98519 164188
rect 101029 164187 101095 164188
rect 108205 164187 108271 164188
rect 122741 164187 122807 164190
rect 123518 164188 123524 164190
rect 123588 164188 123594 164252
rect 145925 164248 145972 164252
rect 146036 164250 146042 164252
rect 145925 164192 145930 164248
rect 145925 164188 145972 164192
rect 146036 164190 146082 164250
rect 148501 164248 148548 164252
rect 148612 164250 148618 164252
rect 148501 164192 148506 164248
rect 146036 164188 146042 164190
rect 148501 164188 148548 164192
rect 148612 164190 148658 164250
rect 150893 164248 150940 164252
rect 151004 164250 151010 164252
rect 150893 164192 150898 164248
rect 148612 164188 148618 164190
rect 150893 164188 150940 164192
rect 151004 164190 151050 164250
rect 151004 164188 151010 164190
rect 203006 164188 203012 164252
rect 203076 164250 203082 164252
rect 296670 164250 296730 164326
rect 203076 164190 296730 164250
rect 298461 164252 298527 164253
rect 300853 164252 300919 164253
rect 303429 164252 303495 164253
rect 313365 164252 313431 164253
rect 418429 164252 418495 164253
rect 421005 164252 421071 164253
rect 428181 164252 428247 164253
rect 430941 164252 431007 164253
rect 473445 164252 473511 164253
rect 475837 164252 475903 164253
rect 478413 164252 478479 164253
rect 483381 164252 483447 164253
rect 298461 164248 298508 164252
rect 298572 164250 298578 164252
rect 298461 164192 298466 164248
rect 203076 164188 203082 164190
rect 298461 164188 298508 164192
rect 298572 164190 298618 164250
rect 300853 164248 300900 164252
rect 300964 164250 300970 164252
rect 300853 164192 300858 164248
rect 298572 164188 298578 164190
rect 300853 164188 300900 164192
rect 300964 164190 301010 164250
rect 303429 164248 303476 164252
rect 303540 164250 303546 164252
rect 303429 164192 303434 164248
rect 300964 164188 300970 164190
rect 303429 164188 303476 164192
rect 303540 164190 303586 164250
rect 313365 164248 313412 164252
rect 313476 164250 313482 164252
rect 313365 164192 313370 164248
rect 303540 164188 303546 164190
rect 313365 164188 313412 164192
rect 313476 164190 313522 164250
rect 418429 164248 418476 164252
rect 418540 164250 418546 164252
rect 418429 164192 418434 164248
rect 313476 164188 313482 164190
rect 418429 164188 418476 164192
rect 418540 164190 418586 164250
rect 421005 164248 421052 164252
rect 421116 164250 421122 164252
rect 421005 164192 421010 164248
rect 418540 164188 418546 164190
rect 421005 164188 421052 164192
rect 421116 164190 421162 164250
rect 428181 164248 428228 164252
rect 428292 164250 428298 164252
rect 428181 164192 428186 164248
rect 421116 164188 421122 164190
rect 428181 164188 428228 164192
rect 428292 164190 428338 164250
rect 430941 164248 430988 164252
rect 431052 164250 431058 164252
rect 430941 164192 430946 164248
rect 428292 164188 428298 164190
rect 430941 164188 430988 164192
rect 431052 164190 431098 164250
rect 473445 164248 473492 164252
rect 473556 164250 473562 164252
rect 473445 164192 473450 164248
rect 431052 164188 431058 164190
rect 473445 164188 473492 164192
rect 473556 164190 473602 164250
rect 475837 164248 475884 164252
rect 475948 164250 475954 164252
rect 475837 164192 475842 164248
rect 473556 164188 473562 164190
rect 475837 164188 475884 164192
rect 475948 164190 475994 164250
rect 478413 164248 478460 164252
rect 478524 164250 478530 164252
rect 478413 164192 478418 164248
rect 475948 164188 475954 164190
rect 478413 164188 478460 164192
rect 478524 164190 478570 164250
rect 483381 164248 483428 164252
rect 483492 164250 483498 164252
rect 483381 164192 483386 164248
rect 478524 164188 478530 164190
rect 483381 164188 483428 164192
rect 483492 164190 483538 164250
rect 483492 164188 483498 164190
rect 145925 164187 145991 164188
rect 148501 164187 148567 164188
rect 150893 164187 150959 164188
rect 298461 164187 298527 164188
rect 300853 164187 300919 164188
rect 303429 164187 303495 164188
rect 313365 164187 313431 164188
rect 418429 164187 418495 164188
rect 421005 164187 421071 164188
rect 428181 164187 428247 164188
rect 430941 164187 431007 164188
rect 473445 164187 473511 164188
rect 475837 164187 475903 164188
rect 478413 164187 478479 164188
rect 483381 164187 483447 164188
rect 198222 164052 198228 164116
rect 198292 164114 198298 164116
rect 308438 164114 308444 164116
rect 198292 164054 308444 164114
rect 198292 164052 198298 164054
rect 308438 164052 308444 164054
rect 308508 164052 308514 164116
rect 369301 164114 369367 164117
rect 485998 164114 486004 164116
rect 369301 164112 486004 164114
rect 369301 164056 369306 164112
rect 369362 164056 486004 164112
rect 369301 164054 486004 164056
rect 369301 164051 369367 164054
rect 485998 164052 486004 164054
rect 486068 164052 486074 164116
rect 111149 163980 111215 163981
rect 111149 163976 111196 163980
rect 111260 163978 111266 163980
rect 111149 163920 111154 163976
rect 111149 163916 111196 163920
rect 111260 163918 111306 163978
rect 111260 163916 111266 163918
rect 202454 163916 202460 163980
rect 202524 163978 202530 163980
rect 295926 163978 295932 163980
rect 202524 163918 295932 163978
rect 202524 163916 202530 163918
rect 295926 163916 295932 163918
rect 295996 163916 296002 163980
rect 111149 163915 111215 163916
rect 285949 163844 286015 163845
rect 196566 163780 196572 163844
rect 196636 163842 196642 163844
rect 270902 163842 270908 163844
rect 196636 163782 270908 163842
rect 196636 163780 196642 163782
rect 270902 163780 270908 163782
rect 270972 163780 270978 163844
rect 285949 163840 285996 163844
rect 286060 163842 286066 163844
rect 285949 163784 285954 163840
rect 285949 163780 285996 163784
rect 286060 163782 286106 163842
rect 286060 163780 286066 163782
rect 285949 163779 286015 163780
rect 113449 163708 113515 163709
rect 113398 163706 113404 163708
rect 113358 163646 113404 163706
rect 113468 163704 113515 163708
rect 113510 163648 113515 163704
rect 113398 163644 113404 163646
rect 113468 163644 113515 163648
rect 113449 163643 113515 163644
rect 218329 163706 218395 163709
rect 218830 163706 218836 163708
rect 218329 163704 218836 163706
rect 218329 163648 218334 163704
rect 218390 163648 218836 163704
rect 218329 163646 218836 163648
rect 218329 163643 218395 163646
rect 218830 163644 218836 163646
rect 218900 163644 218906 163708
rect 99373 163164 99439 163165
rect 128353 163164 128419 163165
rect 235993 163164 236059 163165
rect 95918 163100 95924 163164
rect 95988 163100 95994 163164
rect 99373 163160 99420 163164
rect 99484 163162 99490 163164
rect 128302 163162 128308 163164
rect 99373 163104 99378 163160
rect 99373 163100 99420 163104
rect 99484 163102 99530 163162
rect 128262 163102 128308 163162
rect 128372 163160 128419 163164
rect 235942 163162 235948 163164
rect 128414 163104 128419 163160
rect 99484 163100 99490 163102
rect 128302 163100 128308 163102
rect 128372 163100 128419 163104
rect 235902 163102 235948 163162
rect 236012 163160 236059 163164
rect 236054 163104 236059 163160
rect 235942 163100 235948 163102
rect 236012 163100 236059 163104
rect 261702 163100 261708 163164
rect 261772 163100 261778 163164
rect 264973 163162 265039 163165
rect 276105 163164 276171 163165
rect 265198 163162 265204 163164
rect 264973 163160 265204 163162
rect 264973 163104 264978 163160
rect 265034 163104 265204 163160
rect 264973 163102 265204 163104
rect -960 162740 480 162980
rect 76005 162756 76071 162757
rect 76005 162752 76052 162756
rect 76116 162754 76122 162756
rect 77293 162754 77359 162757
rect 78254 162754 78260 162756
rect 76005 162696 76010 162752
rect 76005 162692 76052 162696
rect 76116 162694 76162 162754
rect 77293 162752 78260 162754
rect 77293 162696 77298 162752
rect 77354 162696 78260 162752
rect 77293 162694 78260 162696
rect 76116 162692 76122 162694
rect 76005 162691 76071 162692
rect 77293 162691 77359 162694
rect 78254 162692 78260 162694
rect 78324 162692 78330 162756
rect 78673 162754 78739 162757
rect 79542 162754 79548 162756
rect 78673 162752 79548 162754
rect 78673 162696 78678 162752
rect 78734 162696 79548 162752
rect 78673 162694 79548 162696
rect 78673 162691 78739 162694
rect 79542 162692 79548 162694
rect 79612 162692 79618 162756
rect 80053 162754 80119 162757
rect 80462 162754 80468 162756
rect 80053 162752 80468 162754
rect 80053 162696 80058 162752
rect 80114 162696 80468 162752
rect 80053 162694 80468 162696
rect 80053 162691 80119 162694
rect 80462 162692 80468 162694
rect 80532 162692 80538 162756
rect 81433 162754 81499 162757
rect 81934 162754 81940 162756
rect 81433 162752 81940 162754
rect 81433 162696 81438 162752
rect 81494 162696 81940 162752
rect 81433 162694 81940 162696
rect 81433 162691 81499 162694
rect 81934 162692 81940 162694
rect 82004 162692 82010 162756
rect 82813 162754 82879 162757
rect 83038 162754 83044 162756
rect 82813 162752 83044 162754
rect 82813 162696 82818 162752
rect 82874 162696 83044 162752
rect 82813 162694 83044 162696
rect 82813 162691 82879 162694
rect 83038 162692 83044 162694
rect 83108 162692 83114 162756
rect 84193 162754 84259 162757
rect 84326 162754 84332 162756
rect 84193 162752 84332 162754
rect 84193 162696 84198 162752
rect 84254 162696 84332 162752
rect 84193 162694 84332 162696
rect 84193 162691 84259 162694
rect 84326 162692 84332 162694
rect 84396 162692 84402 162756
rect 85573 162754 85639 162757
rect 86534 162754 86540 162756
rect 85573 162752 86540 162754
rect 85573 162696 85578 162752
rect 85634 162696 86540 162752
rect 85573 162694 86540 162696
rect 85573 162691 85639 162694
rect 86534 162692 86540 162694
rect 86604 162692 86610 162756
rect 86953 162754 87019 162757
rect 87638 162754 87644 162756
rect 86953 162752 87644 162754
rect 86953 162696 86958 162752
rect 87014 162696 87644 162752
rect 86953 162694 87644 162696
rect 86953 162691 87019 162694
rect 87638 162692 87644 162694
rect 87708 162692 87714 162756
rect 88425 162754 88491 162757
rect 88742 162754 88748 162756
rect 88425 162752 88748 162754
rect 88425 162696 88430 162752
rect 88486 162696 88748 162752
rect 88425 162694 88748 162696
rect 88425 162691 88491 162694
rect 88742 162692 88748 162694
rect 88812 162692 88818 162756
rect 89805 162754 89871 162757
rect 90725 162756 90791 162757
rect 90030 162754 90036 162756
rect 89805 162752 90036 162754
rect 89805 162696 89810 162752
rect 89866 162696 90036 162752
rect 89805 162694 90036 162696
rect 89805 162691 89871 162694
rect 90030 162692 90036 162694
rect 90100 162692 90106 162756
rect 90725 162752 90772 162756
rect 90836 162754 90842 162756
rect 91185 162754 91251 162757
rect 91318 162754 91324 162756
rect 90725 162696 90730 162752
rect 90725 162692 90772 162696
rect 90836 162694 90882 162754
rect 91185 162752 91324 162754
rect 91185 162696 91190 162752
rect 91246 162696 91324 162752
rect 91185 162694 91324 162696
rect 90836 162692 90842 162694
rect 90725 162691 90791 162692
rect 91185 162691 91251 162694
rect 91318 162692 91324 162694
rect 91388 162692 91394 162756
rect 92473 162754 92539 162757
rect 93342 162754 93348 162756
rect 92473 162752 93348 162754
rect 92473 162696 92478 162752
rect 92534 162696 93348 162752
rect 92473 162694 93348 162696
rect 92473 162691 92539 162694
rect 93342 162692 93348 162694
rect 93412 162692 93418 162756
rect 93853 162754 93919 162757
rect 94446 162754 94452 162756
rect 93853 162752 94452 162754
rect 93853 162696 93858 162752
rect 93914 162696 94452 162752
rect 93853 162694 94452 162696
rect 93853 162691 93919 162694
rect 94446 162692 94452 162694
rect 94516 162692 94522 162756
rect 95233 162754 95299 162757
rect 95926 162754 95986 163100
rect 99373 163099 99439 163100
rect 128353 163099 128419 163100
rect 235993 163099 236059 163100
rect 95233 162752 95986 162754
rect 95233 162696 95238 162752
rect 95294 162696 95986 162752
rect 95233 162694 95986 162696
rect 96613 162754 96679 162757
rect 97022 162754 97028 162756
rect 96613 162752 97028 162754
rect 96613 162696 96618 162752
rect 96674 162696 97028 162752
rect 96613 162694 97028 162696
rect 95233 162691 95299 162694
rect 96613 162691 96679 162694
rect 97022 162692 97028 162694
rect 97092 162692 97098 162756
rect 97993 162754 98059 162757
rect 100753 162756 100819 162757
rect 98126 162754 98132 162756
rect 97993 162752 98132 162754
rect 97993 162696 97998 162752
rect 98054 162696 98132 162752
rect 97993 162694 98132 162696
rect 97993 162691 98059 162694
rect 98126 162692 98132 162694
rect 98196 162692 98202 162756
rect 100702 162754 100708 162756
rect 100662 162694 100708 162754
rect 100772 162752 100819 162756
rect 100814 162696 100819 162752
rect 100702 162692 100708 162694
rect 100772 162692 100819 162696
rect 100753 162691 100819 162692
rect 102133 162754 102199 162757
rect 103789 162756 103855 162757
rect 102726 162754 102732 162756
rect 102133 162752 102732 162754
rect 102133 162696 102138 162752
rect 102194 162696 102732 162752
rect 102133 162694 102732 162696
rect 102133 162691 102199 162694
rect 102726 162692 102732 162694
rect 102796 162692 102802 162756
rect 103789 162752 103836 162756
rect 103900 162754 103906 162756
rect 104893 162754 104959 162757
rect 105302 162754 105308 162756
rect 103789 162696 103794 162752
rect 103789 162692 103836 162696
rect 103900 162694 103946 162754
rect 104893 162752 105308 162754
rect 104893 162696 104898 162752
rect 104954 162696 105308 162752
rect 104893 162694 105308 162696
rect 103900 162692 103906 162694
rect 103789 162691 103855 162692
rect 104893 162691 104959 162694
rect 105302 162692 105308 162694
rect 105372 162692 105378 162756
rect 106273 162754 106339 162757
rect 106406 162754 106412 162756
rect 106273 162752 106412 162754
rect 106273 162696 106278 162752
rect 106334 162696 106412 162752
rect 106273 162694 106412 162696
rect 106273 162691 106339 162694
rect 106406 162692 106412 162694
rect 106476 162692 106482 162756
rect 107653 162754 107719 162757
rect 108614 162754 108620 162756
rect 107653 162752 108620 162754
rect 107653 162696 107658 162752
rect 107714 162696 108620 162752
rect 107653 162694 108620 162696
rect 107653 162691 107719 162694
rect 108614 162692 108620 162694
rect 108684 162692 108690 162756
rect 109534 162692 109540 162756
rect 109604 162754 109610 162756
rect 110505 162754 110571 162757
rect 109604 162752 110571 162754
rect 109604 162696 110510 162752
rect 110566 162696 110571 162752
rect 109604 162694 110571 162696
rect 109604 162692 109610 162694
rect 110505 162691 110571 162694
rect 110965 162756 111031 162757
rect 113173 162756 113239 162757
rect 110965 162752 111012 162756
rect 111076 162754 111082 162756
rect 110965 162696 110970 162752
rect 110965 162692 111012 162696
rect 111076 162694 111122 162754
rect 113173 162752 113220 162756
rect 113284 162754 113290 162756
rect 115933 162754 115999 162757
rect 118325 162756 118391 162757
rect 116894 162754 116900 162756
rect 113173 162696 113178 162752
rect 111076 162692 111082 162694
rect 113173 162692 113220 162696
rect 113284 162694 113330 162754
rect 115933 162752 116900 162754
rect 115933 162696 115938 162752
rect 115994 162696 116900 162752
rect 115933 162694 116900 162696
rect 113284 162692 113290 162694
rect 110965 162691 111031 162692
rect 113173 162691 113239 162692
rect 115933 162691 115999 162694
rect 116894 162692 116900 162694
rect 116964 162692 116970 162756
rect 118325 162752 118372 162756
rect 118436 162754 118442 162756
rect 118693 162754 118759 162757
rect 120717 162756 120783 162757
rect 125869 162756 125935 162757
rect 130837 162756 130903 162757
rect 133413 162756 133479 162757
rect 135989 162756 136055 162757
rect 155953 162756 156019 162757
rect 119102 162754 119108 162756
rect 118325 162696 118330 162752
rect 118325 162692 118372 162696
rect 118436 162694 118482 162754
rect 118693 162752 119108 162754
rect 118693 162696 118698 162752
rect 118754 162696 119108 162752
rect 118693 162694 119108 162696
rect 118436 162692 118442 162694
rect 118325 162691 118391 162692
rect 118693 162691 118759 162694
rect 119102 162692 119108 162694
rect 119172 162692 119178 162756
rect 120717 162752 120764 162756
rect 120828 162754 120834 162756
rect 120717 162696 120722 162752
rect 120717 162692 120764 162696
rect 120828 162694 120874 162754
rect 125869 162752 125916 162756
rect 125980 162754 125986 162756
rect 125869 162696 125874 162752
rect 120828 162692 120834 162694
rect 125869 162692 125916 162696
rect 125980 162694 126026 162754
rect 130837 162752 130884 162756
rect 130948 162754 130954 162756
rect 130837 162696 130842 162752
rect 125980 162692 125986 162694
rect 130837 162692 130884 162696
rect 130948 162694 130994 162754
rect 133413 162752 133460 162756
rect 133524 162754 133530 162756
rect 133413 162696 133418 162752
rect 130948 162692 130954 162694
rect 133413 162692 133460 162696
rect 133524 162694 133570 162754
rect 135989 162752 136036 162756
rect 136100 162754 136106 162756
rect 155902 162754 155908 162756
rect 135989 162696 135994 162752
rect 133524 162692 133530 162694
rect 135989 162692 136036 162696
rect 136100 162694 136146 162754
rect 155862 162694 155908 162754
rect 155972 162752 156019 162756
rect 156014 162696 156019 162752
rect 136100 162692 136106 162694
rect 155902 162692 155908 162694
rect 155972 162692 156019 162696
rect 120717 162691 120783 162692
rect 125869 162691 125935 162692
rect 130837 162691 130903 162692
rect 133413 162691 133479 162692
rect 135989 162691 136055 162692
rect 155953 162691 156019 162692
rect 183461 162756 183527 162757
rect 183461 162752 183508 162756
rect 183572 162754 183578 162756
rect 236085 162754 236151 162757
rect 237046 162754 237052 162756
rect 183461 162696 183466 162752
rect 183461 162692 183508 162696
rect 183572 162694 183618 162754
rect 236085 162752 237052 162754
rect 236085 162696 236090 162752
rect 236146 162696 237052 162752
rect 236085 162694 237052 162696
rect 183572 162692 183578 162694
rect 183461 162691 183527 162692
rect 236085 162691 236151 162694
rect 237046 162692 237052 162694
rect 237116 162692 237122 162756
rect 237373 162754 237439 162757
rect 238150 162754 238156 162756
rect 237373 162752 238156 162754
rect 237373 162696 237378 162752
rect 237434 162696 238156 162752
rect 237373 162694 238156 162696
rect 237373 162691 237439 162694
rect 238150 162692 238156 162694
rect 238220 162692 238226 162756
rect 240133 162754 240199 162757
rect 240542 162754 240548 162756
rect 240133 162752 240548 162754
rect 240133 162696 240138 162752
rect 240194 162696 240548 162752
rect 240133 162694 240548 162696
rect 240133 162691 240199 162694
rect 240542 162692 240548 162694
rect 240612 162692 240618 162756
rect 241513 162754 241579 162757
rect 242893 162756 242959 162757
rect 241646 162754 241652 162756
rect 241513 162752 241652 162754
rect 241513 162696 241518 162752
rect 241574 162696 241652 162752
rect 241513 162694 241652 162696
rect 241513 162691 241579 162694
rect 241646 162692 241652 162694
rect 241716 162692 241722 162756
rect 242893 162752 242940 162756
rect 243004 162754 243010 162756
rect 242893 162696 242898 162752
rect 242893 162692 242940 162696
rect 243004 162694 243050 162754
rect 243004 162692 243010 162694
rect 244222 162692 244228 162756
rect 244292 162754 244298 162756
rect 244365 162754 244431 162757
rect 244292 162752 244431 162754
rect 244292 162696 244370 162752
rect 244426 162696 244431 162752
rect 244292 162694 244431 162696
rect 244292 162692 244298 162694
rect 242893 162691 242959 162692
rect 244365 162691 244431 162694
rect 245653 162754 245719 162757
rect 246430 162754 246436 162756
rect 245653 162752 246436 162754
rect 245653 162696 245658 162752
rect 245714 162696 246436 162752
rect 245653 162694 246436 162696
rect 245653 162691 245719 162694
rect 246430 162692 246436 162694
rect 246500 162692 246506 162756
rect 247033 162754 247099 162757
rect 248229 162756 248295 162757
rect 247718 162754 247724 162756
rect 247033 162752 247724 162754
rect 247033 162696 247038 162752
rect 247094 162696 247724 162752
rect 247033 162694 247724 162696
rect 247033 162691 247099 162694
rect 247718 162692 247724 162694
rect 247788 162692 247794 162756
rect 248229 162754 248276 162756
rect 248184 162752 248276 162754
rect 248184 162696 248234 162752
rect 248184 162694 248276 162696
rect 248229 162692 248276 162694
rect 248340 162692 248346 162756
rect 248413 162754 248479 162757
rect 248638 162754 248644 162756
rect 248413 162752 248644 162754
rect 248413 162696 248418 162752
rect 248474 162696 248644 162752
rect 248413 162694 248644 162696
rect 248229 162691 248295 162692
rect 248413 162691 248479 162694
rect 248638 162692 248644 162694
rect 248708 162692 248714 162756
rect 249793 162754 249859 162757
rect 250621 162756 250687 162757
rect 251173 162756 251239 162757
rect 250110 162754 250116 162756
rect 249793 162752 250116 162754
rect 249793 162696 249798 162752
rect 249854 162696 250116 162752
rect 249793 162694 250116 162696
rect 249793 162691 249859 162694
rect 250110 162692 250116 162694
rect 250180 162692 250186 162756
rect 250621 162752 250668 162756
rect 250732 162754 250738 162756
rect 250621 162696 250626 162752
rect 250621 162692 250668 162696
rect 250732 162694 250778 162754
rect 251173 162752 251220 162756
rect 251284 162754 251290 162756
rect 252553 162754 252619 162757
rect 253565 162756 253631 162757
rect 253422 162754 253428 162756
rect 251173 162696 251178 162752
rect 250732 162692 250738 162694
rect 251173 162692 251220 162696
rect 251284 162694 251330 162754
rect 252553 162752 253428 162754
rect 252553 162696 252558 162752
rect 252614 162696 253428 162752
rect 252553 162694 253428 162696
rect 251284 162692 251290 162694
rect 250621 162691 250687 162692
rect 251173 162691 251239 162692
rect 252553 162691 252619 162694
rect 253422 162692 253428 162694
rect 253492 162692 253498 162756
rect 253565 162752 253612 162756
rect 253676 162754 253682 162756
rect 253933 162754 253999 162757
rect 254526 162754 254532 162756
rect 253565 162696 253570 162752
rect 253565 162692 253612 162696
rect 253676 162694 253722 162754
rect 253933 162752 254532 162754
rect 253933 162696 253938 162752
rect 253994 162696 254532 162752
rect 253933 162694 254532 162696
rect 253676 162692 253682 162694
rect 253565 162691 253631 162692
rect 253933 162691 253999 162694
rect 254526 162692 254532 162694
rect 254596 162692 254602 162756
rect 255313 162754 255379 162757
rect 256141 162756 256207 162757
rect 255814 162754 255820 162756
rect 255313 162752 255820 162754
rect 255313 162696 255318 162752
rect 255374 162696 255820 162752
rect 255313 162694 255820 162696
rect 255313 162691 255379 162694
rect 255814 162692 255820 162694
rect 255884 162692 255890 162756
rect 256141 162752 256188 162756
rect 256252 162754 256258 162756
rect 256693 162754 256759 162757
rect 258349 162756 258415 162757
rect 259453 162756 259519 162757
rect 256918 162754 256924 162756
rect 256141 162696 256146 162752
rect 256141 162692 256188 162696
rect 256252 162694 256298 162754
rect 256693 162752 256924 162754
rect 256693 162696 256698 162752
rect 256754 162696 256924 162752
rect 256693 162694 256924 162696
rect 256252 162692 256258 162694
rect 256141 162691 256207 162692
rect 256693 162691 256759 162694
rect 256918 162692 256924 162694
rect 256988 162692 256994 162756
rect 258349 162752 258396 162756
rect 258460 162754 258466 162756
rect 258349 162696 258354 162752
rect 258349 162692 258396 162696
rect 258460 162694 258506 162754
rect 259453 162752 259500 162756
rect 259564 162754 259570 162756
rect 260833 162754 260899 162757
rect 261710 162754 261770 163100
rect 264973 163099 265039 163102
rect 265198 163100 265204 163102
rect 265268 163100 265274 163164
rect 272190 163100 272196 163164
rect 272260 163100 272266 163164
rect 276054 163162 276060 163164
rect 276014 163102 276060 163162
rect 276124 163160 276171 163164
rect 276166 163104 276171 163160
rect 276054 163100 276060 163102
rect 276124 163100 276171 163104
rect 398230 163100 398236 163164
rect 398300 163100 398306 163164
rect 401593 163162 401659 163165
rect 416037 163164 416103 163165
rect 455781 163164 455847 163165
rect 401726 163162 401732 163164
rect 401593 163160 401732 163162
rect 401593 163104 401598 163160
rect 401654 163104 401732 163160
rect 401593 163102 401732 163104
rect 263542 162828 263548 162892
rect 263612 162890 263618 162892
rect 263685 162890 263751 162893
rect 263612 162888 263751 162890
rect 263612 162832 263690 162888
rect 263746 162832 263751 162888
rect 263612 162830 263751 162832
rect 263612 162828 263618 162830
rect 263685 162827 263751 162830
rect 268285 162892 268351 162893
rect 268285 162888 268332 162892
rect 268396 162890 268402 162892
rect 268285 162832 268290 162888
rect 268285 162828 268332 162832
rect 268396 162830 268442 162890
rect 268396 162828 268402 162830
rect 268285 162827 268351 162828
rect 259453 162696 259458 162752
rect 258460 162692 258466 162694
rect 259453 162692 259500 162696
rect 259564 162694 259610 162754
rect 260833 162752 261770 162754
rect 260833 162696 260838 162752
rect 260894 162696 261770 162752
rect 260833 162694 261770 162696
rect 262213 162754 262279 162757
rect 262806 162754 262812 162756
rect 262213 162752 262812 162754
rect 262213 162696 262218 162752
rect 262274 162696 262812 162752
rect 262213 162694 262812 162696
rect 259564 162692 259570 162694
rect 258349 162691 258415 162692
rect 259453 162691 259519 162692
rect 260833 162691 260899 162694
rect 262213 162691 262279 162694
rect 262806 162692 262812 162694
rect 262876 162692 262882 162756
rect 263593 162754 263659 162757
rect 266353 162756 266419 162757
rect 263910 162754 263916 162756
rect 263593 162752 263916 162754
rect 263593 162696 263598 162752
rect 263654 162696 263916 162752
rect 263593 162694 263916 162696
rect 263593 162691 263659 162694
rect 263910 162692 263916 162694
rect 263980 162692 263986 162756
rect 266302 162754 266308 162756
rect 266262 162694 266308 162754
rect 266372 162752 266419 162756
rect 267549 162756 267615 162757
rect 267549 162754 267596 162756
rect 266414 162696 266419 162752
rect 266302 162692 266308 162694
rect 266372 162692 266419 162696
rect 267504 162752 267596 162754
rect 267504 162696 267554 162752
rect 267504 162694 267596 162696
rect 266353 162691 266419 162692
rect 267549 162692 267596 162694
rect 267660 162692 267666 162756
rect 267733 162754 267799 162757
rect 268694 162754 268700 162756
rect 267733 162752 268700 162754
rect 267733 162696 267738 162752
rect 267794 162696 268700 162752
rect 267733 162694 268700 162696
rect 267549 162691 267615 162692
rect 267733 162691 267799 162694
rect 268694 162692 268700 162694
rect 268764 162692 268770 162756
rect 269113 162754 269179 162757
rect 269798 162754 269804 162756
rect 269113 162752 269804 162754
rect 269113 162696 269118 162752
rect 269174 162696 269804 162752
rect 269113 162694 269804 162696
rect 269113 162691 269179 162694
rect 269798 162692 269804 162694
rect 269868 162692 269874 162756
rect 270493 162754 270559 162757
rect 271086 162754 271092 162756
rect 270493 162752 271092 162754
rect 270493 162696 270498 162752
rect 270554 162696 271092 162752
rect 270493 162694 271092 162696
rect 270493 162691 270559 162694
rect 271086 162692 271092 162694
rect 271156 162692 271162 162756
rect 271873 162754 271939 162757
rect 272198 162754 272258 163100
rect 276105 163099 276171 163100
rect 273437 162892 273503 162893
rect 273437 162888 273484 162892
rect 273548 162890 273554 162892
rect 273437 162832 273442 162888
rect 273437 162828 273484 162832
rect 273548 162830 273594 162890
rect 273548 162828 273554 162830
rect 273437 162827 273503 162828
rect 271873 162752 272258 162754
rect 271873 162696 271878 162752
rect 271934 162696 272258 162752
rect 271873 162694 272258 162696
rect 273253 162754 273319 162757
rect 274398 162754 274404 162756
rect 273253 162752 274404 162754
rect 273253 162696 273258 162752
rect 273314 162696 274404 162752
rect 273253 162694 274404 162696
rect 271873 162691 271939 162694
rect 273253 162691 273319 162694
rect 274398 162692 274404 162694
rect 274468 162692 274474 162756
rect 274817 162754 274883 162757
rect 275318 162754 275324 162756
rect 274817 162752 275324 162754
rect 274817 162696 274822 162752
rect 274878 162696 275324 162752
rect 274817 162694 275324 162696
rect 274817 162691 274883 162694
rect 275318 162692 275324 162694
rect 275388 162692 275394 162756
rect 276013 162754 276079 162757
rect 276974 162754 276980 162756
rect 276013 162752 276980 162754
rect 276013 162696 276018 162752
rect 276074 162696 276980 162752
rect 276013 162694 276980 162696
rect 276013 162691 276079 162694
rect 276974 162692 276980 162694
rect 277044 162692 277050 162756
rect 278998 162692 279004 162756
rect 279068 162754 279074 162756
rect 280061 162754 280127 162757
rect 279068 162752 280127 162754
rect 279068 162696 280066 162752
rect 280122 162696 280127 162752
rect 279068 162694 280127 162696
rect 279068 162692 279074 162694
rect 280061 162691 280127 162694
rect 280797 162756 280863 162757
rect 283741 162756 283807 162757
rect 280797 162752 280844 162756
rect 280908 162754 280914 162756
rect 280797 162696 280802 162752
rect 280797 162692 280844 162696
rect 280908 162694 280954 162754
rect 283741 162752 283788 162756
rect 283852 162754 283858 162756
rect 293217 162754 293283 162757
rect 320909 162756 320975 162757
rect 343449 162756 343515 162757
rect 396073 162756 396139 162757
rect 293350 162754 293356 162756
rect 283741 162696 283746 162752
rect 280908 162692 280914 162694
rect 283741 162692 283788 162696
rect 283852 162694 283898 162754
rect 293217 162752 293356 162754
rect 293217 162696 293222 162752
rect 293278 162696 293356 162752
rect 293217 162694 293356 162696
rect 283852 162692 283858 162694
rect 280797 162691 280863 162692
rect 283741 162691 283807 162692
rect 293217 162691 293283 162694
rect 293350 162692 293356 162694
rect 293420 162692 293426 162756
rect 320909 162752 320956 162756
rect 321020 162754 321026 162756
rect 343398 162754 343404 162756
rect 320909 162696 320914 162752
rect 320909 162692 320956 162696
rect 321020 162694 321066 162754
rect 343358 162694 343404 162754
rect 343468 162752 343515 162756
rect 396022 162754 396028 162756
rect 343510 162696 343515 162752
rect 321020 162692 321026 162694
rect 343398 162692 343404 162694
rect 343468 162692 343515 162696
rect 395982 162694 396028 162754
rect 396092 162752 396139 162756
rect 396134 162696 396139 162752
rect 396022 162692 396028 162694
rect 396092 162692 396139 162696
rect 320909 162691 320975 162692
rect 343449 162691 343515 162692
rect 396073 162691 396139 162692
rect 397453 162754 397519 162757
rect 398238 162754 398298 163100
rect 401593 163099 401659 163102
rect 401726 163100 401732 163102
rect 401796 163100 401802 163164
rect 416037 163160 416084 163164
rect 416148 163162 416154 163164
rect 416037 163104 416042 163160
rect 416037 163100 416084 163104
rect 416148 163102 416194 163162
rect 455781 163160 455828 163164
rect 455892 163162 455898 163164
rect 455781 163104 455786 163160
rect 416148 163100 416154 163102
rect 455781 163100 455828 163104
rect 455892 163102 455938 163162
rect 455892 163100 455898 163102
rect 416037 163099 416103 163100
rect 455781 163099 455847 163100
rect 397453 162752 398298 162754
rect 397453 162696 397458 162752
rect 397514 162696 398298 162752
rect 397453 162694 398298 162696
rect 398833 162754 398899 162757
rect 399518 162754 399524 162756
rect 398833 162752 399524 162754
rect 398833 162696 398838 162752
rect 398894 162696 399524 162752
rect 398833 162694 399524 162696
rect 397453 162691 397519 162694
rect 398833 162691 398899 162694
rect 399518 162692 399524 162694
rect 399588 162692 399594 162756
rect 400213 162754 400279 162757
rect 403065 162756 403131 162757
rect 400438 162754 400444 162756
rect 400213 162752 400444 162754
rect 400213 162696 400218 162752
rect 400274 162696 400444 162752
rect 400213 162694 400444 162696
rect 400213 162691 400279 162694
rect 400438 162692 400444 162694
rect 400508 162692 400514 162756
rect 403014 162754 403020 162756
rect 402974 162694 403020 162754
rect 403084 162752 403131 162756
rect 403126 162696 403131 162752
rect 403014 162692 403020 162694
rect 403084 162692 403131 162696
rect 403065 162691 403131 162692
rect 404353 162754 404419 162757
rect 405038 162754 405044 162756
rect 404353 162752 405044 162754
rect 404353 162696 404358 162752
rect 404414 162696 405044 162752
rect 404353 162694 405044 162696
rect 404353 162691 404419 162694
rect 405038 162692 405044 162694
rect 405108 162692 405114 162756
rect 405733 162754 405799 162757
rect 406510 162754 406516 162756
rect 405733 162752 406516 162754
rect 405733 162696 405738 162752
rect 405794 162696 406516 162752
rect 405733 162694 406516 162696
rect 405733 162691 405799 162694
rect 406510 162692 406516 162694
rect 406580 162692 406586 162756
rect 407205 162754 407271 162757
rect 408309 162756 408375 162757
rect 407614 162754 407620 162756
rect 407205 162752 407620 162754
rect 407205 162696 407210 162752
rect 407266 162696 407620 162752
rect 407205 162694 407620 162696
rect 407205 162691 407271 162694
rect 407614 162692 407620 162694
rect 407684 162692 407690 162756
rect 408309 162754 408356 162756
rect 408264 162752 408356 162754
rect 408264 162696 408314 162752
rect 408264 162694 408356 162696
rect 408309 162692 408356 162694
rect 408420 162692 408426 162756
rect 408493 162754 408559 162757
rect 408718 162754 408724 162756
rect 408493 162752 408724 162754
rect 408493 162696 408498 162752
rect 408554 162696 408724 162752
rect 408493 162694 408724 162696
rect 408309 162691 408375 162692
rect 408493 162691 408559 162694
rect 408718 162692 408724 162694
rect 408788 162692 408794 162756
rect 409873 162754 409939 162757
rect 410006 162754 410012 162756
rect 409873 162752 410012 162754
rect 409873 162696 409878 162752
rect 409934 162696 410012 162752
rect 409873 162694 410012 162696
rect 409873 162691 409939 162694
rect 410006 162692 410012 162694
rect 410076 162692 410082 162756
rect 410609 162754 410675 162757
rect 411345 162756 411411 162757
rect 410742 162754 410748 162756
rect 410609 162752 410748 162754
rect 410609 162696 410614 162752
rect 410670 162696 410748 162752
rect 410609 162694 410748 162696
rect 410609 162691 410675 162694
rect 410742 162692 410748 162694
rect 410812 162692 410818 162756
rect 411294 162754 411300 162756
rect 411254 162694 411300 162754
rect 411364 162752 411411 162756
rect 411406 162696 411411 162752
rect 411294 162692 411300 162694
rect 411364 162692 411411 162696
rect 411345 162691 411411 162692
rect 413553 162754 413619 162757
rect 413686 162754 413692 162756
rect 413553 162752 413692 162754
rect 413553 162696 413558 162752
rect 413614 162696 413692 162752
rect 413553 162694 413692 162696
rect 413553 162691 413619 162694
rect 413686 162692 413692 162694
rect 413756 162692 413762 162756
rect 414013 162754 414079 162757
rect 415485 162756 415551 162757
rect 414606 162754 414612 162756
rect 414013 162752 414612 162754
rect 414013 162696 414018 162752
rect 414074 162696 414612 162752
rect 414013 162694 414612 162696
rect 414013 162691 414079 162694
rect 414606 162692 414612 162694
rect 414676 162692 414682 162756
rect 415485 162752 415532 162756
rect 415596 162754 415602 162756
rect 416773 162754 416839 162757
rect 416998 162754 417004 162756
rect 415485 162696 415490 162752
rect 415485 162692 415532 162696
rect 415596 162694 415642 162754
rect 416773 162752 417004 162754
rect 416773 162696 416778 162752
rect 416834 162696 417004 162752
rect 416773 162694 417004 162696
rect 415596 162692 415602 162694
rect 415485 162691 415551 162692
rect 416773 162691 416839 162694
rect 416998 162692 417004 162694
rect 417068 162692 417074 162756
rect 418153 162754 418219 162757
rect 419206 162754 419212 162756
rect 418153 162752 419212 162754
rect 418153 162696 418158 162752
rect 418214 162696 419212 162752
rect 418153 162694 419212 162696
rect 418153 162691 418219 162694
rect 419206 162692 419212 162694
rect 419276 162692 419282 162756
rect 419533 162754 419599 162757
rect 420678 162754 420684 162756
rect 419533 162752 420684 162754
rect 419533 162696 419538 162752
rect 419594 162696 420684 162752
rect 419533 162694 420684 162696
rect 419533 162691 419599 162694
rect 420678 162692 420684 162694
rect 420748 162692 420754 162756
rect 420913 162754 420979 162757
rect 421782 162754 421788 162756
rect 420913 162752 421788 162754
rect 420913 162696 420918 162752
rect 420974 162696 421788 162752
rect 420913 162694 421788 162696
rect 420913 162691 420979 162694
rect 421782 162692 421788 162694
rect 421852 162692 421858 162756
rect 422293 162754 422359 162757
rect 422886 162754 422892 162756
rect 422293 162752 422892 162754
rect 422293 162696 422298 162752
rect 422354 162696 422892 162752
rect 422293 162694 422892 162696
rect 422293 162691 422359 162694
rect 422886 162692 422892 162694
rect 422956 162692 422962 162756
rect 423673 162754 423739 162757
rect 423990 162754 423996 162756
rect 423673 162752 423996 162754
rect 423673 162696 423678 162752
rect 423734 162696 423996 162752
rect 423673 162694 423996 162696
rect 423673 162691 423739 162694
rect 423990 162692 423996 162694
rect 424060 162692 424066 162756
rect 425053 162754 425119 162757
rect 426433 162756 426499 162757
rect 425278 162754 425284 162756
rect 425053 162752 425284 162754
rect 425053 162696 425058 162752
rect 425114 162696 425284 162752
rect 425053 162694 425284 162696
rect 425053 162691 425119 162694
rect 425278 162692 425284 162694
rect 425348 162692 425354 162756
rect 426382 162754 426388 162756
rect 426342 162694 426388 162754
rect 426452 162752 426499 162756
rect 426494 162696 426499 162752
rect 426382 162692 426388 162694
rect 426452 162692 426499 162696
rect 428774 162692 428780 162756
rect 428844 162754 428850 162756
rect 429101 162754 429167 162757
rect 428844 162752 429167 162754
rect 428844 162696 429106 162752
rect 429162 162696 429167 162752
rect 428844 162694 429167 162696
rect 428844 162692 428850 162694
rect 426433 162691 426499 162692
rect 429101 162691 429167 162694
rect 430573 162754 430639 162757
rect 431166 162754 431172 162756
rect 430573 162752 431172 162754
rect 430573 162696 430578 162752
rect 430634 162696 431172 162752
rect 430573 162694 431172 162696
rect 430573 162691 430639 162694
rect 431166 162692 431172 162694
rect 431236 162692 431242 162756
rect 431718 162692 431724 162756
rect 431788 162754 431794 162756
rect 431953 162754 432019 162757
rect 431788 162752 432019 162754
rect 431788 162696 431958 162752
rect 432014 162696 432019 162752
rect 431788 162694 432019 162696
rect 431788 162692 431794 162694
rect 431953 162691 432019 162694
rect 433333 162754 433399 162757
rect 435725 162756 435791 162757
rect 435909 162756 435975 162757
rect 434662 162754 434668 162756
rect 433333 162752 434668 162754
rect 433333 162696 433338 162752
rect 433394 162696 434668 162752
rect 433333 162694 434668 162696
rect 433333 162691 433399 162694
rect 434662 162692 434668 162694
rect 434732 162692 434738 162756
rect 435725 162754 435772 162756
rect 435680 162752 435772 162754
rect 435680 162696 435730 162752
rect 435680 162694 435772 162696
rect 435725 162692 435772 162694
rect 435836 162692 435842 162756
rect 435909 162752 435956 162756
rect 436020 162754 436026 162756
rect 437473 162754 437539 162757
rect 438485 162756 438551 162757
rect 438342 162754 438348 162756
rect 435909 162696 435914 162752
rect 435909 162692 435956 162696
rect 436020 162694 436066 162754
rect 437473 162752 438348 162754
rect 437473 162696 437478 162752
rect 437534 162696 438348 162752
rect 437473 162694 438348 162696
rect 436020 162692 436026 162694
rect 435725 162691 435791 162692
rect 435909 162691 435975 162692
rect 437473 162691 437539 162694
rect 438342 162692 438348 162694
rect 438412 162692 438418 162756
rect 438485 162752 438532 162756
rect 438596 162754 438602 162756
rect 438853 162754 438919 162757
rect 440877 162756 440943 162757
rect 443453 162756 443519 162757
rect 445845 162756 445911 162757
rect 448237 162756 448303 162757
rect 453389 162756 453455 162757
rect 458357 162756 458423 162757
rect 439078 162754 439084 162756
rect 438485 162696 438490 162752
rect 438485 162692 438532 162696
rect 438596 162694 438642 162754
rect 438853 162752 439084 162754
rect 438853 162696 438858 162752
rect 438914 162696 439084 162752
rect 438853 162694 439084 162696
rect 438596 162692 438602 162694
rect 438485 162691 438551 162692
rect 438853 162691 438919 162694
rect 439078 162692 439084 162694
rect 439148 162692 439154 162756
rect 440877 162752 440924 162756
rect 440988 162754 440994 162756
rect 440877 162696 440882 162752
rect 440877 162692 440924 162696
rect 440988 162694 441034 162754
rect 443453 162752 443500 162756
rect 443564 162754 443570 162756
rect 443453 162696 443458 162752
rect 440988 162692 440994 162694
rect 443453 162692 443500 162696
rect 443564 162694 443610 162754
rect 445845 162752 445892 162756
rect 445956 162754 445962 162756
rect 445845 162696 445850 162752
rect 443564 162692 443570 162694
rect 445845 162692 445892 162696
rect 445956 162694 446002 162754
rect 448237 162752 448284 162756
rect 448348 162754 448354 162756
rect 448237 162696 448242 162752
rect 445956 162692 445962 162694
rect 448237 162692 448284 162696
rect 448348 162694 448394 162754
rect 453389 162752 453436 162756
rect 453500 162754 453506 162756
rect 453389 162696 453394 162752
rect 448348 162692 448354 162694
rect 453389 162692 453436 162696
rect 453500 162694 453546 162754
rect 458357 162752 458404 162756
rect 458468 162754 458474 162756
rect 458357 162696 458362 162752
rect 453500 162692 453506 162694
rect 458357 162692 458404 162696
rect 458468 162694 458514 162754
rect 458468 162692 458474 162694
rect 503110 162692 503116 162756
rect 503180 162754 503186 162756
rect 503253 162754 503319 162757
rect 503180 162752 503319 162754
rect 503180 162696 503258 162752
rect 503314 162696 503319 162752
rect 503180 162694 503319 162696
rect 503180 162692 503186 162694
rect 440877 162691 440943 162692
rect 443453 162691 443519 162692
rect 445845 162691 445911 162692
rect 448237 162691 448303 162692
rect 453389 162691 453455 162692
rect 458357 162691 458423 162692
rect 503253 162691 503319 162694
rect 50705 162618 50771 162621
rect 183185 162620 183251 162621
rect 158478 162618 158484 162620
rect 50705 162616 158484 162618
rect 50705 162560 50710 162616
rect 50766 162560 158484 162616
rect 50705 162558 158484 162560
rect 50705 162555 50771 162558
rect 158478 162556 158484 162558
rect 158548 162556 158554 162620
rect 183134 162618 183140 162620
rect 183094 162558 183140 162618
rect 183204 162616 183251 162620
rect 183246 162560 183251 162616
rect 183134 162556 183140 162558
rect 183204 162556 183251 162560
rect 207974 162556 207980 162620
rect 208044 162618 208050 162620
rect 323342 162618 323348 162620
rect 208044 162558 323348 162618
rect 208044 162556 208050 162558
rect 323342 162556 323348 162558
rect 323412 162556 323418 162620
rect 343214 162556 343220 162620
rect 343284 162618 343290 162620
rect 343357 162618 343423 162621
rect 343284 162616 343423 162618
rect 343284 162560 343362 162616
rect 343418 162560 343423 162616
rect 343284 162558 343423 162560
rect 343284 162556 343290 162558
rect 183185 162555 183251 162556
rect 343357 162555 343423 162558
rect 379053 162618 379119 162621
rect 468518 162618 468524 162620
rect 379053 162616 468524 162618
rect 379053 162560 379058 162616
rect 379114 162560 468524 162616
rect 379053 162558 468524 162560
rect 379053 162555 379119 162558
rect 468518 162556 468524 162558
rect 468588 162556 468594 162620
rect 503478 162556 503484 162620
rect 503548 162618 503554 162620
rect 503621 162618 503687 162621
rect 503548 162616 503687 162618
rect 503548 162560 503626 162616
rect 503682 162560 503687 162616
rect 503548 162558 503687 162560
rect 503548 162556 503554 162558
rect 503621 162555 503687 162558
rect 47894 162420 47900 162484
rect 47964 162482 47970 162484
rect 90909 162482 90975 162485
rect 47964 162480 90975 162482
rect 47964 162424 90914 162480
rect 90970 162424 90975 162480
rect 47964 162422 90975 162424
rect 47964 162420 47970 162422
rect 90909 162419 90975 162422
rect 91093 162482 91159 162485
rect 91502 162482 91508 162484
rect 91093 162480 91508 162482
rect 91093 162424 91098 162480
rect 91154 162424 91508 162480
rect 91093 162422 91508 162424
rect 91093 162419 91159 162422
rect 91502 162420 91508 162422
rect 91572 162420 91578 162484
rect 106365 162482 106431 162485
rect 116025 162484 116091 162485
rect 107510 162482 107516 162484
rect 106365 162480 107516 162482
rect 106365 162424 106370 162480
rect 106426 162424 107516 162480
rect 106365 162422 107516 162424
rect 106365 162419 106431 162422
rect 107510 162420 107516 162422
rect 107580 162420 107586 162484
rect 115974 162482 115980 162484
rect 115934 162422 115980 162482
rect 116044 162480 116091 162484
rect 116086 162424 116091 162480
rect 115974 162420 115980 162422
rect 116044 162420 116091 162424
rect 203190 162420 203196 162484
rect 203260 162482 203266 162484
rect 311014 162482 311020 162484
rect 203260 162422 311020 162482
rect 203260 162420 203266 162422
rect 311014 162420 311020 162422
rect 311084 162420 311090 162484
rect 376109 162482 376175 162485
rect 462630 162482 462636 162484
rect 376109 162480 462636 162482
rect 376109 162424 376114 162480
rect 376170 162424 462636 162480
rect 376109 162422 462636 162424
rect 116025 162419 116091 162420
rect 376109 162419 376175 162422
rect 462630 162420 462636 162422
rect 462700 162420 462706 162484
rect 47710 162284 47716 162348
rect 47780 162346 47786 162348
rect 160870 162346 160876 162348
rect 47780 162286 160876 162346
rect 47780 162284 47786 162286
rect 160870 162284 160876 162286
rect 160940 162284 160946 162348
rect 213310 162284 213316 162348
rect 213380 162346 213386 162348
rect 315062 162346 315068 162348
rect 213380 162286 315068 162346
rect 213380 162284 213386 162286
rect 315062 162284 315068 162286
rect 315132 162284 315138 162348
rect 378869 162346 378935 162349
rect 460974 162346 460980 162348
rect 378869 162344 460980 162346
rect 378869 162288 378874 162344
rect 378930 162288 460980 162344
rect 378869 162286 460980 162288
rect 378869 162283 378935 162286
rect 460974 162284 460980 162286
rect 461044 162284 461050 162348
rect 75913 162210 75979 162213
rect 88333 162212 88399 162213
rect 77150 162210 77156 162212
rect 75913 162208 77156 162210
rect 75913 162152 75918 162208
rect 75974 162152 77156 162208
rect 75913 162150 77156 162152
rect 75913 162147 75979 162150
rect 77150 162148 77156 162150
rect 77220 162148 77226 162212
rect 88333 162208 88380 162212
rect 88444 162210 88450 162212
rect 90909 162210 90975 162213
rect 93710 162210 93716 162212
rect 88333 162152 88338 162208
rect 88333 162148 88380 162152
rect 88444 162150 88490 162210
rect 90909 162208 93716 162210
rect 90909 162152 90914 162208
rect 90970 162152 93716 162208
rect 90909 162150 93716 162152
rect 88444 162148 88450 162150
rect 88333 162147 88399 162148
rect 90909 162147 90975 162150
rect 93710 162148 93716 162150
rect 93780 162148 93786 162212
rect 112294 162148 112300 162212
rect 112364 162210 112370 162212
rect 112805 162210 112871 162213
rect 112364 162208 112871 162210
rect 112364 162152 112810 162208
rect 112866 162152 112871 162208
rect 112364 162150 112871 162152
rect 112364 162148 112370 162150
rect 112805 162147 112871 162150
rect 215886 162148 215892 162212
rect 215956 162210 215962 162212
rect 278446 162210 278452 162212
rect 215956 162150 278452 162210
rect 215956 162148 215962 162150
rect 278446 162148 278452 162150
rect 278516 162148 278522 162212
rect 396165 162210 396231 162213
rect 397126 162210 397132 162212
rect 396165 162208 397132 162210
rect 396165 162152 396170 162208
rect 396226 162152 397132 162208
rect 396165 162150 397132 162152
rect 396165 162147 396231 162150
rect 397126 162148 397132 162150
rect 397196 162148 397202 162212
rect 402973 162210 403039 162213
rect 404118 162210 404124 162212
rect 402973 162208 404124 162210
rect 402973 162152 402978 162208
rect 403034 162152 404124 162208
rect 402973 162150 404124 162152
rect 402973 162147 403039 162150
rect 404118 162148 404124 162150
rect 404188 162148 404194 162212
rect 411253 162210 411319 162213
rect 412398 162210 412404 162212
rect 411253 162208 412404 162210
rect 411253 162152 411258 162208
rect 411314 162152 412404 162208
rect 411253 162150 412404 162152
rect 411253 162147 411319 162150
rect 412398 162148 412404 162150
rect 412468 162148 412474 162212
rect 418102 162148 418108 162212
rect 418172 162210 418178 162212
rect 418245 162210 418311 162213
rect 418172 162208 418311 162210
rect 418172 162152 418250 162208
rect 418306 162152 418311 162208
rect 418172 162150 418311 162152
rect 418172 162148 418178 162150
rect 418245 162147 418311 162150
rect 426525 162210 426591 162213
rect 427670 162210 427676 162212
rect 426525 162208 427676 162210
rect 426525 162152 426530 162208
rect 426586 162152 427676 162208
rect 426525 162150 427676 162152
rect 426525 162147 426591 162150
rect 427670 162148 427676 162150
rect 427740 162148 427746 162212
rect 433374 162148 433380 162212
rect 433444 162210 433450 162212
rect 434621 162210 434687 162213
rect 433444 162208 434687 162210
rect 433444 162152 434626 162208
rect 434682 162152 434687 162208
rect 433444 162150 434687 162152
rect 433444 162148 433450 162150
rect 434621 162147 434687 162150
rect 100753 162074 100819 162077
rect 101806 162074 101812 162076
rect 100753 162072 101812 162074
rect 100753 162016 100758 162072
rect 100814 162016 101812 162072
rect 100753 162014 101812 162016
rect 100753 162011 100819 162014
rect 101806 162012 101812 162014
rect 101876 162012 101882 162076
rect 244273 162074 244339 162077
rect 245326 162074 245332 162076
rect 244273 162072 245332 162074
rect 244273 162016 244278 162072
rect 244334 162016 245332 162072
rect 244273 162014 245332 162016
rect 244273 162011 244339 162014
rect 245326 162012 245332 162014
rect 245396 162012 245402 162076
rect 251265 162074 251331 162077
rect 252318 162074 252324 162076
rect 251265 162072 252324 162074
rect 251265 162016 251270 162072
rect 251326 162016 252324 162072
rect 251265 162014 252324 162016
rect 251265 162011 251331 162014
rect 252318 162012 252324 162014
rect 252388 162012 252394 162076
rect 259545 162074 259611 162077
rect 260598 162074 260604 162076
rect 259545 162072 260604 162074
rect 259545 162016 259550 162072
rect 259606 162016 260604 162072
rect 259545 162014 260604 162016
rect 259545 162011 259611 162014
rect 260598 162012 260604 162014
rect 260668 162012 260674 162076
rect 273294 162012 273300 162076
rect 273364 162074 273370 162076
rect 274541 162074 274607 162077
rect 273364 162072 274607 162074
rect 273364 162016 274546 162072
rect 274602 162016 274607 162072
rect 273364 162014 274607 162016
rect 273364 162012 273370 162014
rect 274541 162011 274607 162014
rect 393957 162074 394023 162077
rect 415301 162074 415367 162077
rect 393957 162072 415367 162074
rect 393957 162016 393962 162072
rect 394018 162016 415306 162072
rect 415362 162016 415367 162072
rect 393957 162014 415367 162016
rect 393957 162011 394023 162014
rect 415301 162011 415367 162014
rect 433517 162076 433583 162077
rect 433517 162072 433564 162076
rect 433628 162074 433634 162076
rect 433517 162016 433522 162072
rect 433517 162012 433564 162016
rect 433628 162014 433674 162074
rect 433628 162012 433634 162014
rect 433517 162011 433583 162012
rect 206318 161740 206324 161804
rect 206388 161802 206394 161804
rect 326654 161802 326660 161804
rect 206388 161742 326660 161802
rect 206388 161740 206394 161742
rect 326654 161740 326660 161742
rect 326724 161740 326730 161804
rect 376293 161802 376359 161805
rect 465942 161802 465948 161804
rect 376293 161800 465948 161802
rect 376293 161744 376298 161800
rect 376354 161744 465948 161800
rect 376293 161742 465948 161744
rect 376293 161739 376359 161742
rect 465942 161740 465948 161742
rect 466012 161740 466018 161804
rect 84101 161666 84167 161669
rect 84285 161666 84351 161669
rect 84101 161664 84351 161666
rect 84101 161608 84106 161664
rect 84162 161608 84290 161664
rect 84346 161608 84351 161664
rect 84101 161606 84351 161608
rect 84101 161603 84167 161606
rect 84285 161603 84351 161606
rect 238753 161532 238819 161533
rect 238702 161468 238708 161532
rect 238772 161530 238819 161532
rect 258073 161530 258139 161533
rect 258390 161530 258396 161532
rect 238772 161528 238864 161530
rect 238814 161472 238864 161528
rect 238772 161470 238864 161472
rect 258073 161528 258396 161530
rect 258073 161472 258078 161528
rect 258134 161472 258396 161528
rect 258073 161470 258396 161472
rect 238772 161468 238819 161470
rect 238753 161467 238819 161468
rect 258073 161467 258139 161470
rect 258390 161468 258396 161470
rect 258460 161468 258466 161532
rect 277342 161468 277348 161532
rect 277412 161530 277418 161532
rect 278037 161530 278103 161533
rect 277412 161528 278103 161530
rect 277412 161472 278042 161528
rect 278098 161472 278103 161528
rect 277412 161470 278103 161472
rect 277412 161468 277418 161470
rect 278037 161467 278103 161470
rect 412541 161530 412607 161533
rect 412725 161530 412791 161533
rect 412541 161528 412791 161530
rect 412541 161472 412546 161528
rect 412602 161472 412730 161528
rect 412786 161472 412791 161528
rect 412541 161470 412791 161472
rect 412541 161467 412607 161470
rect 412725 161467 412791 161470
rect 217542 161060 217548 161124
rect 217612 161122 217618 161124
rect 217869 161122 217935 161125
rect 217612 161120 217935 161122
rect 217612 161064 217874 161120
rect 217930 161064 217935 161120
rect 217612 161062 217935 161064
rect 217612 161060 217618 161062
rect 217869 161059 217935 161062
rect 56869 160170 56935 160173
rect 57830 160170 57836 160172
rect 56869 160168 57836 160170
rect 56869 160112 56874 160168
rect 56930 160112 57836 160168
rect 56869 160110 57836 160112
rect 56869 160107 56935 160110
rect 57830 160108 57836 160110
rect 57900 160108 57906 160172
rect 580257 152690 580323 152693
rect 583520 152690 584960 152780
rect 580257 152688 584960 152690
rect 580257 152632 580262 152688
rect 580318 152632 584960 152688
rect 580257 152630 584960 152632
rect 580257 152627 580323 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect -960 149774 674 149834
rect -960 149698 480 149774
rect 614 149698 674 149774
rect -960 149684 674 149698
rect 246 149638 674 149684
rect 246 149154 306 149638
rect 360878 149154 360884 149156
rect 246 149094 360884 149154
rect 360878 149092 360884 149094
rect 360948 149092 360954 149156
rect 278221 149018 278287 149021
rect 357709 149018 357775 149021
rect 278221 149016 357775 149018
rect 278221 148960 278226 149016
rect 278282 148960 357714 149016
rect 357770 148960 357775 149016
rect 278221 148958 357775 148960
rect 278221 148955 278287 148958
rect 357709 148955 357775 148958
rect 370957 148474 371023 148477
rect 379462 148474 379468 148476
rect 370957 148472 379468 148474
rect 370957 148416 370962 148472
rect 371018 148416 379468 148472
rect 370957 148414 379468 148416
rect 370957 148411 371023 148414
rect 379462 148412 379468 148414
rect 379532 148474 379538 148476
rect 380801 148474 380867 148477
rect 379532 148472 380867 148474
rect 379532 148416 380806 148472
rect 380862 148416 380867 148472
rect 379532 148414 380867 148416
rect 379532 148412 379538 148414
rect 380801 148411 380867 148414
rect 217358 148276 217364 148340
rect 217428 148338 217434 148340
rect 278221 148338 278287 148341
rect 217428 148336 278287 148338
rect 217428 148280 278226 148336
rect 278282 148280 278287 148336
rect 217428 148278 278287 148280
rect 217428 148276 217434 148278
rect 278221 148275 278287 148278
rect 377622 148276 377628 148340
rect 377692 148338 377698 148340
rect 438853 148338 438919 148341
rect 377692 148336 438919 148338
rect 377692 148280 438858 148336
rect 438914 148280 438919 148336
rect 377692 148278 438919 148280
rect 377692 148276 377698 148278
rect 438853 148275 438919 148278
rect 57053 147522 57119 147525
rect 57278 147522 57284 147524
rect 57053 147520 57284 147522
rect 57053 147464 57058 147520
rect 57114 147464 57284 147520
rect 57053 147462 57284 147464
rect 57053 147459 57119 147462
rect 57278 147460 57284 147462
rect 57348 147460 57354 147524
rect 217174 146372 217180 146436
rect 217244 146434 217250 146436
rect 276013 146434 276079 146437
rect 217244 146432 276079 146434
rect 217244 146376 276018 146432
rect 276074 146376 276079 146432
rect 217244 146374 276079 146376
rect 217244 146372 217250 146374
rect 276013 146371 276079 146374
rect 53741 146298 53807 146301
rect 56317 146298 56383 146301
rect 53741 146296 56383 146298
rect 53741 146240 53746 146296
rect 53802 146240 56322 146296
rect 56378 146240 56383 146296
rect 53741 146238 56383 146240
rect 53741 146235 53807 146238
rect 56317 146235 56383 146238
rect 216213 146298 216279 146301
rect 262213 146298 262279 146301
rect 216213 146296 262279 146298
rect 216213 146240 216218 146296
rect 216274 146240 262218 146296
rect 262274 146240 262279 146296
rect 216213 146238 262279 146240
rect 216213 146235 216279 146238
rect 262213 146235 262279 146238
rect 374453 146298 374519 146301
rect 375925 146298 375991 146301
rect 374453 146296 375991 146298
rect 374453 146240 374458 146296
rect 374514 146240 375930 146296
rect 375986 146240 375991 146296
rect 374453 146238 375991 146240
rect 374453 146235 374519 146238
rect 375925 146235 375991 146238
rect 377990 146236 377996 146300
rect 378060 146298 378066 146300
rect 379145 146298 379211 146301
rect 378060 146296 379211 146298
rect 378060 146240 379150 146296
rect 379206 146240 379211 146296
rect 378060 146238 379211 146240
rect 378060 146236 378066 146238
rect 379145 146235 379211 146238
rect 379513 146298 379579 146301
rect 379973 146298 380039 146301
rect 414013 146298 414079 146301
rect 379513 146296 414079 146298
rect 379513 146240 379518 146296
rect 379574 146240 379978 146296
rect 380034 146240 414018 146296
rect 414074 146240 414079 146296
rect 379513 146238 414079 146240
rect 379513 146235 379579 146238
rect 379973 146235 380039 146238
rect 414013 146235 414079 146238
rect 58617 146026 58683 146029
rect 92473 146026 92539 146029
rect 58617 146024 92539 146026
rect 58617 145968 58622 146024
rect 58678 145968 92478 146024
rect 92534 145968 92539 146024
rect 58617 145966 92539 145968
rect 58617 145963 58683 145966
rect 92473 145963 92539 145966
rect 215753 146026 215819 146029
rect 216213 146026 216279 146029
rect 215753 146024 216279 146026
rect 215753 145968 215758 146024
rect 215814 145968 216218 146024
rect 216274 145968 216279 146024
rect 215753 145966 216279 145968
rect 215753 145963 215819 145966
rect 216213 145963 216279 145966
rect 56409 145890 56475 145893
rect 98637 145890 98703 145893
rect 56409 145888 98703 145890
rect 56409 145832 56414 145888
rect 56470 145832 98642 145888
rect 98698 145832 98703 145888
rect 56409 145830 98703 145832
rect 56409 145827 56475 145830
rect 98637 145827 98703 145830
rect 214557 145890 214623 145893
rect 237373 145890 237439 145893
rect 214557 145888 237439 145890
rect 214557 145832 214562 145888
rect 214618 145832 237378 145888
rect 237434 145832 237439 145888
rect 214557 145830 237439 145832
rect 214557 145827 214623 145830
rect 237373 145827 237439 145830
rect 379145 145890 379211 145893
rect 415485 145890 415551 145893
rect 379145 145888 415551 145890
rect 379145 145832 379150 145888
rect 379206 145832 415490 145888
rect 415546 145832 415551 145888
rect 379145 145830 415551 145832
rect 379145 145827 379211 145830
rect 415485 145827 415551 145830
rect 57646 145692 57652 145756
rect 57716 145754 57722 145756
rect 100017 145754 100083 145757
rect 57716 145752 100083 145754
rect 57716 145696 100022 145752
rect 100078 145696 100083 145752
rect 57716 145694 100083 145696
rect 57716 145692 57722 145694
rect 100017 145691 100083 145694
rect 216305 145754 216371 145757
rect 269113 145754 269179 145757
rect 216305 145752 269179 145754
rect 216305 145696 216310 145752
rect 216366 145696 269118 145752
rect 269174 145696 269179 145752
rect 216305 145694 269179 145696
rect 216305 145691 216371 145694
rect 269113 145691 269179 145694
rect 375925 145754 375991 145757
rect 416773 145754 416839 145757
rect 375925 145752 416839 145754
rect 375925 145696 375930 145752
rect 375986 145696 416778 145752
rect 416834 145696 416839 145752
rect 375925 145694 416839 145696
rect 375925 145691 375991 145694
rect 416773 145691 416839 145694
rect 56041 145618 56107 145621
rect 56317 145618 56383 145621
rect 100753 145618 100819 145621
rect 270493 145618 270559 145621
rect 56041 145616 100819 145618
rect 56041 145560 56046 145616
rect 56102 145560 56322 145616
rect 56378 145560 100758 145616
rect 100814 145560 100819 145616
rect 56041 145558 100819 145560
rect 56041 145555 56107 145558
rect 56317 145555 56383 145558
rect 100753 145555 100819 145558
rect 215250 145616 270559 145618
rect 215250 145560 270498 145616
rect 270554 145560 270559 145616
rect 215250 145558 270559 145560
rect 190862 145420 190868 145484
rect 190932 145482 190938 145484
rect 191741 145482 191807 145485
rect 190932 145480 191807 145482
rect 190932 145424 191746 145480
rect 191802 145424 191807 145480
rect 190932 145422 191807 145424
rect 190932 145420 190938 145422
rect 191741 145419 191807 145422
rect 215017 145482 215083 145485
rect 215250 145482 215310 145558
rect 270493 145555 270559 145558
rect 372521 145618 372587 145621
rect 377806 145618 377812 145620
rect 372521 145616 377812 145618
rect 372521 145560 372526 145616
rect 372582 145560 377812 145616
rect 372521 145558 377812 145560
rect 372521 145555 372587 145558
rect 377806 145556 377812 145558
rect 377876 145618 377882 145620
rect 422293 145618 422359 145621
rect 377876 145616 422359 145618
rect 377876 145560 422298 145616
rect 422354 145560 422359 145616
rect 377876 145558 422359 145560
rect 377876 145556 377882 145558
rect 422293 145555 422359 145558
rect 215017 145480 215310 145482
rect 215017 145424 215022 145480
rect 215078 145424 215310 145480
rect 215017 145422 215310 145424
rect 510613 145482 510679 145485
rect 510838 145482 510844 145484
rect 510613 145480 510844 145482
rect 510613 145424 510618 145480
rect 510674 145424 510844 145480
rect 510613 145422 510844 145424
rect 215017 145419 215083 145422
rect 510613 145419 510679 145422
rect 510838 145420 510844 145422
rect 510908 145420 510914 145484
rect 178534 144876 178540 144940
rect 178604 144938 178610 144940
rect 179045 144938 179111 144941
rect 179689 144940 179755 144941
rect 338481 144940 338547 144941
rect 179638 144938 179644 144940
rect 178604 144936 179111 144938
rect 178604 144880 179050 144936
rect 179106 144880 179111 144936
rect 178604 144878 179111 144880
rect 179598 144878 179644 144938
rect 179708 144936 179755 144940
rect 338430 144938 338436 144940
rect 179750 144880 179755 144936
rect 178604 144876 178610 144878
rect 179045 144875 179111 144878
rect 179638 144876 179644 144878
rect 179708 144876 179755 144880
rect 338390 144878 338436 144938
rect 338500 144936 338547 144940
rect 338542 144880 338547 144936
rect 338430 144876 338436 144878
rect 338500 144876 338547 144880
rect 339718 144876 339724 144940
rect 339788 144938 339794 144940
rect 340229 144938 340295 144941
rect 339788 144936 340295 144938
rect 339788 144880 340234 144936
rect 340290 144880 340295 144936
rect 339788 144878 340295 144880
rect 339788 144876 339794 144878
rect 179689 144875 179755 144876
rect 338481 144875 338547 144876
rect 340229 144875 340295 144878
rect 350942 144876 350948 144940
rect 351012 144938 351018 144940
rect 351637 144938 351703 144941
rect 351012 144936 351703 144938
rect 351012 144880 351642 144936
rect 351698 144880 351703 144936
rect 351012 144878 351703 144880
rect 351012 144876 351018 144878
rect 351637 144875 351703 144878
rect 498510 144876 498516 144940
rect 498580 144938 498586 144940
rect 498653 144938 498719 144941
rect 498580 144936 498719 144938
rect 498580 144880 498658 144936
rect 498714 144880 498719 144936
rect 498580 144878 498719 144880
rect 498580 144876 498586 144878
rect 498653 144875 498719 144878
rect 499798 144876 499804 144940
rect 499868 144938 499874 144940
rect 500217 144938 500283 144941
rect 499868 144936 500283 144938
rect 499868 144880 500222 144936
rect 500278 144880 500283 144936
rect 499868 144878 500283 144880
rect 499868 144876 499874 144878
rect 500217 144875 500283 144878
rect 51533 144802 51599 144805
rect 57094 144802 57100 144804
rect 51533 144800 57100 144802
rect 51533 144744 51538 144800
rect 51594 144744 57100 144800
rect 51533 144742 57100 144744
rect 51533 144739 51599 144742
rect 57094 144740 57100 144742
rect 57164 144802 57170 144804
rect 57646 144802 57652 144804
rect 57164 144742 57652 144802
rect 57164 144740 57170 144742
rect 57646 144740 57652 144742
rect 57716 144740 57722 144804
rect 57462 140796 57468 140860
rect 57532 140858 57538 140860
rect 59353 140858 59419 140861
rect 57532 140856 59419 140858
rect 57532 140800 59358 140856
rect 59414 140800 59419 140856
rect 57532 140798 59419 140800
rect 57532 140796 57538 140798
rect 59353 140795 59419 140798
rect 359365 139362 359431 139365
rect 519353 139362 519419 139365
rect 356562 139360 359431 139362
rect 356562 139304 359370 139360
rect 359426 139304 359431 139360
rect 356562 139302 359431 139304
rect 199193 139226 199259 139229
rect 197126 139224 199259 139226
rect 197126 139220 199198 139224
rect 196604 139168 199198 139220
rect 199254 139168 199259 139224
rect 356562 139190 356622 139302
rect 359365 139299 359431 139302
rect 516558 139360 519419 139362
rect 516558 139304 519358 139360
rect 519414 139304 519419 139360
rect 516558 139302 519419 139304
rect 516558 139190 516618 139302
rect 519353 139299 519419 139302
rect 583520 139212 584960 139452
rect 196604 139166 199259 139168
rect 196604 139160 197186 139166
rect 199193 139163 199259 139166
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 580441 112842 580507 112845
rect 583520 112842 584960 112932
rect 580441 112840 584960 112842
rect 580441 112784 580446 112840
rect 580502 112784 584960 112840
rect 580441 112782 584960 112784
rect 580441 112779 580507 112782
rect 583520 112692 584960 112782
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97610 480 97700
rect 3509 97610 3575 97613
rect -960 97608 3575 97610
rect -960 97552 3514 97608
rect 3570 97552 3575 97608
rect -960 97550 3575 97552
rect -960 97460 480 97550
rect 3509 97547 3575 97550
rect 57237 97474 57303 97477
rect 57237 97472 60062 97474
rect 57237 97416 57242 97472
rect 57298 97416 60062 97472
rect 57237 97414 60062 97416
rect 57237 97411 57303 97414
rect 60002 96894 60062 97414
rect 216673 96930 216739 96933
rect 377581 96930 377647 96933
rect 216673 96928 219450 96930
rect 216673 96872 216678 96928
rect 216734 96924 219450 96928
rect 377581 96928 379530 96930
rect 216734 96872 220064 96924
rect 216673 96870 220064 96872
rect 216673 96867 216739 96870
rect 219390 96864 220064 96870
rect 377581 96872 377586 96928
rect 377642 96924 379530 96928
rect 377642 96872 380052 96924
rect 377581 96870 380052 96872
rect 377581 96867 377647 96870
rect 379470 96864 380052 96870
rect 57145 96522 57211 96525
rect 57145 96520 60062 96522
rect 57145 96464 57150 96520
rect 57206 96464 60062 96520
rect 57145 96462 60062 96464
rect 57145 96459 57211 96462
rect 60002 95942 60062 96462
rect 216765 95978 216831 95981
rect 377305 95978 377371 95981
rect 216765 95976 219450 95978
rect 216765 95920 216770 95976
rect 216826 95972 219450 95976
rect 377305 95976 379530 95978
rect 216826 95920 220064 95972
rect 216765 95918 220064 95920
rect 216765 95915 216831 95918
rect 219390 95912 220064 95918
rect 377305 95920 377310 95976
rect 377366 95972 379530 95976
rect 377366 95920 380052 95972
rect 377305 95918 380052 95920
rect 377305 95915 377371 95918
rect 379470 95912 380052 95918
rect 57605 93802 57671 93805
rect 217777 93802 217843 93805
rect 376937 93802 377003 93805
rect 57605 93800 60062 93802
rect 57605 93744 57610 93800
rect 57666 93744 60062 93800
rect 57605 93742 60062 93744
rect 217777 93800 219450 93802
rect 217777 93744 217782 93800
rect 217838 93796 219450 93800
rect 376937 93800 379530 93802
rect 217838 93744 220064 93796
rect 217777 93742 220064 93744
rect 57605 93739 57671 93742
rect 217777 93739 217843 93742
rect 219390 93736 220064 93742
rect 376937 93744 376942 93800
rect 376998 93796 379530 93800
rect 376998 93744 380052 93796
rect 376937 93742 380052 93744
rect 376937 93739 377003 93742
rect 379470 93736 380052 93742
rect 57329 93394 57395 93397
rect 57329 93392 60062 93394
rect 57329 93336 57334 93392
rect 57390 93336 60062 93392
rect 57329 93334 60062 93336
rect 57329 93331 57395 93334
rect 60002 92814 60062 93334
rect 216857 92850 216923 92853
rect 377489 92850 377555 92853
rect 216857 92848 219450 92850
rect 216857 92792 216862 92848
rect 216918 92844 219450 92848
rect 377489 92848 379530 92850
rect 216918 92792 220064 92844
rect 216857 92790 220064 92792
rect 216857 92787 216923 92790
rect 219390 92784 220064 92790
rect 377489 92792 377494 92848
rect 377550 92844 379530 92848
rect 377550 92792 380052 92844
rect 377489 92790 380052 92792
rect 377489 92787 377555 92790
rect 379470 92784 380052 92790
rect 57697 91082 57763 91085
rect 217685 91082 217751 91085
rect 377029 91082 377095 91085
rect 57697 91080 60062 91082
rect 57697 91024 57702 91080
rect 57758 91024 60062 91080
rect 57697 91022 60062 91024
rect 217685 91080 219450 91082
rect 217685 91024 217690 91080
rect 217746 91076 219450 91080
rect 377029 91080 379530 91082
rect 217746 91024 220064 91076
rect 217685 91022 220064 91024
rect 57697 91019 57763 91022
rect 217685 91019 217751 91022
rect 219390 91016 220064 91022
rect 377029 91024 377034 91080
rect 377090 91076 379530 91080
rect 377090 91024 380052 91076
rect 377029 91022 380052 91024
rect 377029 91019 377095 91022
rect 379470 91016 380052 91022
rect 57421 90538 57487 90541
rect 57421 90536 60062 90538
rect 57421 90480 57426 90536
rect 57482 90480 60062 90536
rect 57421 90478 60062 90480
rect 57421 90475 57487 90478
rect 60002 89958 60062 90478
rect 217225 89994 217291 89997
rect 377765 89994 377831 89997
rect 217225 89992 219450 89994
rect 217225 89936 217230 89992
rect 217286 89988 219450 89992
rect 377765 89992 379530 89994
rect 217286 89936 220064 89988
rect 217225 89934 220064 89936
rect 217225 89931 217291 89934
rect 219390 89928 220064 89934
rect 377765 89936 377770 89992
rect 377826 89988 379530 89992
rect 377826 89936 380052 89988
rect 377765 89934 380052 89936
rect 377765 89931 377831 89934
rect 379470 89928 380052 89934
rect 57513 88226 57579 88229
rect 217593 88226 217659 88229
rect 377213 88226 377279 88229
rect 57513 88224 60062 88226
rect 57513 88168 57518 88224
rect 57574 88168 60062 88224
rect 57513 88166 60062 88168
rect 217593 88224 219450 88226
rect 217593 88168 217598 88224
rect 217654 88220 219450 88224
rect 377213 88224 379530 88226
rect 217654 88168 220064 88220
rect 217593 88166 220064 88168
rect 57513 88163 57579 88166
rect 217593 88163 217659 88166
rect 219390 88160 220064 88166
rect 377213 88168 377218 88224
rect 377274 88220 379530 88224
rect 377274 88168 380052 88220
rect 377213 88166 380052 88168
rect 377213 88163 377279 88166
rect 379470 88160 380052 88166
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 359089 79930 359155 79933
rect 519261 79930 519327 79933
rect 520181 79930 520247 79933
rect 356562 79928 359155 79930
rect 356562 79872 359094 79928
rect 359150 79872 359155 79928
rect 356562 79870 359155 79872
rect 199009 79386 199075 79389
rect 197126 79384 199075 79386
rect 197126 79380 199014 79384
rect 196604 79328 199014 79380
rect 199070 79328 199075 79384
rect 356562 79350 356622 79870
rect 359089 79867 359155 79870
rect 516558 79928 520247 79930
rect 516558 79872 519266 79928
rect 519322 79872 520186 79928
rect 520242 79872 520247 79928
rect 516558 79870 520247 79872
rect 516558 79350 516618 79870
rect 519261 79867 519327 79870
rect 520181 79867 520247 79870
rect 196604 79326 199075 79328
rect 196604 79320 197186 79326
rect 199009 79323 199075 79326
rect 358905 78298 358971 78301
rect 519169 78298 519235 78301
rect 356562 78296 358971 78298
rect 356562 78240 358910 78296
rect 358966 78240 358971 78296
rect 356562 78238 358971 78240
rect 199377 77754 199443 77757
rect 197126 77752 199443 77754
rect 197126 77748 199382 77752
rect 196604 77696 199382 77748
rect 199438 77696 199443 77752
rect 356562 77718 356622 78238
rect 358905 78235 358971 78238
rect 516558 78296 519235 78298
rect 516558 78240 519174 78296
rect 519230 78240 519235 78296
rect 516558 78238 519235 78240
rect 516558 77718 516618 78238
rect 519169 78235 519235 78238
rect 196604 77694 199443 77696
rect 196604 77688 197186 77694
rect 199377 77691 199443 77694
rect 359181 76938 359247 76941
rect 356562 76936 359247 76938
rect 356562 76880 359186 76936
rect 359242 76880 359247 76936
rect 356562 76878 359247 76880
rect 198825 76394 198891 76397
rect 197126 76392 198891 76394
rect 197126 76388 198830 76392
rect 196604 76336 198830 76388
rect 198886 76336 198891 76392
rect 356562 76358 356622 76878
rect 359181 76875 359247 76878
rect 519537 76802 519603 76805
rect 516558 76800 519603 76802
rect 516558 76744 519542 76800
rect 519598 76744 519603 76800
rect 516558 76742 519603 76744
rect 516558 76358 516618 76742
rect 519537 76739 519603 76742
rect 196604 76334 198891 76336
rect 196604 76328 197186 76334
rect 198825 76331 198891 76334
rect 359273 75442 359339 75445
rect 518985 75442 519051 75445
rect 356562 75440 359339 75442
rect 356562 75384 359278 75440
rect 359334 75384 359339 75440
rect 356562 75382 359339 75384
rect 198733 74898 198799 74901
rect 197126 74896 198799 74898
rect 197126 74892 198738 74896
rect 196604 74840 198738 74892
rect 198794 74840 198799 74896
rect 356562 74862 356622 75382
rect 359273 75379 359339 75382
rect 516558 75440 519051 75442
rect 516558 75384 518990 75440
rect 519046 75384 519051 75440
rect 516558 75382 519051 75384
rect 516558 74862 516618 75382
rect 518985 75379 519051 75382
rect 196604 74838 198799 74840
rect 196604 74832 197186 74838
rect 198733 74835 198799 74838
rect 518893 74218 518959 74221
rect 516558 74216 518959 74218
rect 516558 74160 518898 74216
rect 518954 74160 518959 74216
rect 516558 74158 518959 74160
rect 358997 74082 359063 74085
rect 356562 74080 359063 74082
rect 356562 74024 359002 74080
rect 359058 74024 359063 74080
rect 356562 74022 359063 74024
rect 198917 73674 198983 73677
rect 197126 73672 198983 73674
rect 197126 73668 198922 73672
rect 196604 73616 198922 73668
rect 198978 73616 198983 73672
rect 356562 73638 356622 74022
rect 358997 74019 359063 74022
rect 516558 73638 516618 74158
rect 518893 74155 518959 74158
rect 196604 73614 198983 73616
rect 196604 73608 197186 73614
rect 198917 73611 198983 73614
rect 580349 72994 580415 72997
rect 583520 72994 584960 73084
rect 580349 72992 584960 72994
rect 580349 72936 580354 72992
rect 580410 72936 584960 72992
rect 580349 72934 584960 72936
rect 580349 72931 580415 72934
rect 583520 72844 584960 72934
rect -960 71484 480 71724
rect 216673 70002 216739 70005
rect 376937 70002 377003 70005
rect 216673 70000 219450 70002
rect 46790 68988 46796 69052
rect 46860 69050 46866 69052
rect 60002 69050 60062 69966
rect 216673 69944 216678 70000
rect 216734 69996 219450 70000
rect 376937 70000 379530 70002
rect 216734 69944 220064 69996
rect 216673 69942 220064 69944
rect 216673 69939 216739 69942
rect 219390 69936 220064 69942
rect 376937 69944 376942 70000
rect 376998 69996 379530 70000
rect 376998 69944 380052 69996
rect 376937 69942 380052 69944
rect 376937 69939 377003 69942
rect 379470 69936 380052 69942
rect 46860 68990 60062 69050
rect 46860 68988 46866 68990
rect 57881 68914 57947 68917
rect 57881 68912 60062 68914
rect 57881 68856 57886 68912
rect 57942 68856 60062 68912
rect 57881 68854 60062 68856
rect 57881 68851 57947 68854
rect 60002 68334 60062 68854
rect 216673 68370 216739 68373
rect 217961 68370 218027 68373
rect 376937 68370 377003 68373
rect 216673 68368 219450 68370
rect 216673 68312 216678 68368
rect 216734 68312 217966 68368
rect 218022 68364 219450 68368
rect 376937 68368 379530 68370
rect 218022 68312 220064 68364
rect 216673 68310 220064 68312
rect 216673 68307 216739 68310
rect 217961 68307 218027 68310
rect 219390 68304 220064 68310
rect 376937 68312 376942 68368
rect 376998 68364 379530 68368
rect 376998 68312 380052 68364
rect 376937 68310 380052 68312
rect 376937 68307 377003 68310
rect 379470 68304 380052 68310
rect 56869 68098 56935 68101
rect 56869 68096 59554 68098
rect 56869 68040 56874 68096
rect 56930 68092 59554 68096
rect 56930 68040 60032 68092
rect 56869 68038 60032 68040
rect 56869 68035 56935 68038
rect 59494 68032 60032 68038
rect 205030 68036 205036 68100
rect 205100 68098 205106 68100
rect 205100 68092 219450 68098
rect 205100 68038 220064 68092
rect 205100 68036 205106 68038
rect 219390 68032 220064 68038
rect 367870 68036 367876 68100
rect 367940 68098 367946 68100
rect 367940 68092 379530 68098
rect 367940 68038 380052 68092
rect 367940 68036 367946 68038
rect 379470 68032 380052 68038
rect 218697 60620 218763 60621
rect 219249 60620 219315 60621
rect 218646 60618 218652 60620
rect 218606 60558 218652 60618
rect 218716 60616 218763 60620
rect 219198 60618 219204 60620
rect 218758 60560 218763 60616
rect 218646 60556 218652 60558
rect 218716 60556 218763 60560
rect 219158 60558 219204 60618
rect 219268 60616 219315 60620
rect 219310 60560 219315 60616
rect 219198 60556 219204 60558
rect 219268 60556 219315 60560
rect 218697 60555 218763 60556
rect 219249 60555 219315 60556
rect 77109 59804 77175 59805
rect 83089 59804 83155 59805
rect 99465 59804 99531 59805
rect 77109 59800 77142 59804
rect 77206 59802 77212 59804
rect 77109 59744 77114 59800
rect 77109 59740 77142 59744
rect 77206 59742 77266 59802
rect 83089 59800 83126 59804
rect 83190 59802 83196 59804
rect 99440 59802 99446 59804
rect 83089 59744 83094 59800
rect 77206 59740 77212 59742
rect 83089 59740 83126 59744
rect 83190 59742 83246 59802
rect 99374 59742 99446 59802
rect 99510 59800 99531 59804
rect 99526 59744 99531 59800
rect 83190 59740 83196 59742
rect 99440 59740 99446 59742
rect 99510 59740 99531 59744
rect 77109 59739 77175 59740
rect 83089 59739 83155 59740
rect 99465 59739 99531 59740
rect 113541 59804 113607 59805
rect 237097 59804 237163 59805
rect 255865 59804 255931 59805
rect 256969 59804 257035 59805
rect 261753 59804 261819 59805
rect 263869 59804 263935 59805
rect 396073 59804 396139 59805
rect 113541 59800 113590 59804
rect 113654 59802 113660 59804
rect 113541 59744 113546 59800
rect 113541 59740 113590 59744
rect 113654 59742 113698 59802
rect 237097 59800 237142 59804
rect 237206 59802 237212 59804
rect 237097 59744 237102 59800
rect 113654 59740 113660 59742
rect 237097 59740 237142 59744
rect 237206 59742 237254 59802
rect 255865 59800 255910 59804
rect 255974 59802 255980 59804
rect 255865 59744 255870 59800
rect 237206 59740 237212 59742
rect 255865 59740 255910 59744
rect 255974 59742 256022 59802
rect 256969 59800 256998 59804
rect 257062 59802 257068 59804
rect 256969 59744 256974 59800
rect 255974 59740 255980 59742
rect 256969 59740 256998 59744
rect 257062 59742 257126 59802
rect 257062 59740 257068 59742
rect 261752 59740 261758 59804
rect 261822 59802 261828 59804
rect 261822 59742 261910 59802
rect 263869 59800 263934 59804
rect 263869 59744 263874 59800
rect 263930 59744 263934 59800
rect 261822 59740 261828 59742
rect 263869 59740 263934 59744
rect 263998 59802 264004 59804
rect 396048 59802 396054 59804
rect 263998 59742 264026 59802
rect 395982 59742 396054 59802
rect 396118 59800 396139 59804
rect 396134 59744 396139 59800
rect 263998 59740 264004 59742
rect 396048 59740 396054 59742
rect 396118 59740 396139 59744
rect 113541 59739 113607 59740
rect 237097 59739 237163 59740
rect 255865 59739 255931 59740
rect 256969 59739 257035 59740
rect 261753 59739 261819 59740
rect 263869 59739 263935 59740
rect 396073 59739 396139 59740
rect 397085 59804 397151 59805
rect 416957 59804 417023 59805
rect 418429 59804 418495 59805
rect 423949 59804 424015 59805
rect 397085 59800 397142 59804
rect 397206 59802 397212 59804
rect 397085 59744 397090 59800
rect 397085 59740 397142 59744
rect 397206 59742 397242 59802
rect 416957 59800 416998 59804
rect 417062 59802 417068 59804
rect 416957 59744 416962 59800
rect 397206 59740 397212 59742
rect 416957 59740 416998 59744
rect 417062 59742 417114 59802
rect 418429 59800 418494 59804
rect 418429 59744 418434 59800
rect 418490 59744 418494 59800
rect 417062 59740 417068 59742
rect 418429 59740 418494 59744
rect 418558 59802 418564 59804
rect 423928 59802 423934 59804
rect 418558 59742 418586 59802
rect 423858 59742 423934 59802
rect 423998 59800 424015 59804
rect 424010 59744 424015 59800
rect 418558 59740 418564 59742
rect 423928 59740 423934 59742
rect 423998 59740 424015 59744
rect 397085 59739 397151 59740
rect 416957 59739 417023 59740
rect 418429 59739 418495 59740
rect 423949 59739 424015 59740
rect 94497 59668 94563 59669
rect 94497 59664 94550 59668
rect 94614 59666 94620 59668
rect 95693 59666 95759 59669
rect 102777 59668 102843 59669
rect 103881 59668 103947 59669
rect 260649 59668 260715 59669
rect 305913 59668 305979 59669
rect 318425 59668 318491 59669
rect 403065 59668 403131 59669
rect 404169 59668 404235 59669
rect 101072 59666 101078 59668
rect 94497 59608 94502 59664
rect 94497 59604 94550 59608
rect 94614 59606 94654 59666
rect 95693 59664 101078 59666
rect 95693 59608 95698 59664
rect 95754 59608 101078 59664
rect 95693 59606 101078 59608
rect 94614 59604 94620 59606
rect 94497 59603 94563 59604
rect 95693 59603 95759 59606
rect 101072 59604 101078 59606
rect 101142 59604 101148 59668
rect 102777 59664 102846 59668
rect 102777 59608 102782 59664
rect 102838 59608 102846 59664
rect 102777 59604 102846 59608
rect 102910 59666 102916 59668
rect 102910 59606 102934 59666
rect 103881 59664 103934 59668
rect 103998 59666 104004 59668
rect 103881 59608 103886 59664
rect 102910 59604 102916 59606
rect 103881 59604 103934 59608
rect 103998 59606 104038 59666
rect 260649 59664 260670 59668
rect 260734 59666 260740 59668
rect 260649 59608 260654 59664
rect 103998 59604 104004 59606
rect 260649 59604 260670 59608
rect 260734 59606 260806 59666
rect 305913 59664 305958 59668
rect 306022 59666 306028 59668
rect 305913 59608 305918 59664
rect 260734 59604 260740 59606
rect 305913 59604 305958 59608
rect 306022 59606 306070 59666
rect 318425 59664 318470 59668
rect 318534 59666 318540 59668
rect 318425 59608 318430 59664
rect 306022 59604 306028 59606
rect 318425 59604 318470 59608
rect 318534 59606 318582 59666
rect 403065 59664 403126 59668
rect 403065 59608 403070 59664
rect 318534 59604 318540 59606
rect 403065 59604 403126 59608
rect 403190 59666 403196 59668
rect 403190 59606 403222 59666
rect 404169 59664 404214 59668
rect 404278 59666 404284 59668
rect 412541 59666 412607 59669
rect 419441 59668 419507 59669
rect 421741 59668 421807 59669
rect 423489 59668 423555 59669
rect 503253 59668 503319 59669
rect 413456 59666 413462 59668
rect 404169 59608 404174 59664
rect 403190 59604 403196 59606
rect 404169 59604 404214 59608
rect 404278 59606 404326 59666
rect 412541 59664 413462 59666
rect 412541 59608 412546 59664
rect 412602 59608 413462 59664
rect 412541 59606 413462 59608
rect 404278 59604 404284 59606
rect 102777 59603 102843 59604
rect 103881 59603 103947 59604
rect 260649 59603 260715 59604
rect 305913 59603 305979 59604
rect 318425 59603 318491 59604
rect 403065 59603 403131 59604
rect 404169 59603 404235 59604
rect 412541 59603 412607 59606
rect 413456 59604 413462 59606
rect 413526 59604 413532 59668
rect 419440 59604 419446 59668
rect 419510 59666 419516 59668
rect 419510 59606 419598 59666
rect 421741 59664 421758 59668
rect 421822 59666 421828 59668
rect 421741 59608 421746 59664
rect 419510 59604 419516 59606
rect 421741 59604 421758 59608
rect 421822 59606 421898 59666
rect 423489 59664 423526 59668
rect 423590 59666 423596 59668
rect 503216 59666 503222 59668
rect 423489 59608 423494 59664
rect 421822 59604 421828 59606
rect 423489 59604 423526 59608
rect 423590 59606 423646 59666
rect 503162 59606 503222 59666
rect 503286 59664 503319 59668
rect 503314 59608 503319 59664
rect 423590 59604 423596 59606
rect 503216 59604 503222 59606
rect 503286 59604 503319 59608
rect 419441 59603 419507 59604
rect 421741 59603 421807 59604
rect 423489 59603 423555 59604
rect 503253 59603 503319 59604
rect 262765 59532 262831 59533
rect 418153 59532 418219 59533
rect 57094 59468 57100 59532
rect 57164 59530 57170 59532
rect 100702 59530 100708 59532
rect 57164 59470 100708 59530
rect 57164 59468 57170 59470
rect 100702 59468 100708 59470
rect 100772 59468 100778 59532
rect 262765 59528 262812 59532
rect 262876 59530 262882 59532
rect 418102 59530 418108 59532
rect 262765 59472 262770 59528
rect 262765 59468 262812 59472
rect 262876 59470 262922 59530
rect 418062 59470 418108 59530
rect 418172 59528 418219 59532
rect 418214 59472 418219 59528
rect 262876 59468 262882 59470
rect 418102 59468 418108 59470
rect 418172 59468 418219 59472
rect 262765 59467 262831 59468
rect 418153 59467 418219 59468
rect 420637 59532 420703 59533
rect 420637 59528 420684 59532
rect 420748 59530 420754 59532
rect 420637 59472 420642 59528
rect 420637 59468 420684 59472
rect 420748 59470 420794 59530
rect 583520 59516 584960 59756
rect 420748 59468 420754 59470
rect 420637 59467 420703 59468
rect 46606 59332 46612 59396
rect 46676 59394 46682 59396
rect 95693 59394 95759 59397
rect 46676 59392 95759 59394
rect 46676 59336 95698 59392
rect 95754 59336 95759 59392
rect 46676 59334 95759 59336
rect 46676 59332 46682 59334
rect 95693 59331 95759 59334
rect 95877 59396 95943 59397
rect 96981 59396 97047 59397
rect 101765 59396 101831 59397
rect 111149 59396 111215 59397
rect 115933 59396 115999 59397
rect 425237 59396 425303 59397
rect 425973 59396 426039 59397
rect 428181 59396 428247 59397
rect 465901 59396 465967 59397
rect 95877 59392 95924 59396
rect 95988 59394 95994 59396
rect 95877 59336 95882 59392
rect 95877 59332 95924 59336
rect 95988 59334 96034 59394
rect 96981 59392 97028 59396
rect 97092 59394 97098 59396
rect 96981 59336 96986 59392
rect 95988 59332 95994 59334
rect 96981 59332 97028 59336
rect 97092 59334 97138 59394
rect 101765 59392 101812 59396
rect 101876 59394 101882 59396
rect 101765 59336 101770 59392
rect 97092 59332 97098 59334
rect 101765 59332 101812 59336
rect 101876 59334 101922 59394
rect 111149 59392 111196 59396
rect 111260 59394 111266 59396
rect 111149 59336 111154 59392
rect 101876 59332 101882 59334
rect 111149 59332 111196 59336
rect 111260 59334 111306 59394
rect 115933 59392 115980 59396
rect 116044 59394 116050 59396
rect 115933 59336 115938 59392
rect 111260 59332 111266 59334
rect 115933 59332 115980 59336
rect 116044 59334 116090 59394
rect 116044 59332 116050 59334
rect 198038 59332 198044 59396
rect 198108 59394 198114 59396
rect 263542 59394 263548 59396
rect 198108 59334 263548 59394
rect 198108 59332 198114 59334
rect 263542 59332 263548 59334
rect 263612 59332 263618 59396
rect 377806 59332 377812 59396
rect 377876 59394 377882 59396
rect 422886 59394 422892 59396
rect 377876 59334 422892 59394
rect 377876 59332 377882 59334
rect 422886 59332 422892 59334
rect 422956 59332 422962 59396
rect 425237 59392 425284 59396
rect 425348 59394 425354 59396
rect 425237 59336 425242 59392
rect 425237 59332 425284 59336
rect 425348 59334 425394 59394
rect 425973 59392 426020 59396
rect 426084 59394 426090 59396
rect 425973 59336 425978 59392
rect 425348 59332 425354 59334
rect 425973 59332 426020 59336
rect 426084 59334 426130 59394
rect 428181 59392 428228 59396
rect 428292 59394 428298 59396
rect 428181 59336 428186 59392
rect 426084 59332 426090 59334
rect 428181 59332 428228 59336
rect 428292 59334 428338 59394
rect 465901 59392 465948 59396
rect 466012 59394 466018 59396
rect 465901 59336 465906 59392
rect 428292 59332 428298 59334
rect 465901 59332 465948 59336
rect 466012 59334 466058 59394
rect 466012 59332 466018 59334
rect 95877 59331 95943 59332
rect 96981 59331 97047 59332
rect 101765 59331 101831 59332
rect 111149 59331 111215 59332
rect 115933 59331 115999 59332
rect 425237 59331 425303 59332
rect 425973 59331 426039 59332
rect 428181 59331 428247 59332
rect 465901 59331 465967 59332
rect 148501 59260 148567 59261
rect 150893 59260 150959 59261
rect 279233 59260 279299 59261
rect 52310 59196 52316 59260
rect 52380 59258 52386 59260
rect 143574 59258 143580 59260
rect 52380 59198 143580 59258
rect 52380 59196 52386 59198
rect 143574 59196 143580 59198
rect 143644 59196 143650 59260
rect 148501 59256 148548 59260
rect 148612 59258 148618 59260
rect 148501 59200 148506 59256
rect 148501 59196 148548 59200
rect 148612 59198 148658 59258
rect 150893 59256 150940 59260
rect 151004 59258 151010 59260
rect 150893 59200 150898 59256
rect 148612 59196 148618 59198
rect 150893 59196 150940 59200
rect 151004 59198 151050 59258
rect 151004 59196 151010 59198
rect 201350 59196 201356 59260
rect 201420 59258 201426 59260
rect 279182 59258 279188 59260
rect 201420 59198 277410 59258
rect 279142 59198 279188 59258
rect 279252 59256 279299 59260
rect 279294 59200 279299 59256
rect 201420 59196 201426 59198
rect 148501 59195 148567 59196
rect 150893 59195 150959 59196
rect 54702 59060 54708 59124
rect 54772 59122 54778 59124
rect 140814 59122 140820 59124
rect 54772 59062 140820 59122
rect 54772 59060 54778 59062
rect 140814 59060 140820 59062
rect 140884 59060 140890 59124
rect 198590 59060 198596 59124
rect 198660 59122 198666 59124
rect 273478 59122 273484 59124
rect 198660 59062 273484 59122
rect 198660 59060 198666 59062
rect 273478 59060 273484 59062
rect 273548 59060 273554 59124
rect 277350 59122 277410 59198
rect 279182 59196 279188 59198
rect 279252 59196 279299 59200
rect 279233 59195 279299 59196
rect 290917 59260 290983 59261
rect 298461 59260 298527 59261
rect 313365 59260 313431 59261
rect 325877 59260 325943 59261
rect 485957 59260 486023 59261
rect 290917 59256 290964 59260
rect 291028 59258 291034 59260
rect 290917 59200 290922 59256
rect 290917 59196 290964 59200
rect 291028 59198 291074 59258
rect 298461 59256 298508 59260
rect 298572 59258 298578 59260
rect 298461 59200 298466 59256
rect 291028 59196 291034 59198
rect 298461 59196 298508 59200
rect 298572 59198 298618 59258
rect 313365 59256 313412 59260
rect 313476 59258 313482 59260
rect 313365 59200 313370 59256
rect 298572 59196 298578 59198
rect 313365 59196 313412 59200
rect 313476 59198 313522 59258
rect 325877 59256 325924 59260
rect 325988 59258 325994 59260
rect 325877 59200 325882 59256
rect 313476 59196 313482 59198
rect 325877 59196 325924 59200
rect 325988 59198 326034 59258
rect 325988 59196 325994 59198
rect 360694 59196 360700 59260
rect 360764 59258 360770 59260
rect 483422 59258 483428 59260
rect 360764 59198 483428 59258
rect 360764 59196 360770 59198
rect 483422 59196 483428 59198
rect 483492 59196 483498 59260
rect 485957 59256 486004 59260
rect 486068 59258 486074 59260
rect 485957 59200 485962 59256
rect 485957 59196 486004 59200
rect 486068 59198 486114 59258
rect 486068 59196 486074 59198
rect 290917 59195 290983 59196
rect 298461 59195 298527 59196
rect 313365 59195 313431 59196
rect 325877 59195 325943 59196
rect 485957 59195 486023 59196
rect 285990 59122 285996 59124
rect 277350 59062 285996 59122
rect 285990 59060 285996 59062
rect 286060 59060 286066 59124
rect 357934 59060 357940 59124
rect 358004 59122 358010 59124
rect 475878 59122 475884 59124
rect 358004 59062 475884 59122
rect 358004 59060 358010 59062
rect 475878 59060 475884 59062
rect 475948 59060 475954 59124
rect 53414 58924 53420 58988
rect 53484 58986 53490 58988
rect 138422 58986 138428 58988
rect 53484 58926 138428 58986
rect 53484 58924 53490 58926
rect 138422 58924 138428 58926
rect 138492 58924 138498 58988
rect 206870 58924 206876 58988
rect 206940 58986 206946 58988
rect 276054 58986 276060 58988
rect 206940 58926 276060 58986
rect 206940 58924 206946 58926
rect 276054 58924 276060 58926
rect 276124 58924 276130 58988
rect 371734 58924 371740 58988
rect 371804 58986 371810 58988
rect 480846 58986 480852 58988
rect 371804 58926 480852 58986
rect 371804 58924 371810 58926
rect 480846 58924 480852 58926
rect 480916 58924 480922 58988
rect 51942 58788 51948 58852
rect 52012 58850 52018 58852
rect 135846 58850 135852 58852
rect 52012 58790 135852 58850
rect 52012 58788 52018 58790
rect 135846 58788 135852 58790
rect 135916 58788 135922 58852
rect 213678 58788 213684 58852
rect 213748 58850 213754 58852
rect 278446 58850 278452 58852
rect 213748 58790 278452 58850
rect 213748 58788 213754 58790
rect 278446 58788 278452 58790
rect 278516 58788 278522 58852
rect 375966 58788 375972 58852
rect 376036 58850 376042 58852
rect 470910 58850 470916 58852
rect 376036 58790 470916 58850
rect 376036 58788 376042 58790
rect 470910 58788 470916 58790
rect 470980 58788 470986 58852
rect 259453 58716 259519 58717
rect -960 58578 480 58668
rect 59302 58652 59308 58716
rect 59372 58714 59378 58716
rect 120942 58714 120948 58716
rect 59372 58654 120948 58714
rect 59372 58652 59378 58654
rect 120942 58652 120948 58654
rect 121012 58652 121018 58716
rect 197854 58652 197860 58716
rect 197924 58714 197930 58716
rect 253606 58714 253612 58716
rect 197924 58654 253612 58714
rect 197924 58652 197930 58654
rect 253606 58652 253612 58654
rect 253676 58652 253682 58716
rect 259453 58712 259500 58716
rect 259564 58714 259570 58716
rect 259453 58656 259458 58712
rect 259453 58652 259500 58656
rect 259564 58654 259610 58714
rect 259564 58652 259570 58654
rect 370446 58652 370452 58716
rect 370516 58714 370522 58716
rect 458398 58714 458404 58716
rect 370516 58654 458404 58714
rect 370516 58652 370522 58654
rect 458398 58652 458404 58654
rect 458468 58652 458474 58716
rect 259453 58651 259519 58652
rect 3417 58578 3483 58581
rect -960 58576 3483 58578
rect -960 58520 3422 58576
rect 3478 58520 3483 58576
rect -960 58518 3483 58520
rect -960 58428 480 58518
rect 3417 58515 3483 58518
rect 48078 58516 48084 58580
rect 48148 58578 48154 58580
rect 108246 58578 108252 58580
rect 48148 58518 108252 58578
rect 48148 58516 48154 58518
rect 108246 58516 108252 58518
rect 108316 58516 108322 58580
rect 202086 58516 202092 58580
rect 202156 58578 202162 58580
rect 250662 58578 250668 58580
rect 202156 58518 250668 58578
rect 202156 58516 202162 58518
rect 250662 58516 250668 58518
rect 250732 58516 250738 58580
rect 374678 58516 374684 58580
rect 374748 58578 374754 58580
rect 463550 58578 463556 58580
rect 374748 58518 463556 58578
rect 374748 58516 374754 58518
rect 463550 58516 463556 58518
rect 463620 58516 463626 58580
rect 52126 58380 52132 58444
rect 52196 58442 52202 58444
rect 111006 58442 111012 58444
rect 52196 58382 111012 58442
rect 52196 58380 52202 58382
rect 111006 58380 111012 58382
rect 111076 58380 111082 58444
rect 217542 58380 217548 58444
rect 217612 58442 217618 58444
rect 257838 58442 257844 58444
rect 217612 58382 257844 58442
rect 217612 58380 217618 58382
rect 257838 58380 257844 58382
rect 257908 58380 257914 58444
rect 367686 58380 367692 58444
rect 367756 58442 367762 58444
rect 453430 58442 453436 58444
rect 367756 58382 453436 58442
rect 367756 58380 367762 58382
rect 453430 58380 453436 58382
rect 453500 58380 453506 58444
rect 85430 58108 85436 58172
rect 85500 58108 85506 58172
rect 92238 58108 92244 58172
rect 92308 58108 92314 58172
rect 153326 58108 153332 58172
rect 153396 58108 153402 58172
rect 235942 58108 235948 58172
rect 236012 58108 236018 58172
rect 265198 58108 265204 58172
rect 265268 58108 265274 58172
rect 272190 58108 272196 58172
rect 272260 58108 272266 58172
rect 275686 58108 275692 58172
rect 275756 58108 275762 58172
rect 300894 58108 300900 58172
rect 300964 58108 300970 58172
rect 315798 58108 315804 58172
rect 315868 58108 315874 58172
rect 398230 58108 398236 58172
rect 398300 58108 398306 58172
rect 401726 58108 401732 58172
rect 401796 58108 401802 58172
rect 405406 58108 405412 58172
rect 405476 58108 405482 58172
rect 416078 58108 416084 58172
rect 416148 58108 416154 58172
rect 83958 57972 83964 58036
rect 84028 58034 84034 58036
rect 84193 58034 84259 58037
rect 84028 58032 84259 58034
rect 84028 57976 84198 58032
rect 84254 57976 84259 58032
rect 84028 57974 84259 57976
rect 84028 57972 84034 57974
rect 84193 57971 84259 57974
rect 85438 57901 85498 58108
rect 76005 57900 76071 57901
rect 78213 57900 78279 57901
rect 79501 57900 79567 57901
rect 76005 57896 76052 57900
rect 76116 57898 76122 57900
rect 76005 57840 76010 57896
rect 76005 57836 76052 57840
rect 76116 57838 76162 57898
rect 78213 57896 78260 57900
rect 78324 57898 78330 57900
rect 78213 57840 78218 57896
rect 76116 57836 76122 57838
rect 78213 57836 78260 57840
rect 78324 57838 78370 57898
rect 79501 57896 79548 57900
rect 79612 57898 79618 57900
rect 80053 57898 80119 57901
rect 80462 57898 80468 57900
rect 79501 57840 79506 57896
rect 78324 57836 78330 57838
rect 79501 57836 79548 57840
rect 79612 57838 79658 57898
rect 80053 57896 80468 57898
rect 80053 57840 80058 57896
rect 80114 57840 80468 57896
rect 80053 57838 80468 57840
rect 79612 57836 79618 57838
rect 76005 57835 76071 57836
rect 78213 57835 78279 57836
rect 79501 57835 79567 57836
rect 80053 57835 80119 57838
rect 80462 57836 80468 57838
rect 80532 57836 80538 57900
rect 81801 57898 81867 57901
rect 81934 57898 81940 57900
rect 81801 57896 81940 57898
rect 81801 57840 81806 57896
rect 81862 57840 81940 57896
rect 81801 57838 81940 57840
rect 81801 57835 81867 57838
rect 81934 57836 81940 57838
rect 82004 57836 82010 57900
rect 85389 57896 85498 57901
rect 85389 57840 85394 57896
rect 85450 57840 85498 57896
rect 85389 57838 85498 57840
rect 86493 57900 86559 57901
rect 86493 57896 86540 57900
rect 86604 57898 86610 57900
rect 86953 57898 87019 57901
rect 88333 57900 88399 57901
rect 88701 57900 88767 57901
rect 87638 57898 87644 57900
rect 86493 57840 86498 57896
rect 85389 57835 85455 57838
rect 86493 57836 86540 57840
rect 86604 57838 86650 57898
rect 86953 57896 87644 57898
rect 86953 57840 86958 57896
rect 87014 57840 87644 57896
rect 86953 57838 87644 57840
rect 86604 57836 86610 57838
rect 86493 57835 86559 57836
rect 86953 57835 87019 57838
rect 87638 57836 87644 57838
rect 87708 57836 87714 57900
rect 88333 57896 88380 57900
rect 88444 57898 88450 57900
rect 88333 57840 88338 57896
rect 88333 57836 88380 57840
rect 88444 57838 88490 57898
rect 88701 57896 88748 57900
rect 88812 57898 88818 57900
rect 89713 57898 89779 57901
rect 90725 57900 90791 57901
rect 90030 57898 90036 57900
rect 88701 57840 88706 57896
rect 88444 57836 88450 57838
rect 88701 57836 88748 57840
rect 88812 57838 88858 57898
rect 89713 57896 90036 57898
rect 89713 57840 89718 57896
rect 89774 57840 90036 57896
rect 89713 57838 90036 57840
rect 88812 57836 88818 57838
rect 88333 57835 88399 57836
rect 88701 57835 88767 57836
rect 89713 57835 89779 57838
rect 90030 57836 90036 57838
rect 90100 57836 90106 57900
rect 90725 57896 90772 57900
rect 90836 57898 90842 57900
rect 91185 57898 91251 57901
rect 91318 57898 91324 57900
rect 90725 57840 90730 57896
rect 90725 57836 90772 57840
rect 90836 57838 90882 57898
rect 91185 57896 91324 57898
rect 91185 57840 91190 57896
rect 91246 57840 91324 57896
rect 91185 57838 91324 57840
rect 90836 57836 90842 57838
rect 90725 57835 90791 57836
rect 91185 57835 91251 57838
rect 91318 57836 91324 57838
rect 91388 57836 91394 57900
rect 92105 57898 92171 57901
rect 92246 57898 92306 58108
rect 153334 57901 153394 58108
rect 235950 57901 236010 58108
rect 92105 57896 92306 57898
rect 92105 57840 92110 57896
rect 92166 57840 92306 57896
rect 92105 57838 92306 57840
rect 92473 57898 92539 57901
rect 93669 57900 93735 57901
rect 98085 57900 98151 57901
rect 106365 57900 106431 57901
rect 93342 57898 93348 57900
rect 92473 57896 93348 57898
rect 92473 57840 92478 57896
rect 92534 57840 93348 57896
rect 92473 57838 93348 57840
rect 92105 57835 92171 57838
rect 92473 57835 92539 57838
rect 93342 57836 93348 57838
rect 93412 57836 93418 57900
rect 93669 57896 93716 57900
rect 93780 57898 93786 57900
rect 93669 57840 93674 57896
rect 93669 57836 93716 57840
rect 93780 57838 93826 57898
rect 98085 57896 98132 57900
rect 98196 57898 98202 57900
rect 98085 57840 98090 57896
rect 93780 57836 93786 57838
rect 98085 57836 98132 57840
rect 98196 57838 98242 57898
rect 106365 57896 106412 57900
rect 106476 57898 106482 57900
rect 107377 57898 107443 57901
rect 107510 57898 107516 57900
rect 106365 57840 106370 57896
rect 98196 57836 98202 57838
rect 106365 57836 106412 57840
rect 106476 57838 106522 57898
rect 107377 57896 107516 57898
rect 107377 57840 107382 57896
rect 107438 57840 107516 57896
rect 107377 57838 107516 57840
rect 106476 57836 106482 57838
rect 93669 57835 93735 57836
rect 98085 57835 98151 57836
rect 106365 57835 106431 57836
rect 107377 57835 107443 57838
rect 107510 57836 107516 57838
rect 107580 57836 107586 57900
rect 108021 57898 108087 57901
rect 112069 57900 112135 57901
rect 113173 57900 113239 57901
rect 123477 57900 123543 57901
rect 130837 57900 130903 57901
rect 108614 57898 108620 57900
rect 108021 57896 108620 57898
rect 108021 57840 108026 57896
rect 108082 57840 108620 57896
rect 108021 57838 108620 57840
rect 108021 57835 108087 57838
rect 108614 57836 108620 57838
rect 108684 57836 108690 57900
rect 112069 57896 112116 57900
rect 112180 57898 112186 57900
rect 112069 57840 112074 57896
rect 112069 57836 112116 57840
rect 112180 57838 112226 57898
rect 113173 57896 113220 57900
rect 113284 57898 113290 57900
rect 113173 57840 113178 57896
rect 112180 57836 112186 57838
rect 113173 57836 113220 57840
rect 113284 57838 113330 57898
rect 123477 57896 123524 57900
rect 123588 57898 123594 57900
rect 123477 57840 123482 57896
rect 113284 57836 113290 57838
rect 123477 57836 123524 57840
rect 123588 57838 123634 57898
rect 130837 57896 130884 57900
rect 130948 57898 130954 57900
rect 133229 57898 133295 57901
rect 145557 57900 145623 57901
rect 133454 57898 133460 57900
rect 130837 57840 130842 57896
rect 123588 57836 123594 57838
rect 130837 57836 130884 57840
rect 130948 57838 130994 57898
rect 133229 57896 133460 57898
rect 133229 57840 133234 57896
rect 133290 57840 133460 57896
rect 133229 57838 133460 57840
rect 130948 57836 130954 57838
rect 112069 57835 112135 57836
rect 113173 57835 113239 57836
rect 123477 57835 123543 57836
rect 130837 57835 130903 57836
rect 133229 57835 133295 57838
rect 133454 57836 133460 57838
rect 133524 57836 133530 57900
rect 145557 57896 145604 57900
rect 145668 57898 145674 57900
rect 145557 57840 145562 57896
rect 145557 57836 145604 57840
rect 145668 57838 145714 57898
rect 153285 57896 153394 57901
rect 153285 57840 153290 57896
rect 153346 57840 153394 57896
rect 153285 57838 153394 57840
rect 157425 57898 157491 57901
rect 158478 57898 158484 57900
rect 157425 57896 158484 57898
rect 157425 57840 157430 57896
rect 157486 57840 158484 57896
rect 157425 57838 158484 57840
rect 145668 57836 145674 57838
rect 145557 57835 145623 57836
rect 153285 57835 153351 57838
rect 157425 57835 157491 57838
rect 158478 57836 158484 57838
rect 158548 57836 158554 57900
rect 183134 57836 183140 57900
rect 183204 57898 183210 57900
rect 183277 57898 183343 57901
rect 183204 57896 183343 57898
rect 183204 57840 183282 57896
rect 183338 57840 183343 57896
rect 183204 57838 183343 57840
rect 235950 57896 236059 57901
rect 235950 57840 235998 57896
rect 236054 57840 236059 57896
rect 235950 57838 236059 57840
rect 183204 57836 183210 57838
rect 183277 57835 183343 57838
rect 235993 57835 236059 57838
rect 237373 57898 237439 57901
rect 239213 57900 239279 57901
rect 238150 57898 238156 57900
rect 237373 57896 238156 57898
rect 237373 57840 237378 57896
rect 237434 57840 238156 57896
rect 237373 57838 238156 57840
rect 237373 57835 237439 57838
rect 238150 57836 238156 57838
rect 238220 57836 238226 57900
rect 239213 57896 239260 57900
rect 239324 57898 239330 57900
rect 240133 57898 240199 57901
rect 241605 57900 241671 57901
rect 242893 57900 242959 57901
rect 240542 57898 240548 57900
rect 239213 57840 239218 57896
rect 239213 57836 239260 57840
rect 239324 57838 239370 57898
rect 240133 57896 240548 57898
rect 240133 57840 240138 57896
rect 240194 57840 240548 57896
rect 240133 57838 240548 57840
rect 239324 57836 239330 57838
rect 239213 57835 239279 57836
rect 240133 57835 240199 57838
rect 240542 57836 240548 57838
rect 240612 57836 240618 57900
rect 241605 57896 241652 57900
rect 241716 57898 241722 57900
rect 241605 57840 241610 57896
rect 241605 57836 241652 57840
rect 241716 57838 241762 57898
rect 242893 57896 242940 57900
rect 243004 57898 243010 57900
rect 242893 57840 242898 57896
rect 241716 57836 241722 57838
rect 242893 57836 242940 57840
rect 243004 57838 243050 57898
rect 243004 57836 243010 57838
rect 244222 57836 244228 57900
rect 244292 57898 244298 57900
rect 244365 57898 244431 57901
rect 244292 57896 244431 57898
rect 244292 57840 244370 57896
rect 244426 57840 244431 57896
rect 244292 57838 244431 57840
rect 244292 57836 244298 57838
rect 241605 57835 241671 57836
rect 242893 57835 242959 57836
rect 244365 57835 244431 57838
rect 245285 57900 245351 57901
rect 245285 57896 245332 57900
rect 245396 57898 245402 57900
rect 245653 57898 245719 57901
rect 246430 57898 246436 57900
rect 245285 57840 245290 57896
rect 245285 57836 245332 57840
rect 245396 57838 245442 57898
rect 245653 57896 246436 57898
rect 245653 57840 245658 57896
rect 245714 57840 246436 57896
rect 245653 57838 246436 57840
rect 245396 57836 245402 57838
rect 245285 57835 245351 57836
rect 245653 57835 245719 57838
rect 246430 57836 246436 57838
rect 246500 57836 246506 57900
rect 247033 57898 247099 57901
rect 248597 57900 248663 57901
rect 247718 57898 247724 57900
rect 247033 57896 247724 57898
rect 247033 57840 247038 57896
rect 247094 57840 247724 57896
rect 247033 57838 247724 57840
rect 247033 57835 247099 57838
rect 247718 57836 247724 57838
rect 247788 57836 247794 57900
rect 248597 57896 248644 57900
rect 248708 57898 248714 57900
rect 249793 57898 249859 57901
rect 251173 57900 251239 57901
rect 250110 57898 250116 57900
rect 248597 57840 248602 57896
rect 248597 57836 248644 57840
rect 248708 57838 248754 57898
rect 249793 57896 250116 57898
rect 249793 57840 249798 57896
rect 249854 57840 250116 57896
rect 249793 57838 250116 57840
rect 248708 57836 248714 57838
rect 248597 57835 248663 57836
rect 249793 57835 249859 57838
rect 250110 57836 250116 57838
rect 250180 57836 250186 57900
rect 251173 57898 251220 57900
rect 251128 57896 251220 57898
rect 251128 57840 251178 57896
rect 251128 57838 251220 57840
rect 251173 57836 251220 57838
rect 251284 57836 251290 57900
rect 251357 57898 251423 57901
rect 253381 57900 253447 57901
rect 252318 57898 252324 57900
rect 251357 57896 252324 57898
rect 251357 57840 251362 57896
rect 251418 57840 252324 57896
rect 251357 57838 252324 57840
rect 251173 57835 251239 57836
rect 251357 57835 251423 57838
rect 252318 57836 252324 57838
rect 252388 57836 252394 57900
rect 253381 57896 253428 57900
rect 253492 57898 253498 57900
rect 253933 57898 253999 57901
rect 254526 57898 254532 57900
rect 253381 57840 253386 57896
rect 253381 57836 253428 57840
rect 253492 57838 253538 57898
rect 253933 57896 254532 57898
rect 253933 57840 253938 57896
rect 253994 57840 254532 57896
rect 253933 57838 254532 57840
rect 253492 57836 253498 57838
rect 253381 57835 253447 57836
rect 253933 57835 253999 57838
rect 254526 57836 254532 57838
rect 254596 57836 254602 57900
rect 264973 57898 265039 57901
rect 265206 57898 265266 58108
rect 264973 57896 265266 57898
rect 264973 57840 264978 57896
rect 265034 57840 265266 57896
rect 264973 57838 265266 57840
rect 265893 57900 265959 57901
rect 266353 57900 266419 57901
rect 265893 57896 265940 57900
rect 266004 57898 266010 57900
rect 266302 57898 266308 57900
rect 265893 57840 265898 57896
rect 264973 57835 265039 57838
rect 265893 57836 265940 57840
rect 266004 57838 266050 57898
rect 266262 57838 266308 57898
rect 266372 57896 266419 57900
rect 266414 57840 266419 57896
rect 266004 57836 266010 57838
rect 266302 57836 266308 57838
rect 266372 57836 266419 57840
rect 265893 57835 265959 57836
rect 266353 57835 266419 57836
rect 268469 57898 268535 57901
rect 271229 57900 271295 57901
rect 268694 57898 268700 57900
rect 268469 57896 268700 57898
rect 268469 57840 268474 57896
rect 268530 57840 268700 57896
rect 268469 57838 268700 57840
rect 268469 57835 268535 57838
rect 268694 57836 268700 57838
rect 268764 57836 268770 57900
rect 271229 57896 271276 57900
rect 271340 57898 271346 57900
rect 271873 57898 271939 57901
rect 272198 57898 272258 58108
rect 271229 57840 271234 57896
rect 271229 57836 271276 57840
rect 271340 57838 271386 57898
rect 271873 57896 272258 57898
rect 271873 57840 271878 57896
rect 271934 57840 272258 57896
rect 271873 57838 272258 57840
rect 273253 57900 273319 57901
rect 273253 57896 273300 57900
rect 273364 57898 273370 57900
rect 275461 57898 275527 57901
rect 275694 57898 275754 58108
rect 300902 57901 300962 58108
rect 315806 57901 315866 58108
rect 273253 57840 273258 57896
rect 271340 57836 271346 57838
rect 271229 57835 271295 57836
rect 271873 57835 271939 57838
rect 273253 57836 273300 57840
rect 273364 57838 273410 57898
rect 275461 57896 275754 57898
rect 275461 57840 275466 57896
rect 275522 57840 275754 57896
rect 275461 57838 275754 57840
rect 287605 57898 287671 57901
rect 293309 57900 293375 57901
rect 295885 57900 295951 57901
rect 288198 57898 288204 57900
rect 287605 57896 288204 57898
rect 287605 57840 287610 57896
rect 287666 57840 288204 57896
rect 287605 57838 288204 57840
rect 273364 57836 273370 57838
rect 273253 57835 273319 57836
rect 275461 57835 275527 57838
rect 287605 57835 287671 57838
rect 288198 57836 288204 57838
rect 288268 57836 288274 57900
rect 293309 57896 293356 57900
rect 293420 57898 293426 57900
rect 293309 57840 293314 57896
rect 293309 57836 293356 57840
rect 293420 57838 293466 57898
rect 295885 57896 295932 57900
rect 295996 57898 296002 57900
rect 295885 57840 295890 57896
rect 293420 57836 293426 57838
rect 295885 57836 295932 57840
rect 295996 57838 296042 57898
rect 300853 57896 300962 57901
rect 300853 57840 300858 57896
rect 300914 57840 300962 57896
rect 300853 57838 300962 57840
rect 303429 57900 303495 57901
rect 303429 57896 303476 57900
rect 303540 57898 303546 57900
rect 308489 57898 308555 57901
rect 310973 57900 311039 57901
rect 308622 57898 308628 57900
rect 303429 57840 303434 57896
rect 295996 57836 296002 57838
rect 293309 57835 293375 57836
rect 295885 57835 295951 57836
rect 300853 57835 300919 57838
rect 303429 57836 303476 57840
rect 303540 57838 303586 57898
rect 308489 57896 308628 57898
rect 308489 57840 308494 57896
rect 308550 57840 308628 57896
rect 308489 57838 308628 57840
rect 303540 57836 303546 57838
rect 303429 57835 303495 57836
rect 308489 57835 308555 57838
rect 308622 57836 308628 57838
rect 308692 57836 308698 57900
rect 310973 57896 311020 57900
rect 311084 57898 311090 57900
rect 310973 57840 310978 57896
rect 310973 57836 311020 57840
rect 311084 57838 311130 57898
rect 315757 57896 315866 57901
rect 315757 57840 315762 57896
rect 315818 57840 315866 57896
rect 315757 57838 315866 57840
rect 320909 57900 320975 57901
rect 323301 57900 323367 57901
rect 343173 57900 343239 57901
rect 343449 57900 343515 57901
rect 320909 57896 320956 57900
rect 321020 57898 321026 57900
rect 320909 57840 320914 57896
rect 311084 57836 311090 57838
rect 310973 57835 311039 57836
rect 315757 57835 315823 57838
rect 320909 57836 320956 57840
rect 321020 57838 321066 57898
rect 323301 57896 323348 57900
rect 323412 57898 323418 57900
rect 343173 57898 343220 57900
rect 323301 57840 323306 57896
rect 321020 57836 321026 57838
rect 323301 57836 323348 57840
rect 323412 57838 323458 57898
rect 343128 57896 343220 57898
rect 343128 57840 343178 57896
rect 343128 57838 343220 57840
rect 323412 57836 323418 57838
rect 343173 57836 343220 57838
rect 343284 57836 343290 57900
rect 343398 57898 343404 57900
rect 343358 57838 343404 57898
rect 343468 57896 343515 57900
rect 343510 57840 343515 57896
rect 343398 57836 343404 57838
rect 343468 57836 343515 57840
rect 320909 57835 320975 57836
rect 323301 57835 323367 57836
rect 343173 57835 343239 57836
rect 343449 57835 343515 57836
rect 397453 57898 397519 57901
rect 398238 57898 398298 58108
rect 401734 57901 401794 58108
rect 397453 57896 398298 57898
rect 397453 57840 397458 57896
rect 397514 57840 398298 57896
rect 397453 57838 398298 57840
rect 399477 57900 399543 57901
rect 399477 57896 399524 57900
rect 399588 57898 399594 57900
rect 400213 57898 400279 57901
rect 400438 57898 400444 57900
rect 399477 57840 399482 57896
rect 397453 57835 397519 57838
rect 399477 57836 399524 57840
rect 399588 57838 399634 57898
rect 400213 57896 400444 57898
rect 400213 57840 400218 57896
rect 400274 57840 400444 57896
rect 400213 57838 400444 57840
rect 399588 57836 399594 57838
rect 399477 57835 399543 57836
rect 400213 57835 400279 57838
rect 400438 57836 400444 57838
rect 400508 57836 400514 57900
rect 401685 57896 401794 57901
rect 401685 57840 401690 57896
rect 401746 57840 401794 57896
rect 401685 57838 401794 57840
rect 404353 57898 404419 57901
rect 405414 57898 405474 58108
rect 416086 57901 416146 58108
rect 404353 57896 405474 57898
rect 404353 57840 404358 57896
rect 404414 57840 405474 57896
rect 404353 57838 405474 57840
rect 405825 57898 405891 57901
rect 406510 57898 406516 57900
rect 405825 57896 406516 57898
rect 405825 57840 405830 57896
rect 405886 57840 406516 57896
rect 405825 57838 406516 57840
rect 401685 57835 401751 57838
rect 404353 57835 404419 57838
rect 405825 57835 405891 57838
rect 406510 57836 406516 57838
rect 406580 57836 406586 57900
rect 407205 57898 407271 57901
rect 408309 57900 408375 57901
rect 408677 57900 408743 57901
rect 407614 57898 407620 57900
rect 407205 57896 407620 57898
rect 407205 57840 407210 57896
rect 407266 57840 407620 57896
rect 407205 57838 407620 57840
rect 407205 57835 407271 57838
rect 407614 57836 407620 57838
rect 407684 57836 407690 57900
rect 408309 57896 408356 57900
rect 408420 57898 408426 57900
rect 408309 57840 408314 57896
rect 408309 57836 408356 57840
rect 408420 57838 408466 57898
rect 408677 57896 408724 57900
rect 408788 57898 408794 57900
rect 409873 57898 409939 57901
rect 410006 57898 410012 57900
rect 408677 57840 408682 57896
rect 408420 57836 408426 57838
rect 408677 57836 408724 57840
rect 408788 57838 408834 57898
rect 409873 57896 410012 57898
rect 409873 57840 409878 57896
rect 409934 57840 410012 57896
rect 409873 57838 410012 57840
rect 408788 57836 408794 57838
rect 408309 57835 408375 57836
rect 408677 57835 408743 57836
rect 409873 57835 409939 57838
rect 410006 57836 410012 57838
rect 410076 57836 410082 57900
rect 411345 57898 411411 57901
rect 414565 57900 414631 57901
rect 415485 57900 415551 57901
rect 412398 57898 412404 57900
rect 411345 57896 412404 57898
rect 411345 57840 411350 57896
rect 411406 57840 412404 57896
rect 411345 57838 412404 57840
rect 411345 57835 411411 57838
rect 412398 57836 412404 57838
rect 412468 57836 412474 57900
rect 414565 57896 414612 57900
rect 414676 57898 414682 57900
rect 414565 57840 414570 57896
rect 414565 57836 414612 57840
rect 414676 57838 414722 57898
rect 415485 57896 415532 57900
rect 415596 57898 415602 57900
rect 415485 57840 415490 57896
rect 414676 57836 414682 57838
rect 415485 57836 415532 57840
rect 415596 57838 415642 57898
rect 416037 57896 416146 57901
rect 426433 57900 426499 57901
rect 426382 57898 426388 57900
rect 416037 57840 416042 57896
rect 416098 57840 416146 57896
rect 416037 57838 416146 57840
rect 426342 57838 426388 57898
rect 426452 57896 426499 57900
rect 427629 57900 427695 57901
rect 427629 57898 427676 57900
rect 426494 57840 426499 57896
rect 415596 57836 415602 57838
rect 414565 57835 414631 57836
rect 415485 57835 415551 57836
rect 416037 57835 416103 57838
rect 426382 57836 426388 57838
rect 426452 57836 426499 57840
rect 427584 57896 427676 57898
rect 427584 57840 427634 57896
rect 427584 57838 427676 57840
rect 426433 57835 426499 57836
rect 427629 57836 427676 57838
rect 427740 57836 427746 57900
rect 427813 57898 427879 57901
rect 428590 57898 428596 57900
rect 427813 57896 428596 57898
rect 427813 57840 427818 57896
rect 427874 57840 428596 57896
rect 427813 57838 428596 57840
rect 427629 57835 427695 57836
rect 427813 57835 427879 57838
rect 428590 57836 428596 57838
rect 428660 57836 428666 57900
rect 429193 57898 429259 57901
rect 429694 57898 429700 57900
rect 429193 57896 429700 57898
rect 429193 57840 429198 57896
rect 429254 57840 429700 57896
rect 429193 57838 429700 57840
rect 429193 57835 429259 57838
rect 429694 57836 429700 57838
rect 429764 57836 429770 57900
rect 430573 57898 430639 57901
rect 431166 57898 431172 57900
rect 430573 57896 431172 57898
rect 430573 57840 430578 57896
rect 430634 57840 431172 57896
rect 430573 57838 431172 57840
rect 430573 57835 430639 57838
rect 431166 57836 431172 57838
rect 431236 57836 431242 57900
rect 431953 57898 432019 57901
rect 432270 57898 432276 57900
rect 431953 57896 432276 57898
rect 431953 57840 431958 57896
rect 432014 57840 432276 57896
rect 431953 57838 432276 57840
rect 431953 57835 432019 57838
rect 432270 57836 432276 57838
rect 432340 57836 432346 57900
rect 433425 57898 433491 57901
rect 435909 57900 435975 57901
rect 434662 57898 434668 57900
rect 433425 57896 434668 57898
rect 433425 57840 433430 57896
rect 433486 57840 434668 57896
rect 433425 57838 434668 57840
rect 433425 57835 433491 57838
rect 434662 57836 434668 57838
rect 434732 57836 434738 57900
rect 435909 57898 435956 57900
rect 435864 57896 435956 57898
rect 435864 57840 435914 57896
rect 435864 57838 435956 57840
rect 435909 57836 435956 57838
rect 436020 57836 436026 57900
rect 436093 57898 436159 57901
rect 438301 57900 438367 57901
rect 438485 57900 438551 57901
rect 436870 57898 436876 57900
rect 436093 57896 436876 57898
rect 436093 57840 436098 57896
rect 436154 57840 436876 57896
rect 436093 57838 436876 57840
rect 435909 57835 435975 57836
rect 436093 57835 436159 57838
rect 436870 57836 436876 57838
rect 436940 57836 436946 57900
rect 438301 57898 438348 57900
rect 438256 57896 438348 57898
rect 438256 57840 438306 57896
rect 438256 57838 438348 57840
rect 438301 57836 438348 57838
rect 438412 57836 438418 57900
rect 438485 57896 438532 57900
rect 438596 57898 438602 57900
rect 438853 57898 438919 57901
rect 440877 57900 440943 57901
rect 443453 57900 443519 57901
rect 445845 57900 445911 57901
rect 450997 57900 451063 57901
rect 478413 57900 478479 57901
rect 503345 57900 503411 57901
rect 439078 57898 439084 57900
rect 438485 57840 438490 57896
rect 438485 57836 438532 57840
rect 438596 57838 438642 57898
rect 438853 57896 439084 57898
rect 438853 57840 438858 57896
rect 438914 57840 439084 57896
rect 438853 57838 439084 57840
rect 438596 57836 438602 57838
rect 438301 57835 438367 57836
rect 438485 57835 438551 57836
rect 438853 57835 438919 57838
rect 439078 57836 439084 57838
rect 439148 57836 439154 57900
rect 440877 57896 440924 57900
rect 440988 57898 440994 57900
rect 440877 57840 440882 57896
rect 440877 57836 440924 57840
rect 440988 57838 441034 57898
rect 443453 57896 443500 57900
rect 443564 57898 443570 57900
rect 443453 57840 443458 57896
rect 440988 57836 440994 57838
rect 443453 57836 443500 57840
rect 443564 57838 443610 57898
rect 445845 57896 445892 57900
rect 445956 57898 445962 57900
rect 445845 57840 445850 57896
rect 443564 57836 443570 57838
rect 445845 57836 445892 57840
rect 445956 57838 446002 57898
rect 450997 57896 451044 57900
rect 451108 57898 451114 57900
rect 450997 57840 451002 57896
rect 445956 57836 445962 57838
rect 450997 57836 451044 57840
rect 451108 57838 451154 57898
rect 478413 57896 478460 57900
rect 478524 57898 478530 57900
rect 503294 57898 503300 57900
rect 478413 57840 478418 57896
rect 451108 57836 451114 57838
rect 478413 57836 478460 57840
rect 478524 57838 478570 57898
rect 503254 57838 503300 57898
rect 503364 57896 503411 57900
rect 503406 57840 503411 57896
rect 478524 57836 478530 57838
rect 503294 57836 503300 57838
rect 503364 57836 503411 57840
rect 440877 57835 440943 57836
rect 443453 57835 443519 57836
rect 445845 57835 445911 57836
rect 450997 57835 451063 57836
rect 478413 57835 478479 57836
rect 503345 57835 503411 57836
rect 183461 57764 183527 57765
rect 60222 57700 60228 57764
rect 60292 57762 60298 57764
rect 125910 57762 125916 57764
rect 60292 57702 125916 57762
rect 60292 57700 60298 57702
rect 125910 57700 125916 57702
rect 125980 57700 125986 57764
rect 183461 57760 183508 57764
rect 183572 57762 183578 57764
rect 183461 57704 183466 57760
rect 183461 57700 183508 57704
rect 183572 57702 183618 57762
rect 183572 57700 183578 57702
rect 214414 57700 214420 57764
rect 214484 57762 214490 57764
rect 280838 57762 280844 57764
rect 214484 57702 280844 57762
rect 214484 57700 214490 57702
rect 280838 57700 280844 57702
rect 280908 57700 280914 57764
rect 378726 57700 378732 57764
rect 378796 57762 378802 57764
rect 473302 57762 473308 57764
rect 378796 57702 473308 57762
rect 378796 57700 378802 57702
rect 473302 57700 473308 57702
rect 473372 57700 473378 57764
rect 183461 57699 183527 57700
rect 55070 57564 55076 57628
rect 55140 57626 55146 57628
rect 109033 57626 109099 57629
rect 109534 57626 109540 57628
rect 55140 57566 103530 57626
rect 55140 57564 55146 57566
rect 58934 57428 58940 57492
rect 59004 57490 59010 57492
rect 98637 57490 98703 57493
rect 59004 57488 98703 57490
rect 59004 57432 98642 57488
rect 98698 57432 98703 57488
rect 59004 57430 98703 57432
rect 103470 57490 103530 57566
rect 109033 57624 109540 57626
rect 109033 57568 109038 57624
rect 109094 57568 109540 57624
rect 109033 57566 109540 57568
rect 109033 57563 109099 57566
rect 109534 57564 109540 57566
rect 109604 57564 109610 57628
rect 113265 57626 113331 57629
rect 114318 57626 114324 57628
rect 113265 57624 114324 57626
rect 113265 57568 113270 57624
rect 113326 57568 114324 57624
rect 113265 57566 114324 57568
rect 113265 57563 113331 57566
rect 114318 57564 114324 57566
rect 114388 57564 114394 57628
rect 114553 57626 114619 57629
rect 115790 57626 115796 57628
rect 114553 57624 115796 57626
rect 114553 57568 114558 57624
rect 114614 57568 115796 57624
rect 114553 57566 115796 57568
rect 114553 57563 114619 57566
rect 115790 57564 115796 57566
rect 115860 57564 115866 57628
rect 116117 57626 116183 57629
rect 116894 57626 116900 57628
rect 116117 57624 116900 57626
rect 116117 57568 116122 57624
rect 116178 57568 116900 57624
rect 116117 57566 116900 57568
rect 116117 57563 116183 57566
rect 116894 57564 116900 57566
rect 116964 57564 116970 57628
rect 117313 57626 117379 57629
rect 117998 57626 118004 57628
rect 117313 57624 118004 57626
rect 117313 57568 117318 57624
rect 117374 57568 118004 57624
rect 117313 57566 118004 57568
rect 117313 57563 117379 57566
rect 117998 57564 118004 57566
rect 118068 57564 118074 57628
rect 118693 57626 118759 57629
rect 155953 57628 156019 57629
rect 119102 57626 119108 57628
rect 118693 57624 119108 57626
rect 118693 57568 118698 57624
rect 118754 57568 119108 57624
rect 118693 57566 119108 57568
rect 118693 57563 118759 57566
rect 119102 57564 119108 57566
rect 119172 57564 119178 57628
rect 155902 57626 155908 57628
rect 155862 57566 155908 57626
rect 155972 57624 156019 57628
rect 156014 57568 156019 57624
rect 155902 57564 155908 57566
rect 155972 57564 156019 57568
rect 155953 57563 156019 57564
rect 160093 57626 160159 57629
rect 160870 57626 160876 57628
rect 160093 57624 160876 57626
rect 160093 57568 160098 57624
rect 160154 57568 160876 57624
rect 160093 57566 160876 57568
rect 160093 57563 160159 57566
rect 160870 57564 160876 57566
rect 160940 57564 160946 57628
rect 165613 57626 165679 57629
rect 165838 57626 165844 57628
rect 165613 57624 165844 57626
rect 165613 57568 165618 57624
rect 165674 57568 165844 57624
rect 165613 57566 165844 57568
rect 165613 57563 165679 57566
rect 165838 57564 165844 57566
rect 165908 57564 165914 57628
rect 209078 57564 209084 57628
rect 209148 57626 209154 57628
rect 266445 57626 266511 57629
rect 267590 57626 267596 57628
rect 209148 57566 262908 57626
rect 209148 57564 209154 57566
rect 118366 57490 118372 57492
rect 103470 57430 118372 57490
rect 59004 57428 59010 57430
rect 98637 57427 98703 57430
rect 118366 57428 118372 57430
rect 118436 57428 118442 57492
rect 202270 57428 202276 57492
rect 202340 57490 202346 57492
rect 258390 57490 258396 57492
rect 202340 57430 258396 57490
rect 202340 57428 202346 57430
rect 258390 57428 258396 57430
rect 258460 57428 258466 57492
rect 262848 57490 262908 57566
rect 266445 57624 267596 57626
rect 266445 57568 266450 57624
rect 266506 57568 267596 57624
rect 266445 57566 267596 57568
rect 266445 57563 266511 57566
rect 267590 57564 267596 57566
rect 267660 57564 267666 57628
rect 269113 57626 269179 57629
rect 269798 57626 269804 57628
rect 269113 57624 269804 57626
rect 269113 57568 269118 57624
rect 269174 57568 269804 57624
rect 269113 57566 269804 57568
rect 269113 57563 269179 57566
rect 269798 57564 269804 57566
rect 269868 57564 269874 57628
rect 273345 57626 273411 57629
rect 274398 57626 274404 57628
rect 273345 57624 274404 57626
rect 273345 57568 273350 57624
rect 273406 57568 274404 57624
rect 273345 57566 274404 57568
rect 273345 57563 273411 57566
rect 274398 57564 274404 57566
rect 274468 57564 274474 57628
rect 276013 57626 276079 57629
rect 276974 57626 276980 57628
rect 276013 57624 276980 57626
rect 276013 57568 276018 57624
rect 276074 57568 276980 57624
rect 276013 57566 276980 57568
rect 276013 57563 276079 57566
rect 276974 57564 276980 57566
rect 277044 57564 277050 57628
rect 371918 57564 371924 57628
rect 371988 57626 371994 57628
rect 460974 57626 460980 57628
rect 371988 57566 460980 57626
rect 371988 57564 371994 57566
rect 460974 57564 460980 57566
rect 461044 57564 461050 57628
rect 270902 57490 270908 57492
rect 262848 57430 270908 57490
rect 270902 57428 270908 57430
rect 270972 57428 270978 57492
rect 378910 57428 378916 57492
rect 378980 57490 378986 57492
rect 456374 57490 456380 57492
rect 378980 57430 456380 57490
rect 378980 57428 378986 57430
rect 456374 57428 456380 57430
rect 456444 57428 456450 57492
rect 58750 57292 58756 57356
rect 58820 57354 58826 57356
rect 103830 57354 103836 57356
rect 58820 57294 103836 57354
rect 58820 57292 58826 57294
rect 103830 57292 103836 57294
rect 103900 57292 103906 57356
rect 204846 57292 204852 57356
rect 204916 57354 204922 57356
rect 255998 57354 256004 57356
rect 204916 57294 256004 57354
rect 204916 57292 204922 57294
rect 255998 57292 256004 57294
rect 256068 57292 256074 57356
rect 376150 57292 376156 57356
rect 376220 57354 376226 57356
rect 448278 57354 448284 57356
rect 376220 57294 448284 57354
rect 376220 57292 376226 57294
rect 448278 57292 448284 57294
rect 448348 57292 448354 57356
rect 430941 57220 431007 57221
rect 433333 57220 433399 57221
rect 433517 57220 433583 57221
rect 435725 57220 435791 57221
rect 59118 57156 59124 57220
rect 59188 57218 59194 57220
rect 98494 57218 98500 57220
rect 59188 57158 98500 57218
rect 59188 57156 59194 57158
rect 98494 57156 98500 57158
rect 98564 57156 98570 57220
rect 213126 57156 213132 57220
rect 213196 57218 213202 57220
rect 260966 57218 260972 57220
rect 213196 57158 260972 57218
rect 213196 57156 213202 57158
rect 260966 57156 260972 57158
rect 261036 57156 261042 57220
rect 379278 57156 379284 57220
rect 379348 57218 379354 57220
rect 421046 57218 421052 57220
rect 379348 57158 421052 57218
rect 379348 57156 379354 57158
rect 421046 57156 421052 57158
rect 421116 57156 421122 57220
rect 430941 57216 430988 57220
rect 431052 57218 431058 57220
rect 433333 57218 433380 57220
rect 430941 57160 430946 57216
rect 430941 57156 430988 57160
rect 431052 57158 431098 57218
rect 433288 57216 433380 57218
rect 433288 57160 433338 57216
rect 433288 57158 433380 57160
rect 431052 57156 431058 57158
rect 433333 57156 433380 57158
rect 433444 57156 433450 57220
rect 433517 57216 433564 57220
rect 433628 57218 433634 57220
rect 433517 57160 433522 57216
rect 433517 57156 433564 57160
rect 433628 57158 433674 57218
rect 435725 57216 435772 57220
rect 435836 57218 435842 57220
rect 435725 57160 435730 57216
rect 433628 57156 433634 57158
rect 435725 57156 435772 57160
rect 435836 57158 435882 57218
rect 435836 57156 435842 57158
rect 430941 57155 431007 57156
rect 433333 57155 433399 57156
rect 433517 57155 433583 57156
rect 435725 57155 435791 57156
rect 58566 57020 58572 57084
rect 58636 57082 58642 57084
rect 96286 57082 96292 57084
rect 58636 57022 96292 57082
rect 58636 57020 58642 57022
rect 96286 57020 96292 57022
rect 96356 57020 96362 57084
rect 98637 57082 98703 57085
rect 105854 57082 105860 57084
rect 98637 57080 105860 57082
rect 98637 57024 98642 57080
rect 98698 57024 105860 57080
rect 98637 57022 105860 57024
rect 98637 57019 98703 57022
rect 105854 57020 105860 57022
rect 105924 57020 105930 57084
rect 211654 57020 211660 57084
rect 211724 57082 211730 57084
rect 248270 57082 248276 57084
rect 211724 57022 248276 57082
rect 211724 57020 211730 57022
rect 248270 57020 248276 57022
rect 248340 57020 248346 57084
rect 379094 57020 379100 57084
rect 379164 57082 379170 57084
rect 413502 57082 413508 57084
rect 379164 57022 413508 57082
rect 379164 57020 379170 57022
rect 413502 57020 413508 57022
rect 413572 57020 413578 57084
rect 411253 56948 411319 56949
rect 411253 56944 411300 56948
rect 411364 56946 411370 56948
rect 412541 56946 412607 56949
rect 411253 56888 411258 56944
rect 411253 56884 411300 56888
rect 411364 56886 411410 56946
rect 412541 56944 412650 56946
rect 412541 56888 412546 56944
rect 412602 56888 412650 56944
rect 411364 56884 411370 56886
rect 411253 56883 411319 56884
rect 412541 56883 412650 56888
rect 412590 56813 412650 56883
rect 412590 56808 412699 56813
rect 412590 56752 412638 56808
rect 412694 56752 412699 56808
rect 412590 56750 412699 56752
rect 412633 56747 412699 56750
rect 54886 56612 54892 56676
rect 54956 56674 54962 56676
rect 128670 56674 128676 56676
rect 54956 56614 128676 56674
rect 54956 56612 54962 56614
rect 128670 56612 128676 56614
rect 128740 56612 128746 56676
rect 163262 56612 163268 56676
rect 163332 56612 163338 56676
rect 214598 56612 214604 56676
rect 214668 56674 214674 56676
rect 283782 56674 283788 56676
rect 214668 56614 283788 56674
rect 214668 56612 214674 56614
rect 283782 56612 283788 56614
rect 283852 56612 283858 56676
rect 363638 56612 363644 56676
rect 363708 56674 363714 56676
rect 468518 56674 468524 56676
rect 363708 56614 468524 56674
rect 363708 56612 363714 56614
rect 468518 56612 468524 56614
rect 468588 56612 468594 56676
rect 53598 56476 53604 56540
rect 53668 56538 53674 56540
rect 163270 56538 163330 56612
rect 53668 56478 163330 56538
rect 53668 56476 53674 56478
rect 219934 56476 219940 56540
rect 220004 56538 220010 56540
rect 410742 56538 410748 56540
rect 220004 56478 410748 56538
rect 220004 56476 220010 56478
rect 410742 56476 410748 56478
rect 410812 56476 410818 56540
rect 55622 56340 55628 56404
rect 55692 56402 55698 56404
rect 153285 56402 153351 56405
rect 55692 56400 153351 56402
rect 55692 56344 153290 56400
rect 153346 56344 153351 56400
rect 55692 56342 153351 56344
rect 55692 56340 55698 56342
rect 153285 56339 153351 56342
rect 200614 56340 200620 56404
rect 200684 56402 200690 56404
rect 268326 56402 268332 56404
rect 200684 56342 268332 56402
rect 200684 56340 200690 56342
rect 268326 56340 268332 56342
rect 268396 56340 268402 56404
rect 57646 56204 57652 56268
rect 57716 56266 57722 56268
rect 105302 56266 105308 56268
rect 57716 56206 105308 56266
rect 57716 56204 57722 56206
rect 105302 56204 105308 56206
rect 105372 56204 105378 56268
rect 217358 56204 217364 56268
rect 217428 56266 217434 56268
rect 277158 56266 277164 56268
rect 217428 56206 277164 56266
rect 217428 56204 217434 56206
rect 277158 56204 277164 56206
rect 277228 56204 277234 56268
rect 50470 55116 50476 55180
rect 50540 55178 50546 55180
rect 165613 55178 165679 55181
rect 50540 55176 165679 55178
rect 50540 55120 165618 55176
rect 165674 55120 165679 55176
rect 50540 55118 165679 55120
rect 50540 55116 50546 55118
rect 165613 55115 165679 55118
rect 217174 55116 217180 55180
rect 217244 55178 217250 55180
rect 276013 55178 276079 55181
rect 217244 55176 276079 55178
rect 217244 55120 276018 55176
rect 276074 55120 276079 55176
rect 217244 55118 276079 55120
rect 217244 55116 217250 55118
rect 276013 55115 276079 55118
rect 377622 55116 377628 55180
rect 377692 55178 377698 55180
rect 438853 55178 438919 55181
rect 377692 55176 438919 55178
rect 377692 55120 438858 55176
rect 438914 55120 438919 55176
rect 377692 55118 438919 55120
rect 377692 55116 377698 55118
rect 438853 55115 438919 55118
rect 50838 54980 50844 55044
rect 50908 55042 50914 55044
rect 160093 55042 160159 55045
rect 50908 55040 160159 55042
rect 50908 54984 160098 55040
rect 160154 54984 160159 55040
rect 50908 54982 160159 54984
rect 50908 54980 50914 54982
rect 160093 54979 160159 54982
rect 379462 54980 379468 55044
rect 379532 55042 379538 55044
rect 427813 55042 427879 55045
rect 379532 55040 427879 55042
rect 379532 54984 427818 55040
rect 427874 54984 427879 55040
rect 379532 54982 427879 54984
rect 379532 54980 379538 54982
rect 427813 54979 427879 54982
rect 50654 54844 50660 54908
rect 50724 54906 50730 54908
rect 155953 54906 156019 54909
rect 50724 54904 156019 54906
rect 50724 54848 155958 54904
rect 156014 54848 156019 54904
rect 50724 54846 156019 54848
rect 50724 54844 50730 54846
rect 155953 54843 156019 54846
rect 57462 54708 57468 54772
rect 57532 54770 57538 54772
rect 118693 54770 118759 54773
rect 57532 54768 118759 54770
rect 57532 54712 118698 54768
rect 118754 54712 118759 54768
rect 57532 54710 118759 54712
rect 57532 54708 57538 54710
rect 118693 54707 118759 54710
rect 57830 54572 57836 54636
rect 57900 54634 57906 54636
rect 116117 54634 116183 54637
rect 57900 54632 116183 54634
rect 57900 54576 116122 54632
rect 116178 54576 116183 54632
rect 57900 54574 116183 54576
rect 57900 54572 57906 54574
rect 116117 54571 116183 54574
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 580257 33146 580323 33149
rect 583520 33146 584960 33236
rect 580257 33144 584960 33146
rect 580257 33088 580262 33144
rect 580318 33088 584960 33144
rect 580257 33086 584960 33088
rect 580257 33083 580323 33086
rect 583520 32996 584960 33086
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19410 480 19500
rect 2773 19410 2839 19413
rect -960 19408 2839 19410
rect -960 19352 2778 19408
rect 2834 19352 2839 19408
rect -960 19350 2839 19352
rect -960 19260 480 19350
rect 2773 19347 2839 19350
rect -960 6340 480 6580
rect 583520 6476 584960 6716
rect 136449 4042 136515 4045
rect 208894 4042 208900 4044
rect 136449 4040 208900 4042
rect 136449 3984 136454 4040
rect 136510 3984 208900 4040
rect 136449 3982 208900 3984
rect 136449 3979 136515 3982
rect 208894 3980 208900 3982
rect 208964 3980 208970 4044
rect 132953 3906 133019 3909
rect 206134 3906 206140 3908
rect 132953 3904 206140 3906
rect 132953 3848 132958 3904
rect 133014 3848 206140 3904
rect 132953 3846 206140 3848
rect 132953 3843 133019 3846
rect 206134 3844 206140 3846
rect 206204 3844 206210 3908
rect 147121 3770 147187 3773
rect 365110 3770 365116 3772
rect 147121 3768 365116 3770
rect 147121 3712 147126 3768
rect 147182 3712 365116 3768
rect 147121 3710 365116 3712
rect 147121 3707 147187 3710
rect 365110 3708 365116 3710
rect 365180 3708 365186 3772
rect 143533 3634 143599 3637
rect 363454 3634 363460 3636
rect 143533 3632 363460 3634
rect 143533 3576 143538 3632
rect 143594 3576 363460 3632
rect 143533 3574 363460 3576
rect 143533 3571 143599 3574
rect 363454 3572 363460 3574
rect 363524 3572 363530 3636
rect 150617 3498 150683 3501
rect 374494 3498 374500 3500
rect 150617 3496 374500 3498
rect 150617 3440 150622 3496
rect 150678 3440 374500 3496
rect 150617 3438 374500 3440
rect 150617 3435 150683 3438
rect 374494 3436 374500 3438
rect 374564 3436 374570 3500
rect 129365 3362 129431 3365
rect 364926 3362 364932 3364
rect 129365 3360 364932 3362
rect 129365 3304 129370 3360
rect 129426 3304 364932 3360
rect 129365 3302 364932 3304
rect 129365 3299 129431 3302
rect 364926 3300 364932 3302
rect 364996 3300 365002 3364
rect 140037 3226 140103 3229
rect 210366 3226 210372 3228
rect 140037 3224 210372 3226
rect 140037 3168 140042 3224
rect 140098 3168 210372 3224
rect 140037 3166 210372 3168
rect 140037 3163 140103 3166
rect 210366 3164 210372 3166
rect 210436 3164 210442 3228
<< via3 >>
rect 280660 633388 280724 633452
rect 53052 630804 53116 630868
rect 54340 630668 54404 630732
rect 476068 619924 476132 619988
rect 488580 619924 488644 619988
rect 506612 619924 506676 619988
rect 430620 601700 430684 601764
rect 430804 597620 430868 597684
rect 430988 592180 431052 592244
rect 280660 542948 280724 543012
rect 299980 542540 300044 542604
rect 320588 541044 320652 541108
rect 430620 520100 430684 520164
rect 430804 518740 430868 518804
rect 320772 518604 320836 518668
rect 299980 517244 300044 517308
rect 430988 517244 431052 517308
rect 360884 485012 360948 485076
rect 363460 483652 363524 483716
rect 488580 483652 488644 483716
rect 364932 482156 364996 482220
rect 506612 480796 506676 480860
rect 365116 479708 365180 479772
rect 208900 479572 208964 479636
rect 206140 479436 206204 479500
rect 476068 479436 476132 479500
rect 55076 478756 55140 478820
rect 54892 478620 54956 478684
rect 198780 478892 198844 478956
rect 198228 478756 198292 478820
rect 360700 478756 360764 478820
rect 196572 478620 196636 478684
rect 206876 478620 206940 478684
rect 214788 478620 214852 478684
rect 371740 478620 371804 478684
rect 55444 478484 55508 478548
rect 54708 478348 54772 478412
rect 198044 478484 198108 478548
rect 205404 478484 205468 478548
rect 209268 478484 209332 478548
rect 367692 478484 367756 478548
rect 52316 478212 52380 478276
rect 200620 478348 200684 478412
rect 206508 478348 206572 478412
rect 370452 478348 370516 478412
rect 374500 478348 374564 478412
rect 197860 478212 197924 478276
rect 200988 478212 201052 478276
rect 219204 478212 219268 478276
rect 375972 478212 376036 478276
rect 46796 478076 46860 478140
rect 202092 478076 202156 478140
rect 213684 478076 213748 478140
rect 374684 478076 374748 478140
rect 59308 477940 59372 478004
rect 196756 477940 196820 478004
rect 202644 477940 202708 478004
rect 357940 477940 358004 478004
rect 358124 477804 358188 477868
rect 198596 477668 198660 477732
rect 201356 477668 201420 477732
rect 216996 477668 217060 477732
rect 50844 477592 50908 477596
rect 50844 477536 50894 477592
rect 50894 477536 50908 477592
rect 50844 477532 50908 477536
rect 53236 477532 53300 477596
rect 217548 477532 217612 477596
rect 219940 477532 220004 477596
rect 359412 476852 359476 476916
rect 209820 476716 209884 476780
rect 367876 476716 367940 476780
rect 57100 475764 57164 475828
rect 215340 475492 215404 475556
rect 371924 475492 371988 475556
rect 213316 474268 213380 474332
rect 377260 474268 377324 474332
rect 214420 474132 214484 474196
rect 363644 474132 363708 474196
rect 198964 473996 199028 474060
rect 210372 473996 210436 474060
rect 57284 472636 57348 472700
rect 217180 472636 217244 472700
rect 212028 472500 212092 472564
rect 379468 472500 379532 472564
rect 204852 471276 204916 471340
rect 215524 471140 215588 471204
rect 378732 471140 378796 471204
rect 206324 470052 206388 470116
rect 44772 469916 44836 469980
rect 211844 469916 211908 469980
rect 44956 469780 45020 469844
rect 212580 469780 212644 469844
rect 359596 469780 359660 469844
rect 210004 468692 210068 468756
rect 214604 468556 214668 468620
rect 211660 468420 211724 468484
rect 378916 468420 378980 468484
rect 207060 467196 207124 467260
rect 209084 467060 209148 467124
rect 203196 466108 203260 466172
rect 47900 465836 47964 465900
rect 377444 465836 377508 465900
rect 57836 465700 57900 465764
rect 376156 465700 376220 465764
rect 207980 464340 208044 464404
rect 52132 463388 52196 463452
rect 217364 463252 217428 463316
rect 203012 463116 203076 463180
rect 202276 462980 202340 463044
rect 47716 462844 47780 462908
rect 213132 462844 213196 462908
rect 376892 462844 376956 462908
rect 59124 461620 59188 461684
rect 179644 461620 179708 461684
rect 60228 461484 60292 461548
rect 359780 461484 359844 461548
rect 178356 461408 178420 461412
rect 178356 461352 178370 461408
rect 178370 461352 178420 461408
rect 178356 461348 178420 461352
rect 190868 461000 190932 461004
rect 190868 460944 190918 461000
rect 190918 460944 190932 461000
rect 190868 460940 190932 460944
rect 338252 461000 338316 461004
rect 338252 460944 338302 461000
rect 338302 460944 338316 461000
rect 338252 460940 338316 460944
rect 339724 461000 339788 461004
rect 339724 460944 339774 461000
rect 339774 460944 339788 461000
rect 339724 460940 339788 460944
rect 350948 461000 351012 461004
rect 350948 460944 350998 461000
rect 350998 460944 351012 461000
rect 350948 460940 351012 460944
rect 498516 460940 498580 461004
rect 499804 461000 499868 461004
rect 499804 460944 499854 461000
rect 499854 460944 499868 461000
rect 499804 460940 499868 460944
rect 510844 461000 510908 461004
rect 510844 460944 510894 461000
rect 510894 460944 510908 461000
rect 510844 460940 510908 460944
rect 48084 460804 48148 460868
rect 202460 460804 202524 460868
rect 46612 460668 46676 460732
rect 205220 460668 205284 460732
rect 55628 460532 55692 460596
rect 215892 460532 215956 460596
rect 51948 460396 52012 460460
rect 218652 460396 218716 460460
rect 51764 460260 51828 460324
rect 205036 460260 205100 460324
rect 359964 460260 360028 460324
rect 50660 460124 50724 460188
rect 218836 460124 218900 460188
rect 377628 460124 377692 460188
rect 53420 459988 53484 460052
rect 50476 459580 50540 459644
rect 53604 459580 53668 459644
rect 200804 459444 200868 459508
rect 58572 459036 58636 459100
rect 58940 458900 59004 458964
rect 379100 458900 379164 458964
rect 58756 458764 58820 458828
rect 199148 458764 199212 458828
rect 379284 458764 379348 458828
rect 205404 456860 205468 456924
rect 56548 415244 56612 415308
rect 56548 407764 56612 407828
rect 207060 407764 207124 407828
rect 358124 407764 358188 407828
rect 198780 394572 198844 394636
rect 199332 392124 199396 392188
rect 198780 391988 198844 392052
rect 199148 390628 199212 390692
rect 199148 388996 199212 389060
rect 198964 388452 199028 388516
rect 212028 382332 212092 382396
rect 51764 375260 51828 375324
rect 53236 375260 53300 375324
rect 55444 375320 55508 375324
rect 55444 375264 55494 375320
rect 55494 375264 55508 375320
rect 55444 375260 55508 375264
rect 200988 375260 201052 375324
rect 202644 375260 202708 375324
rect 206508 375260 206572 375324
rect 209820 375260 209884 375324
rect 211844 375260 211908 375324
rect 244780 375048 244844 375052
rect 244780 374992 244794 375048
rect 244794 374992 244844 375048
rect 244780 374988 244844 374992
rect 270540 375048 270604 375052
rect 270540 374992 270554 375048
rect 270554 374992 270604 375048
rect 270540 374988 270604 374992
rect 283052 375048 283116 375052
rect 283052 374992 283066 375048
rect 283066 374992 283116 375048
rect 283052 374988 283116 374992
rect 315252 374988 315316 375052
rect 407804 375048 407868 375052
rect 407804 374992 407818 375048
rect 407818 374992 407868 375048
rect 407804 374988 407868 374992
rect 425100 375048 425164 375052
rect 425100 374992 425114 375048
rect 425114 374992 425164 375048
rect 425100 374988 425164 374992
rect 440372 375048 440436 375052
rect 440372 374992 440386 375048
rect 440386 374992 440436 375048
rect 440372 374988 440436 374992
rect 443132 375048 443196 375052
rect 443132 374992 443146 375048
rect 443146 374992 443196 375048
rect 443132 374988 443196 374992
rect 404214 374776 404278 374780
rect 404214 374720 404230 374776
rect 404230 374720 404278 374776
rect 404214 374716 404278 374720
rect 158484 374640 158548 374644
rect 158484 374584 158534 374640
rect 158534 374584 158548 374640
rect 158484 374580 158548 374584
rect 165950 374640 166014 374644
rect 165950 374584 165986 374640
rect 165986 374584 166014 374640
rect 165950 374580 166014 374584
rect 320918 374640 320982 374644
rect 320918 374584 320970 374640
rect 320970 374584 320982 374640
rect 320918 374580 320982 374584
rect 359964 374580 360028 374644
rect 410742 374640 410806 374644
rect 410742 374584 410762 374640
rect 410762 374584 410806 374640
rect 105492 374504 105556 374508
rect 105492 374448 105506 374504
rect 105506 374448 105556 374504
rect 105492 374444 105556 374448
rect 116038 374504 116102 374508
rect 116038 374448 116086 374504
rect 116086 374448 116102 374504
rect 116038 374444 116102 374448
rect 140926 374504 140990 374508
rect 140926 374448 140962 374504
rect 140962 374448 140990 374504
rect 140926 374444 140990 374448
rect 143510 374504 143574 374508
rect 143510 374448 143538 374504
rect 143538 374448 143574 374504
rect 143510 374444 143574 374448
rect 156460 374504 156524 374508
rect 156460 374448 156510 374504
rect 156510 374448 156524 374504
rect 156460 374444 156524 374448
rect 160918 374504 160982 374508
rect 160918 374448 160926 374504
rect 160926 374448 160982 374504
rect 160918 374444 160982 374448
rect 163366 374504 163430 374508
rect 163366 374448 163410 374504
rect 163410 374448 163430 374504
rect 163366 374444 163430 374448
rect 244228 374504 244292 374508
rect 244228 374448 244278 374504
rect 244278 374448 244292 374504
rect 244228 374444 244292 374448
rect 247614 374504 247678 374508
rect 247614 374448 247646 374504
rect 247646 374448 247678 374504
rect 247614 374444 247678 374448
rect 253462 374504 253526 374508
rect 253462 374448 253478 374504
rect 253478 374448 253526 374504
rect 253462 374444 253526 374448
rect 265294 374504 265358 374508
rect 265294 374448 265310 374504
rect 265310 374448 265358 374504
rect 265294 374444 265358 374448
rect 146156 374368 146220 374372
rect 146156 374312 146206 374368
rect 146206 374312 146220 374368
rect 146156 374308 146220 374312
rect 148916 374368 148980 374372
rect 148916 374312 148966 374368
rect 148966 374312 148980 374368
rect 148916 374308 148980 374312
rect 262260 374308 262324 374372
rect 273852 374172 273916 374236
rect 139164 374096 139228 374100
rect 139164 374040 139214 374096
rect 139214 374040 139228 374096
rect 139164 374036 139228 374040
rect 271276 374036 271340 374100
rect 410742 374580 410806 374584
rect 450998 374640 451062 374644
rect 450998 374584 451002 374640
rect 451002 374584 451058 374640
rect 451058 374584 451062 374640
rect 450998 374580 451062 374584
rect 433590 374504 433654 374508
rect 433590 374448 433614 374504
rect 433614 374448 433654 374504
rect 433590 374444 433654 374448
rect 436038 374504 436102 374508
rect 436038 374448 436062 374504
rect 436062 374448 436102 374504
rect 436038 374444 436102 374448
rect 438486 374504 438550 374508
rect 438486 374448 438490 374504
rect 438490 374448 438546 374504
rect 438546 374448 438550 374504
rect 438486 374444 438550 374448
rect 429148 374036 429212 374100
rect 199148 373900 199212 373964
rect 279188 373900 279252 373964
rect 377628 373900 377692 373964
rect 475332 373900 475396 373964
rect 199332 373764 199396 373828
rect 258028 373824 258092 373828
rect 258028 373768 258078 373824
rect 258078 373768 258092 373824
rect 258028 373764 258092 373768
rect 268516 373764 268580 373828
rect 416084 373824 416148 373828
rect 416084 373768 416098 373824
rect 416098 373768 416148 373824
rect 416084 373764 416148 373768
rect 421052 373824 421116 373828
rect 421052 373768 421066 373824
rect 421066 373768 421116 373824
rect 421052 373764 421116 373768
rect 423076 373824 423140 373828
rect 423076 373768 423090 373824
rect 423090 373768 423140 373824
rect 423076 373764 423140 373768
rect 426940 373824 427004 373828
rect 426940 373768 426954 373824
rect 426954 373768 427004 373824
rect 426940 373764 427004 373768
rect 430620 373824 430684 373828
rect 430620 373768 430634 373824
rect 430634 373768 430684 373824
rect 430620 373764 430684 373768
rect 95004 373688 95068 373692
rect 95004 373632 95054 373688
rect 95054 373632 95068 373688
rect 95004 373628 95068 373632
rect 96108 373688 96172 373692
rect 96108 373632 96122 373688
rect 96122 373632 96172 373688
rect 96108 373628 96172 373632
rect 103284 373628 103348 373692
rect 107884 373688 107948 373692
rect 107884 373632 107898 373688
rect 107898 373632 107948 373688
rect 107884 373628 107948 373632
rect 113588 373688 113652 373692
rect 113588 373632 113602 373688
rect 113602 373632 113652 373688
rect 113588 373628 113652 373632
rect 118372 373688 118436 373692
rect 118372 373632 118386 373688
rect 118386 373632 118436 373688
rect 118372 373628 118436 373632
rect 121316 373688 121380 373692
rect 121316 373632 121366 373688
rect 121366 373632 121380 373688
rect 121316 373628 121380 373632
rect 110460 373552 110524 373556
rect 110460 373496 110474 373552
rect 110474 373496 110524 373552
rect 110460 373492 110524 373496
rect 119844 373492 119908 373556
rect 217548 373628 217612 373692
rect 266308 373628 266372 373692
rect 445892 373688 445956 373692
rect 445892 373632 445906 373688
rect 445906 373632 445956 373688
rect 445892 373628 445956 373632
rect 455460 373688 455524 373692
rect 455460 373632 455474 373688
rect 455474 373632 455524 373688
rect 455460 373628 455524 373632
rect 124076 373552 124140 373556
rect 124076 373496 124126 373552
rect 124126 373496 124140 373552
rect 124076 373492 124140 373496
rect 125732 373552 125796 373556
rect 125732 373496 125746 373552
rect 125746 373496 125796 373552
rect 125732 373492 125796 373496
rect 128860 373552 128924 373556
rect 128860 373496 128910 373552
rect 128910 373496 128924 373552
rect 128860 373492 128924 373496
rect 131068 373552 131132 373556
rect 131068 373496 131082 373552
rect 131082 373496 131132 373552
rect 131068 373492 131132 373496
rect 133644 373552 133708 373556
rect 133644 373496 133694 373552
rect 133694 373496 133708 373552
rect 133644 373492 133708 373496
rect 136404 373552 136468 373556
rect 136404 373496 136454 373552
rect 136454 373496 136468 373552
rect 136404 373492 136468 373496
rect 151676 373552 151740 373556
rect 151676 373496 151726 373552
rect 151726 373496 151740 373552
rect 151676 373492 151740 373496
rect 154068 373552 154132 373556
rect 154068 373496 154118 373552
rect 154118 373496 154132 373552
rect 154068 373492 154132 373496
rect 263732 373552 263796 373556
rect 263732 373496 263746 373552
rect 263746 373496 263796 373552
rect 263732 373492 263796 373496
rect 447732 373552 447796 373556
rect 447732 373496 447746 373552
rect 447746 373496 447796 373552
rect 447732 373492 447796 373496
rect 458220 373552 458284 373556
rect 458220 373496 458234 373552
rect 458234 373496 458284 373552
rect 458220 373492 458284 373496
rect 93716 373416 93780 373420
rect 93716 373360 93730 373416
rect 93730 373360 93780 373416
rect 93716 373356 93780 373360
rect 98316 373416 98380 373420
rect 98316 373360 98330 373416
rect 98330 373360 98380 373416
rect 98316 373356 98380 373360
rect 269252 373416 269316 373420
rect 269252 373360 269266 373416
rect 269266 373360 269316 373416
rect 269252 373356 269316 373360
rect 452884 373416 452948 373420
rect 452884 373360 452898 373416
rect 452898 373360 452948 373416
rect 452884 373356 452948 373360
rect 485820 373416 485884 373420
rect 485820 373360 485834 373416
rect 485834 373360 485884 373416
rect 485820 373356 485884 373360
rect 88380 373280 88444 373284
rect 88380 373224 88394 373280
rect 88394 373224 88444 373280
rect 88380 373220 88444 373224
rect 95924 373280 95988 373284
rect 95924 373224 95974 373280
rect 95974 373224 95988 373280
rect 95924 373220 95988 373224
rect 100892 373280 100956 373284
rect 100892 373224 100906 373280
rect 100906 373224 100956 373280
rect 100892 373220 100956 373224
rect 242940 373280 243004 373284
rect 242940 373224 242954 373280
rect 242954 373224 243004 373280
rect 242940 373220 243004 373224
rect 261340 373280 261404 373284
rect 261340 373224 261354 373280
rect 261354 373224 261404 373280
rect 261340 373220 261404 373224
rect 279188 373220 279252 373284
rect 90220 373144 90284 373148
rect 90220 373088 90234 373144
rect 90234 373088 90284 373144
rect 90220 373084 90284 373088
rect 92428 373144 92492 373148
rect 92428 373088 92442 373144
rect 92442 373088 92492 373144
rect 92428 373084 92492 373088
rect 235948 373144 236012 373148
rect 235948 373088 235998 373144
rect 235998 373088 236012 373144
rect 235948 373084 236012 373088
rect 253980 373144 254044 373148
rect 253980 373088 253994 373144
rect 253994 373088 254044 373144
rect 253980 373084 254044 373088
rect 255452 373144 255516 373148
rect 255452 373088 255466 373144
rect 255466 373088 255516 373144
rect 255452 373084 255516 373088
rect 272012 373144 272076 373148
rect 272012 373088 272026 373144
rect 272026 373088 272076 373144
rect 272012 373084 272076 373088
rect 300900 373144 300964 373148
rect 300900 373088 300914 373144
rect 300914 373088 300964 373144
rect 300900 373084 300964 373088
rect 57100 372812 57164 372876
rect 57284 372676 57348 372740
rect 199148 372676 199212 372740
rect 210004 372676 210068 372740
rect 216996 372736 217060 372740
rect 216996 372680 217046 372736
rect 217046 372680 217060 372736
rect 216996 372676 217060 372680
rect 77156 372600 77220 372604
rect 77156 372544 77206 372600
rect 77206 372544 77220 372600
rect 77156 372540 77220 372544
rect 84516 372540 84580 372604
rect 86540 372600 86604 372604
rect 86540 372544 86590 372600
rect 86590 372544 86604 372600
rect 86540 372540 86604 372544
rect 88012 372600 88076 372604
rect 88012 372544 88062 372600
rect 88062 372544 88076 372600
rect 88012 372540 88076 372544
rect 89300 372600 89364 372604
rect 89300 372544 89350 372600
rect 89350 372544 89364 372600
rect 89300 372540 89364 372544
rect 90036 372600 90100 372604
rect 90036 372544 90086 372600
rect 90086 372544 90100 372600
rect 90036 372540 90100 372544
rect 91508 372540 91572 372604
rect 93348 372540 93412 372604
rect 108804 372600 108868 372604
rect 108804 372544 108854 372600
rect 108854 372544 108868 372600
rect 108804 372540 108868 372544
rect 113220 372540 113284 372604
rect 183140 372600 183204 372604
rect 183140 372544 183190 372600
rect 183190 372544 183204 372600
rect 183140 372540 183204 372544
rect 236500 372540 236564 372604
rect 238156 372600 238220 372604
rect 238156 372544 238170 372600
rect 238170 372544 238220 372600
rect 238156 372540 238220 372544
rect 239260 372600 239324 372604
rect 239260 372544 239310 372600
rect 239310 372544 239324 372600
rect 239260 372540 239324 372544
rect 240364 372600 240428 372604
rect 240364 372544 240414 372600
rect 240414 372544 240428 372600
rect 240364 372540 240428 372544
rect 241468 372600 241532 372604
rect 241468 372544 241518 372600
rect 241518 372544 241532 372600
rect 241468 372540 241532 372544
rect 245884 372540 245948 372604
rect 248460 372600 248524 372604
rect 248460 372544 248474 372600
rect 248474 372544 248524 372600
rect 248460 372540 248524 372544
rect 251220 372600 251284 372604
rect 251220 372544 251234 372600
rect 251234 372544 251284 372600
rect 251220 372540 251284 372544
rect 256740 372600 256804 372604
rect 256740 372544 256754 372600
rect 256754 372544 256804 372600
rect 256740 372540 256804 372544
rect 259500 372600 259564 372604
rect 259500 372544 259514 372600
rect 259514 372544 259564 372600
rect 259500 372540 259564 372544
rect 260052 372540 260116 372604
rect 273300 372600 273364 372604
rect 273300 372544 273314 372600
rect 273314 372544 273364 372600
rect 273300 372540 273364 372544
rect 310652 372540 310716 372604
rect 313412 372540 313476 372604
rect 78444 372464 78508 372468
rect 78444 372408 78494 372464
rect 78494 372408 78508 372464
rect 78444 372404 78508 372408
rect 79916 372464 79980 372468
rect 79916 372408 79966 372464
rect 79966 372408 79980 372464
rect 79916 372404 79980 372408
rect 84700 372404 84764 372468
rect 102732 372464 102796 372468
rect 102732 372408 102782 372464
rect 102782 372408 102796 372464
rect 102732 372404 102796 372408
rect 117084 372404 117148 372468
rect 277164 372404 277228 372468
rect 305316 372404 305380 372468
rect 376892 372676 376956 372740
rect 408540 372600 408604 372604
rect 408540 372544 408554 372600
rect 408554 372544 408604 372600
rect 408540 372540 408604 372544
rect 426388 372600 426452 372604
rect 426388 372544 426438 372600
rect 426438 372544 426452 372600
rect 426388 372540 426452 372544
rect 433564 372540 433628 372604
rect 438348 372540 438412 372604
rect 431172 372404 431236 372468
rect 80468 372328 80532 372332
rect 80468 372272 80518 372328
rect 80518 372272 80532 372328
rect 80468 372268 80532 372272
rect 81940 372328 82004 372332
rect 81940 372272 81954 372328
rect 81954 372272 82004 372328
rect 81940 372268 82004 372272
rect 101996 372328 102060 372332
rect 101996 372272 102046 372328
rect 102046 372272 102060 372328
rect 101996 372268 102060 372272
rect 109540 372268 109604 372332
rect 118188 372268 118252 372332
rect 277532 372268 277596 372332
rect 470732 372268 470796 372332
rect 76604 372132 76668 372196
rect 111748 372132 111812 372196
rect 404860 372132 404924 372196
rect 503116 372192 503180 372196
rect 503116 372136 503166 372192
rect 503166 372136 503180 372192
rect 503116 372132 503180 372136
rect 503484 372192 503548 372196
rect 503484 372136 503534 372192
rect 503534 372136 503548 372192
rect 503484 372132 503548 372136
rect 83780 371920 83844 371924
rect 83780 371864 83830 371920
rect 83830 371864 83844 371920
rect 83780 371860 83844 371864
rect 104572 371920 104636 371924
rect 104572 371864 104622 371920
rect 104622 371864 104636 371920
rect 104572 371860 104636 371864
rect 112852 371860 112916 371924
rect 105308 371724 105372 371788
rect 114508 371724 114572 371788
rect 396212 371996 396276 372060
rect 397500 372056 397564 372060
rect 397500 372000 397514 372056
rect 397514 372000 397564 372056
rect 397500 371996 397564 372000
rect 398972 371996 399036 372060
rect 400260 372056 400324 372060
rect 400260 372000 400274 372056
rect 400274 372000 400324 372056
rect 400260 371996 400324 372000
rect 410012 371996 410076 372060
rect 97580 371588 97644 371652
rect 98132 371588 98196 371652
rect 99972 371588 100036 371652
rect 377444 371860 377508 371924
rect 433380 371860 433444 371924
rect 275324 371784 275388 371788
rect 275324 371728 275374 371784
rect 275374 371728 275388 371784
rect 275324 371724 275388 371728
rect 317828 371724 317892 371788
rect 439452 371724 439516 371788
rect 247908 371588 247972 371652
rect 250300 371588 250364 371652
rect 251956 371588 252020 371652
rect 326660 371588 326724 371652
rect 402284 371588 402348 371652
rect 411300 371648 411364 371652
rect 411300 371592 411314 371648
rect 411314 371592 411364 371648
rect 411300 371588 411364 371592
rect 418844 371588 418908 371652
rect 423996 371588 424060 371652
rect 427860 371648 427924 371652
rect 427860 371592 427874 371648
rect 427874 371592 427924 371648
rect 427860 371588 427924 371592
rect 462636 371588 462700 371652
rect 465396 371588 465460 371652
rect 478092 371588 478156 371652
rect 100708 371452 100772 371516
rect 183324 371452 183388 371516
rect 265756 371452 265820 371516
rect 273668 371452 273732 371516
rect 407252 371452 407316 371516
rect 411852 371452 411916 371516
rect 418108 371452 418172 371516
rect 421236 371452 421300 371516
rect 480300 371512 480364 371516
rect 480300 371456 480314 371512
rect 480314 371456 480364 371512
rect 480300 371452 480364 371456
rect 106964 371316 107028 371380
rect 107516 371376 107580 371380
rect 107516 371320 107566 371376
rect 107566 371320 107580 371376
rect 107516 371316 107580 371320
rect 115796 371316 115860 371380
rect 249932 371316 249996 371380
rect 253612 371316 253676 371380
rect 256188 371316 256252 371380
rect 258396 371316 258460 371380
rect 260972 371316 261036 371380
rect 263548 371376 263612 371380
rect 263548 371320 263598 371376
rect 263598 371320 263612 371376
rect 263548 371316 263612 371320
rect 267044 371316 267108 371380
rect 267780 371376 267844 371380
rect 267780 371320 267794 371376
rect 267794 371320 267844 371376
rect 267780 371316 267844 371320
rect 276244 371316 276308 371380
rect 278268 371316 278332 371380
rect 280292 371316 280356 371380
rect 285812 371316 285876 371380
rect 287652 371316 287716 371380
rect 290596 371316 290660 371380
rect 292804 371316 292868 371380
rect 295380 371376 295444 371380
rect 295380 371320 295394 371376
rect 295394 371320 295444 371376
rect 295380 371316 295444 371320
rect 298140 371376 298204 371380
rect 298140 371320 298154 371376
rect 298154 371320 298204 371376
rect 298140 371316 298204 371320
rect 302924 371316 302988 371380
rect 308628 371316 308692 371380
rect 322980 371376 323044 371380
rect 322980 371320 322994 371376
rect 322994 371320 323044 371376
rect 322980 371316 323044 371320
rect 343220 371316 343284 371380
rect 343404 371376 343468 371380
rect 343404 371320 343454 371376
rect 343454 371320 343468 371376
rect 343404 371316 343468 371320
rect 396580 371316 396644 371380
rect 403020 371376 403084 371380
rect 403020 371320 403034 371376
rect 403034 371320 403084 371376
rect 403020 371316 403084 371320
rect 406148 371316 406212 371380
rect 412772 371316 412836 371380
rect 413692 371316 413756 371380
rect 414060 371376 414124 371380
rect 414060 371320 414074 371376
rect 414074 371320 414124 371376
rect 414060 371316 414124 371320
rect 415532 371316 415596 371380
rect 416820 371376 416884 371380
rect 416820 371320 416834 371376
rect 416834 371320 416884 371376
rect 416820 371316 416884 371320
rect 418292 371316 418356 371380
rect 420316 371316 420380 371380
rect 422340 371376 422404 371380
rect 422340 371320 422354 371376
rect 422354 371320 422404 371376
rect 422340 371316 422404 371320
rect 425652 371316 425716 371380
rect 428596 371316 428660 371380
rect 432092 371316 432156 371380
rect 434852 371316 434916 371380
rect 436324 371316 436388 371380
rect 460980 371376 461044 371380
rect 460980 371320 460994 371376
rect 460994 371320 461044 371376
rect 460980 371316 461044 371320
rect 467972 371316 468036 371380
rect 473308 371376 473372 371380
rect 473308 371320 473358 371376
rect 473358 371320 473372 371376
rect 473308 371316 473372 371320
rect 483244 371316 483308 371380
rect 216996 370908 217060 370972
rect 217548 370908 217612 370972
rect 214788 369820 214852 369884
rect 209268 369140 209332 369204
rect 212580 369140 212644 369204
rect 376892 368520 376956 368524
rect 376892 368464 376942 368520
rect 376942 368464 376956 368520
rect 376892 368460 376956 368464
rect 179644 355268 179708 355332
rect 190868 355268 190932 355332
rect 339724 354996 339788 355060
rect 350948 354996 351012 355060
rect 498516 354996 498580 355060
rect 499804 354860 499868 354924
rect 178540 354784 178604 354788
rect 178540 354728 178590 354784
rect 178590 354728 178604 354784
rect 178540 354724 178604 354728
rect 338068 354784 338132 354788
rect 338068 354728 338118 354784
rect 338118 354728 338132 354784
rect 338068 354724 338132 354728
rect 510844 354784 510908 354788
rect 510844 354728 510894 354784
rect 510894 354728 510908 354784
rect 510844 354724 510908 354728
rect 54340 304948 54404 305012
rect 359780 279924 359844 279988
rect 111006 269920 111070 269924
rect 111006 269864 111026 269920
rect 111026 269864 111070 269920
rect 111006 269860 111070 269864
rect 148542 269920 148606 269924
rect 148542 269864 148562 269920
rect 148562 269864 148606 269920
rect 148542 269860 148606 269864
rect 133446 269784 133510 269788
rect 133446 269728 133474 269784
rect 133474 269728 133510 269784
rect 133446 269724 133510 269728
rect 135894 269784 135958 269788
rect 135894 269728 135902 269784
rect 135902 269728 135958 269784
rect 135894 269724 135958 269728
rect 138478 269784 138542 269788
rect 138478 269728 138534 269784
rect 138534 269728 138542 269784
rect 138478 269724 138542 269728
rect 140926 269724 140990 269788
rect 250742 269784 250806 269788
rect 250742 269728 250774 269784
rect 250774 269728 250806 269784
rect 250742 269724 250806 269728
rect 416046 269784 416110 269788
rect 416046 269728 416098 269784
rect 416098 269728 416110 269784
rect 416046 269724 416110 269728
rect 425294 269784 425358 269788
rect 425294 269728 425298 269784
rect 425298 269728 425358 269784
rect 425294 269724 425358 269728
rect 433318 269784 433382 269788
rect 433318 269728 433338 269784
rect 433338 269728 433382 269784
rect 433318 269724 433382 269728
rect 434406 269724 434470 269788
rect 83126 269648 83190 269652
rect 83126 269592 83150 269648
rect 83150 269592 83190 269648
rect 83126 269588 83190 269592
rect 91286 269648 91350 269652
rect 91286 269592 91338 269648
rect 91338 269592 91350 269648
rect 91286 269588 91350 269592
rect 93598 269648 93662 269652
rect 93598 269592 93638 269648
rect 93638 269592 93662 269648
rect 93598 269588 93662 269592
rect 94550 269648 94614 269652
rect 94550 269592 94558 269648
rect 94558 269592 94614 269648
rect 94550 269588 94614 269592
rect 143510 269648 143574 269652
rect 143510 269592 143538 269648
rect 143538 269592 143574 269648
rect 143510 269588 143574 269592
rect 145958 269648 146022 269652
rect 145958 269592 145986 269648
rect 145986 269592 146022 269648
rect 145958 269588 146022 269592
rect 283518 269648 283582 269652
rect 283518 269592 283526 269648
rect 283526 269592 283582 269648
rect 283518 269588 283582 269592
rect 288278 269648 288342 269652
rect 288278 269592 288310 269648
rect 288310 269592 288342 269648
rect 288278 269588 288342 269592
rect 290998 269648 291062 269652
rect 290998 269592 291014 269648
rect 291014 269592 291062 269648
rect 290998 269588 291062 269592
rect 293446 269648 293510 269652
rect 293446 269592 293462 269648
rect 293462 269592 293510 269648
rect 293446 269588 293510 269592
rect 305958 269648 306022 269652
rect 305958 269592 305974 269648
rect 305974 269592 306022 269648
rect 305958 269588 306022 269592
rect 318470 269648 318534 269652
rect 318470 269592 318486 269648
rect 318486 269592 318534 269648
rect 318470 269588 318534 269592
rect 429782 269648 429846 269652
rect 429782 269592 429806 269648
rect 429806 269592 429846 269648
rect 429782 269588 429846 269592
rect 436038 269648 436102 269652
rect 436038 269592 436062 269648
rect 436062 269592 436102 269648
rect 436038 269588 436102 269592
rect 468542 269588 468606 269652
rect 470990 269648 471054 269652
rect 470990 269592 471022 269648
rect 471022 269592 471054 269648
rect 470990 269588 471054 269592
rect 480918 269648 480982 269652
rect 480918 269592 480958 269648
rect 480958 269592 480982 269648
rect 480918 269588 480982 269592
rect 376892 269316 376956 269380
rect 377996 269316 378060 269380
rect 359596 269180 359660 269244
rect 473492 269180 473556 269244
rect 115796 269044 115860 269108
rect 196756 269044 196820 269108
rect 311020 269044 311084 269108
rect 323348 269104 323412 269108
rect 323348 269048 323362 269104
rect 323362 269048 323412 269104
rect 323348 269044 323412 269048
rect 486004 269044 486068 269108
rect 116900 268908 116964 268972
rect 217364 268908 217428 268972
rect 320956 268908 321020 268972
rect 359412 268908 359476 268972
rect 76052 268832 76116 268836
rect 76052 268776 76066 268832
rect 76066 268776 76116 268832
rect 76052 268772 76116 268776
rect 77156 268832 77220 268836
rect 77156 268776 77170 268832
rect 77170 268776 77220 268832
rect 77156 268772 77220 268776
rect 90772 268832 90836 268836
rect 90772 268776 90786 268832
rect 90786 268776 90836 268832
rect 90772 268772 90836 268776
rect 95924 268832 95988 268836
rect 95924 268776 95938 268832
rect 95938 268776 95988 268832
rect 95924 268772 95988 268776
rect 96108 268832 96172 268836
rect 96108 268776 96122 268832
rect 96122 268776 96172 268832
rect 96108 268772 96172 268776
rect 98500 268832 98564 268836
rect 98500 268776 98514 268832
rect 98514 268776 98564 268832
rect 98500 268772 98564 268776
rect 99420 268832 99484 268836
rect 99420 268776 99434 268832
rect 99434 268776 99484 268832
rect 99420 268772 99484 268776
rect 100708 268832 100772 268836
rect 100708 268776 100758 268832
rect 100758 268776 100772 268832
rect 100708 268772 100772 268776
rect 106412 268832 106476 268836
rect 106412 268776 106426 268832
rect 106426 268776 106476 268832
rect 106412 268772 106476 268776
rect 217548 268772 217612 268836
rect 243124 268832 243188 268836
rect 243124 268776 243138 268832
rect 243138 268776 243188 268832
rect 243124 268772 243188 268776
rect 257844 268772 257908 268836
rect 261708 268832 261772 268836
rect 261708 268776 261722 268832
rect 261722 268776 261772 268832
rect 261708 268772 261772 268776
rect 295932 268832 295996 268836
rect 295932 268776 295946 268832
rect 295946 268776 295996 268832
rect 295932 268772 295996 268776
rect 298508 268832 298572 268836
rect 298508 268776 298522 268832
rect 298522 268776 298572 268832
rect 298508 268772 298572 268776
rect 300900 268832 300964 268836
rect 300900 268776 300914 268832
rect 300914 268776 300964 268832
rect 300900 268772 300964 268776
rect 303476 268832 303540 268836
rect 303476 268776 303490 268832
rect 303490 268776 303540 268832
rect 303476 268772 303540 268776
rect 377996 268772 378060 268836
rect 417004 268832 417068 268836
rect 417004 268776 417018 268832
rect 417018 268776 417068 268832
rect 417004 268772 417068 268776
rect 421052 268832 421116 268836
rect 422892 268968 422956 268972
rect 422892 268912 422906 268968
rect 422906 268912 422956 268968
rect 422892 268908 422956 268912
rect 426020 268968 426084 268972
rect 426020 268912 426034 268968
rect 426034 268912 426084 268968
rect 426020 268908 426084 268912
rect 430988 268968 431052 268972
rect 430988 268912 431002 268968
rect 431002 268912 431052 268968
rect 430988 268908 431052 268912
rect 432276 268968 432340 268972
rect 432276 268912 432290 268968
rect 432290 268912 432340 268968
rect 432276 268908 432340 268912
rect 475884 268968 475948 268972
rect 475884 268912 475898 268968
rect 475898 268912 475948 268968
rect 475884 268908 475948 268912
rect 478460 268968 478524 268972
rect 478460 268912 478474 268968
rect 478474 268912 478524 268968
rect 478460 268908 478524 268912
rect 483428 268968 483492 268972
rect 483428 268912 483442 268968
rect 483442 268912 483492 268968
rect 483428 268908 483492 268912
rect 421052 268776 421066 268832
rect 421066 268776 421116 268832
rect 421052 268772 421116 268776
rect 423444 268772 423508 268836
rect 423996 268636 424060 268700
rect 101812 268500 101876 268564
rect 103836 268364 103900 268428
rect 85436 268152 85500 268156
rect 85436 268096 85450 268152
rect 85450 268096 85500 268152
rect 85436 268092 85500 268096
rect 92428 268152 92492 268156
rect 92428 268096 92442 268152
rect 92442 268096 92492 268152
rect 92428 268092 92492 268096
rect 103284 268092 103348 268156
rect 113588 268152 113652 268156
rect 113588 268096 113602 268152
rect 113602 268096 113652 268152
rect 113588 268092 113652 268096
rect 128308 268152 128372 268156
rect 128308 268096 128358 268152
rect 128358 268096 128372 268152
rect 128308 268092 128372 268096
rect 265204 268152 265268 268156
rect 265204 268096 265218 268152
rect 265218 268096 265268 268152
rect 265204 268092 265268 268096
rect 275876 268152 275940 268156
rect 275876 268096 275926 268152
rect 275926 268096 275940 268152
rect 275876 268092 275940 268096
rect 398236 268152 398300 268156
rect 398236 268096 398250 268152
rect 398250 268096 398300 268152
rect 398236 268092 398300 268096
rect 401732 268152 401796 268156
rect 401732 268096 401746 268152
rect 401746 268096 401796 268152
rect 401732 268092 401796 268096
rect 455828 268152 455892 268156
rect 455828 268096 455842 268152
rect 455842 268096 455892 268152
rect 455828 268092 455892 268096
rect 463556 268092 463620 268156
rect 217548 267956 217612 268020
rect 216996 267820 217060 267884
rect 83964 267684 84028 267748
rect 97028 267744 97092 267748
rect 97028 267688 97042 267744
rect 97042 267688 97092 267744
rect 97028 267684 97092 267688
rect 98132 267684 98196 267748
rect 102732 267744 102796 267748
rect 102732 267688 102746 267744
rect 102746 267688 102796 267744
rect 102732 267684 102796 267688
rect 111196 267744 111260 267748
rect 111196 267688 111246 267744
rect 111246 267688 111260 267744
rect 111196 267684 111260 267688
rect 112300 267744 112364 267748
rect 112300 267688 112350 267744
rect 112350 267688 112364 267744
rect 112300 267684 112364 267688
rect 119108 267744 119172 267748
rect 119108 267688 119122 267744
rect 119122 267688 119172 267744
rect 119108 267684 119172 267688
rect 120764 267684 120828 267748
rect 125916 267684 125980 267748
rect 150940 267744 151004 267748
rect 150940 267688 150990 267744
rect 150990 267688 151004 267744
rect 150940 267684 151004 267688
rect 158484 267744 158548 267748
rect 158484 267688 158534 267744
rect 158534 267688 158548 267744
rect 158484 267684 158548 267688
rect 163452 267744 163516 267748
rect 163452 267688 163502 267744
rect 163502 267688 163516 267744
rect 163452 267684 163516 267688
rect 255820 267684 255884 267748
rect 258396 267684 258460 267748
rect 260972 267684 261036 267748
rect 263548 267744 263612 267748
rect 263548 267688 263598 267744
rect 263598 267688 263612 267744
rect 263548 267684 263612 267688
rect 265940 267684 266004 267748
rect 268332 267684 268396 267748
rect 270908 267684 270972 267748
rect 273484 267684 273548 267748
rect 276244 267684 276308 267748
rect 276980 267744 277044 267748
rect 276980 267688 277030 267744
rect 277030 267688 277044 267744
rect 276980 267684 277044 267688
rect 278084 267744 278148 267748
rect 278084 267688 278134 267744
rect 278134 267688 278148 267744
rect 278084 267684 278148 267688
rect 280844 267684 280908 267748
rect 403020 267744 403084 267748
rect 403020 267688 403034 267744
rect 403034 267688 403084 267744
rect 403020 267684 403084 267688
rect 414428 267744 414492 267748
rect 414428 267688 414442 267744
rect 414442 267688 414492 267744
rect 414428 267684 414492 267688
rect 415532 267684 415596 267748
rect 428596 267744 428660 267748
rect 428596 267688 428646 267744
rect 428646 267688 428660 267744
rect 428596 267684 428660 267688
rect 435588 267684 435652 267748
rect 451044 267684 451108 267748
rect 453436 267684 453500 267748
rect 458404 267684 458468 267748
rect 460980 267744 461044 267748
rect 460980 267688 460994 267744
rect 460994 267688 461044 267744
rect 460980 267684 461044 267688
rect 57836 267548 57900 267612
rect 123524 267548 123588 267612
rect 130884 267548 130948 267612
rect 155908 267608 155972 267612
rect 155908 267552 155958 267608
rect 155958 267552 155972 267608
rect 155908 267548 155972 267552
rect 160876 267608 160940 267612
rect 160876 267552 160926 267608
rect 160926 267552 160940 267608
rect 160876 267548 160940 267552
rect 80468 267412 80532 267476
rect 115980 267472 116044 267476
rect 115980 267416 115994 267472
rect 115994 267416 116044 267472
rect 115980 267412 116044 267416
rect 118372 267412 118436 267476
rect 154068 267412 154132 267476
rect 198780 267548 198844 267612
rect 315988 267548 316052 267612
rect 313412 267412 313476 267476
rect 343220 267412 343284 267476
rect 379468 267412 379532 267476
rect 428228 267412 428292 267476
rect 443500 267412 443564 267476
rect 503116 267472 503180 267476
rect 503116 267416 503166 267472
rect 503166 267416 503180 267472
rect 503116 267412 503180 267416
rect 503484 267472 503548 267476
rect 503484 267416 503534 267472
rect 503534 267416 503548 267472
rect 503484 267412 503548 267416
rect 81940 267276 82004 267340
rect 108252 267276 108316 267340
rect 183140 267276 183204 267340
rect 308628 267276 308692 267340
rect 377260 267276 377324 267340
rect 408172 267276 408236 267340
rect 439268 267276 439332 267340
rect 440924 267276 440988 267340
rect 448284 267276 448348 267340
rect 105860 267140 105924 267204
rect 217180 267140 217244 267204
rect 278452 267140 278516 267204
rect 279004 267140 279068 267204
rect 397132 267140 397196 267204
rect 418476 267140 418540 267204
rect 438532 267140 438596 267204
rect 445892 267140 445956 267204
rect 78260 267004 78324 267068
rect 79548 267004 79612 267068
rect 88380 267064 88444 267068
rect 88380 267008 88394 267064
rect 88394 267008 88444 267064
rect 88380 267004 88444 267008
rect 101076 267004 101140 267068
rect 109540 267004 109604 267068
rect 183508 267064 183572 267068
rect 183508 267008 183522 267064
rect 183522 267008 183572 267064
rect 183508 267004 183572 267008
rect 236500 267004 236564 267068
rect 256188 267004 256252 267068
rect 273300 267064 273364 267068
rect 273300 267008 273314 267064
rect 273314 267008 273364 267064
rect 273300 267004 273364 267008
rect 343404 267064 343468 267068
rect 343404 267008 343454 267064
rect 343454 267008 343468 267064
rect 343404 267004 343468 267008
rect 410748 267004 410812 267068
rect 413692 267004 413756 267068
rect 433564 267004 433628 267068
rect 165844 266868 165908 266932
rect 237052 266868 237116 266932
rect 248276 266868 248340 266932
rect 253612 266868 253676 266932
rect 285996 266868 286060 266932
rect 465948 266868 466012 266932
rect 326660 266732 326724 266796
rect 113220 266596 113284 266660
rect 118004 266596 118068 266660
rect 250116 266596 250180 266660
rect 408724 266596 408788 266660
rect 438348 266596 438412 266660
rect 105308 266460 105372 266524
rect 215340 266460 215404 266524
rect 244228 266460 244292 266524
rect 252324 266460 252388 266524
rect 260604 266460 260668 266524
rect 267596 266460 267660 266524
rect 412404 266460 412468 266524
rect 419212 266460 419276 266524
rect 86540 266324 86604 266388
rect 87460 266324 87524 266388
rect 88748 266324 88812 266388
rect 90036 266324 90100 266388
rect 93348 266324 93412 266388
rect 107516 266324 107580 266388
rect 108620 266324 108684 266388
rect 114324 266324 114388 266388
rect 215524 266324 215588 266388
rect 245332 266324 245396 266388
rect 246436 266324 246500 266388
rect 247724 266324 247788 266388
rect 248644 266324 248708 266388
rect 251220 266384 251284 266388
rect 251220 266328 251234 266384
rect 251234 266328 251284 266384
rect 251220 266324 251284 266328
rect 253428 266324 253492 266388
rect 254532 266324 254596 266388
rect 256924 266324 256988 266388
rect 259500 266384 259564 266388
rect 259500 266328 259514 266384
rect 259514 266328 259564 266384
rect 259500 266324 259564 266328
rect 262812 266324 262876 266388
rect 263916 266324 263980 266388
rect 266308 266324 266372 266388
rect 268700 266324 268764 266388
rect 269804 266324 269868 266388
rect 271276 266324 271340 266388
rect 274404 266324 274468 266388
rect 396028 266384 396092 266388
rect 396028 266328 396078 266384
rect 396078 266328 396092 266384
rect 396028 266324 396092 266328
rect 399524 266324 399588 266388
rect 400444 266324 400508 266388
rect 404124 266324 404188 266388
rect 405044 266324 405108 266388
rect 406516 266324 406580 266388
rect 407620 266324 407684 266388
rect 410012 266324 410076 266388
rect 411300 266384 411364 266388
rect 411300 266328 411314 266384
rect 411314 266328 411364 266384
rect 411300 266324 411364 266328
rect 413324 266324 413388 266388
rect 418108 266384 418172 266388
rect 418108 266328 418158 266384
rect 418158 266328 418172 266384
rect 418108 266324 418172 266328
rect 420684 266324 420748 266388
rect 421788 266324 421852 266388
rect 427676 266324 427740 266388
rect 436876 266324 436940 266388
rect 272564 266188 272628 266252
rect 240548 266052 240612 266116
rect 241652 265916 241716 265980
rect 239260 265644 239324 265708
rect 426388 265644 426452 265708
rect 238156 265508 238220 265572
rect 431172 265508 431236 265572
rect 57100 262244 57164 262308
rect 53052 253948 53116 254012
rect 377996 250956 378060 251020
rect 178540 249868 178604 249932
rect 179644 249868 179708 249932
rect 190868 249928 190932 249932
rect 190868 249872 190918 249928
rect 190918 249872 190932 249928
rect 190868 249868 190932 249872
rect 338436 249928 338500 249932
rect 338436 249872 338486 249928
rect 338486 249872 338500 249928
rect 338436 249868 338500 249872
rect 339724 249868 339788 249932
rect 350948 249868 351012 249932
rect 498516 249868 498580 249932
rect 499804 249868 499868 249932
rect 510844 249928 510908 249932
rect 510844 249872 510894 249928
rect 510894 249872 510908 249928
rect 510844 249868 510908 249872
rect 44772 249732 44836 249796
rect 44956 249052 45020 249116
rect 200804 174932 200868 174996
rect 96108 164928 96172 164932
rect 96108 164872 96122 164928
rect 96122 164872 96172 164928
rect 96108 164868 96172 164872
rect 115766 164928 115830 164932
rect 115766 164872 115810 164928
rect 115810 164872 115830 164928
rect 115766 164868 115830 164872
rect 413462 164868 413526 164932
rect 138478 164792 138542 164796
rect 138478 164736 138534 164792
rect 138534 164736 138542 164792
rect 138478 164732 138542 164736
rect 140926 164732 140990 164796
rect 143510 164792 143574 164796
rect 143510 164736 143538 164792
rect 143538 164736 143574 164792
rect 143510 164732 143574 164736
rect 163366 164792 163430 164796
rect 163366 164736 163374 164792
rect 163374 164736 163430 164792
rect 163366 164732 163430 164736
rect 261078 164732 261142 164796
rect 425974 164792 426038 164796
rect 425974 164736 425978 164792
rect 425978 164736 426034 164792
rect 426034 164736 426038 164792
rect 425974 164732 426038 164736
rect 450998 164792 451062 164796
rect 450998 164736 451002 164792
rect 451002 164736 451058 164792
rect 451058 164736 451062 164792
rect 450998 164732 451062 164736
rect 85438 164596 85502 164660
rect 103526 164656 103590 164660
rect 103526 164600 103574 164656
rect 103574 164600 103590 164656
rect 103526 164596 103590 164600
rect 105974 164596 106038 164660
rect 114406 164656 114470 164660
rect 114406 164600 114430 164656
rect 114430 164600 114470 164656
rect 114406 164596 114470 164600
rect 118078 164656 118142 164660
rect 118078 164600 118110 164656
rect 118110 164600 118142 164656
rect 118078 164596 118142 164600
rect 153438 164596 153502 164660
rect 165950 164596 166014 164660
rect 288278 164656 288342 164660
rect 288278 164600 288310 164656
rect 288310 164600 288342 164656
rect 288278 164596 288342 164600
rect 305958 164656 306022 164660
rect 305958 164600 305974 164656
rect 305974 164600 306022 164656
rect 305958 164596 306022 164600
rect 318470 164596 318534 164660
rect 423526 164656 423590 164660
rect 423526 164600 423550 164656
rect 423550 164600 423590 164656
rect 423526 164596 423590 164600
rect 429782 164656 429846 164660
rect 429782 164600 429806 164656
rect 429806 164600 429846 164656
rect 429782 164596 429846 164600
rect 436990 164596 437054 164660
rect 470990 164656 471054 164660
rect 470990 164600 471022 164656
rect 471022 164600 471054 164656
rect 470990 164596 471054 164600
rect 480918 164656 480982 164660
rect 480918 164600 480958 164656
rect 480958 164600 480982 164656
rect 480918 164596 480982 164600
rect 265940 164520 266004 164524
rect 265940 164464 265954 164520
rect 265954 164464 266004 164520
rect 265940 164460 266004 164464
rect 205220 164324 205284 164388
rect 290964 164324 291028 164388
rect 98500 164248 98564 164252
rect 98500 164192 98514 164248
rect 98514 164192 98564 164248
rect 98500 164188 98564 164192
rect 101076 164248 101140 164252
rect 101076 164192 101090 164248
rect 101090 164192 101140 164248
rect 101076 164188 101140 164192
rect 108252 164248 108316 164252
rect 108252 164192 108266 164248
rect 108266 164192 108316 164248
rect 108252 164188 108316 164192
rect 123524 164188 123588 164252
rect 145972 164248 146036 164252
rect 145972 164192 145986 164248
rect 145986 164192 146036 164248
rect 145972 164188 146036 164192
rect 148548 164248 148612 164252
rect 148548 164192 148562 164248
rect 148562 164192 148612 164248
rect 148548 164188 148612 164192
rect 150940 164248 151004 164252
rect 150940 164192 150954 164248
rect 150954 164192 151004 164248
rect 150940 164188 151004 164192
rect 203012 164188 203076 164252
rect 298508 164248 298572 164252
rect 298508 164192 298522 164248
rect 298522 164192 298572 164248
rect 298508 164188 298572 164192
rect 300900 164248 300964 164252
rect 300900 164192 300914 164248
rect 300914 164192 300964 164248
rect 300900 164188 300964 164192
rect 303476 164248 303540 164252
rect 303476 164192 303490 164248
rect 303490 164192 303540 164248
rect 303476 164188 303540 164192
rect 313412 164248 313476 164252
rect 313412 164192 313426 164248
rect 313426 164192 313476 164248
rect 313412 164188 313476 164192
rect 418476 164248 418540 164252
rect 418476 164192 418490 164248
rect 418490 164192 418540 164248
rect 418476 164188 418540 164192
rect 421052 164248 421116 164252
rect 421052 164192 421066 164248
rect 421066 164192 421116 164248
rect 421052 164188 421116 164192
rect 428228 164248 428292 164252
rect 428228 164192 428242 164248
rect 428242 164192 428292 164248
rect 428228 164188 428292 164192
rect 430988 164248 431052 164252
rect 430988 164192 431002 164248
rect 431002 164192 431052 164248
rect 430988 164188 431052 164192
rect 473492 164248 473556 164252
rect 473492 164192 473506 164248
rect 473506 164192 473556 164248
rect 473492 164188 473556 164192
rect 475884 164248 475948 164252
rect 475884 164192 475898 164248
rect 475898 164192 475948 164248
rect 475884 164188 475948 164192
rect 478460 164248 478524 164252
rect 478460 164192 478474 164248
rect 478474 164192 478524 164248
rect 478460 164188 478524 164192
rect 483428 164248 483492 164252
rect 483428 164192 483442 164248
rect 483442 164192 483492 164248
rect 483428 164188 483492 164192
rect 198228 164052 198292 164116
rect 308444 164052 308508 164116
rect 486004 164052 486068 164116
rect 111196 163976 111260 163980
rect 111196 163920 111210 163976
rect 111210 163920 111260 163976
rect 111196 163916 111260 163920
rect 202460 163916 202524 163980
rect 295932 163916 295996 163980
rect 196572 163780 196636 163844
rect 270908 163780 270972 163844
rect 285996 163840 286060 163844
rect 285996 163784 286010 163840
rect 286010 163784 286060 163840
rect 285996 163780 286060 163784
rect 113404 163704 113468 163708
rect 113404 163648 113454 163704
rect 113454 163648 113468 163704
rect 113404 163644 113468 163648
rect 218836 163644 218900 163708
rect 95924 163100 95988 163164
rect 99420 163160 99484 163164
rect 99420 163104 99434 163160
rect 99434 163104 99484 163160
rect 99420 163100 99484 163104
rect 128308 163160 128372 163164
rect 128308 163104 128358 163160
rect 128358 163104 128372 163160
rect 128308 163100 128372 163104
rect 235948 163160 236012 163164
rect 235948 163104 235998 163160
rect 235998 163104 236012 163160
rect 235948 163100 236012 163104
rect 261708 163100 261772 163164
rect 76052 162752 76116 162756
rect 76052 162696 76066 162752
rect 76066 162696 76116 162752
rect 76052 162692 76116 162696
rect 78260 162692 78324 162756
rect 79548 162692 79612 162756
rect 80468 162692 80532 162756
rect 81940 162692 82004 162756
rect 83044 162692 83108 162756
rect 84332 162692 84396 162756
rect 86540 162692 86604 162756
rect 87644 162692 87708 162756
rect 88748 162692 88812 162756
rect 90036 162692 90100 162756
rect 90772 162752 90836 162756
rect 90772 162696 90786 162752
rect 90786 162696 90836 162752
rect 90772 162692 90836 162696
rect 91324 162692 91388 162756
rect 93348 162692 93412 162756
rect 94452 162692 94516 162756
rect 97028 162692 97092 162756
rect 98132 162692 98196 162756
rect 100708 162752 100772 162756
rect 100708 162696 100758 162752
rect 100758 162696 100772 162752
rect 100708 162692 100772 162696
rect 102732 162692 102796 162756
rect 103836 162752 103900 162756
rect 103836 162696 103850 162752
rect 103850 162696 103900 162752
rect 103836 162692 103900 162696
rect 105308 162692 105372 162756
rect 106412 162692 106476 162756
rect 108620 162692 108684 162756
rect 109540 162692 109604 162756
rect 111012 162752 111076 162756
rect 111012 162696 111026 162752
rect 111026 162696 111076 162752
rect 111012 162692 111076 162696
rect 113220 162752 113284 162756
rect 113220 162696 113234 162752
rect 113234 162696 113284 162752
rect 113220 162692 113284 162696
rect 116900 162692 116964 162756
rect 118372 162752 118436 162756
rect 118372 162696 118386 162752
rect 118386 162696 118436 162752
rect 118372 162692 118436 162696
rect 119108 162692 119172 162756
rect 120764 162752 120828 162756
rect 120764 162696 120778 162752
rect 120778 162696 120828 162752
rect 120764 162692 120828 162696
rect 125916 162752 125980 162756
rect 125916 162696 125930 162752
rect 125930 162696 125980 162752
rect 125916 162692 125980 162696
rect 130884 162752 130948 162756
rect 130884 162696 130898 162752
rect 130898 162696 130948 162752
rect 130884 162692 130948 162696
rect 133460 162752 133524 162756
rect 133460 162696 133474 162752
rect 133474 162696 133524 162752
rect 133460 162692 133524 162696
rect 136036 162752 136100 162756
rect 136036 162696 136050 162752
rect 136050 162696 136100 162752
rect 136036 162692 136100 162696
rect 155908 162752 155972 162756
rect 155908 162696 155958 162752
rect 155958 162696 155972 162752
rect 155908 162692 155972 162696
rect 183508 162752 183572 162756
rect 183508 162696 183522 162752
rect 183522 162696 183572 162752
rect 183508 162692 183572 162696
rect 237052 162692 237116 162756
rect 238156 162692 238220 162756
rect 240548 162692 240612 162756
rect 241652 162692 241716 162756
rect 242940 162752 243004 162756
rect 242940 162696 242954 162752
rect 242954 162696 243004 162752
rect 242940 162692 243004 162696
rect 244228 162692 244292 162756
rect 246436 162692 246500 162756
rect 247724 162692 247788 162756
rect 248276 162752 248340 162756
rect 248276 162696 248290 162752
rect 248290 162696 248340 162752
rect 248276 162692 248340 162696
rect 248644 162692 248708 162756
rect 250116 162692 250180 162756
rect 250668 162752 250732 162756
rect 250668 162696 250682 162752
rect 250682 162696 250732 162752
rect 250668 162692 250732 162696
rect 251220 162752 251284 162756
rect 251220 162696 251234 162752
rect 251234 162696 251284 162752
rect 251220 162692 251284 162696
rect 253428 162692 253492 162756
rect 253612 162752 253676 162756
rect 253612 162696 253626 162752
rect 253626 162696 253676 162752
rect 253612 162692 253676 162696
rect 254532 162692 254596 162756
rect 255820 162692 255884 162756
rect 256188 162752 256252 162756
rect 256188 162696 256202 162752
rect 256202 162696 256252 162752
rect 256188 162692 256252 162696
rect 256924 162692 256988 162756
rect 258396 162752 258460 162756
rect 258396 162696 258410 162752
rect 258410 162696 258460 162752
rect 258396 162692 258460 162696
rect 259500 162752 259564 162756
rect 265204 163100 265268 163164
rect 272196 163100 272260 163164
rect 276060 163160 276124 163164
rect 276060 163104 276110 163160
rect 276110 163104 276124 163160
rect 276060 163100 276124 163104
rect 398236 163100 398300 163164
rect 263548 162828 263612 162892
rect 268332 162888 268396 162892
rect 268332 162832 268346 162888
rect 268346 162832 268396 162888
rect 268332 162828 268396 162832
rect 259500 162696 259514 162752
rect 259514 162696 259564 162752
rect 259500 162692 259564 162696
rect 262812 162692 262876 162756
rect 263916 162692 263980 162756
rect 266308 162752 266372 162756
rect 266308 162696 266358 162752
rect 266358 162696 266372 162752
rect 266308 162692 266372 162696
rect 267596 162752 267660 162756
rect 267596 162696 267610 162752
rect 267610 162696 267660 162752
rect 267596 162692 267660 162696
rect 268700 162692 268764 162756
rect 269804 162692 269868 162756
rect 271092 162692 271156 162756
rect 273484 162888 273548 162892
rect 273484 162832 273498 162888
rect 273498 162832 273548 162888
rect 273484 162828 273548 162832
rect 274404 162692 274468 162756
rect 275324 162692 275388 162756
rect 276980 162692 277044 162756
rect 279004 162692 279068 162756
rect 280844 162752 280908 162756
rect 280844 162696 280858 162752
rect 280858 162696 280908 162752
rect 280844 162692 280908 162696
rect 283788 162752 283852 162756
rect 283788 162696 283802 162752
rect 283802 162696 283852 162752
rect 283788 162692 283852 162696
rect 293356 162692 293420 162756
rect 320956 162752 321020 162756
rect 320956 162696 320970 162752
rect 320970 162696 321020 162752
rect 320956 162692 321020 162696
rect 343404 162752 343468 162756
rect 343404 162696 343454 162752
rect 343454 162696 343468 162752
rect 343404 162692 343468 162696
rect 396028 162752 396092 162756
rect 396028 162696 396078 162752
rect 396078 162696 396092 162752
rect 396028 162692 396092 162696
rect 401732 163100 401796 163164
rect 416084 163160 416148 163164
rect 416084 163104 416098 163160
rect 416098 163104 416148 163160
rect 416084 163100 416148 163104
rect 455828 163160 455892 163164
rect 455828 163104 455842 163160
rect 455842 163104 455892 163160
rect 455828 163100 455892 163104
rect 399524 162692 399588 162756
rect 400444 162692 400508 162756
rect 403020 162752 403084 162756
rect 403020 162696 403070 162752
rect 403070 162696 403084 162752
rect 403020 162692 403084 162696
rect 405044 162692 405108 162756
rect 406516 162692 406580 162756
rect 407620 162692 407684 162756
rect 408356 162752 408420 162756
rect 408356 162696 408370 162752
rect 408370 162696 408420 162752
rect 408356 162692 408420 162696
rect 408724 162692 408788 162756
rect 410012 162692 410076 162756
rect 410748 162692 410812 162756
rect 411300 162752 411364 162756
rect 411300 162696 411350 162752
rect 411350 162696 411364 162752
rect 411300 162692 411364 162696
rect 413692 162692 413756 162756
rect 414612 162692 414676 162756
rect 415532 162752 415596 162756
rect 415532 162696 415546 162752
rect 415546 162696 415596 162752
rect 415532 162692 415596 162696
rect 417004 162692 417068 162756
rect 419212 162692 419276 162756
rect 420684 162692 420748 162756
rect 421788 162692 421852 162756
rect 422892 162692 422956 162756
rect 423996 162692 424060 162756
rect 425284 162692 425348 162756
rect 426388 162752 426452 162756
rect 426388 162696 426438 162752
rect 426438 162696 426452 162752
rect 426388 162692 426452 162696
rect 428780 162692 428844 162756
rect 431172 162692 431236 162756
rect 431724 162692 431788 162756
rect 434668 162692 434732 162756
rect 435772 162752 435836 162756
rect 435772 162696 435786 162752
rect 435786 162696 435836 162752
rect 435772 162692 435836 162696
rect 435956 162752 436020 162756
rect 435956 162696 435970 162752
rect 435970 162696 436020 162752
rect 435956 162692 436020 162696
rect 438348 162692 438412 162756
rect 438532 162752 438596 162756
rect 438532 162696 438546 162752
rect 438546 162696 438596 162752
rect 438532 162692 438596 162696
rect 439084 162692 439148 162756
rect 440924 162752 440988 162756
rect 440924 162696 440938 162752
rect 440938 162696 440988 162752
rect 440924 162692 440988 162696
rect 443500 162752 443564 162756
rect 443500 162696 443514 162752
rect 443514 162696 443564 162752
rect 443500 162692 443564 162696
rect 445892 162752 445956 162756
rect 445892 162696 445906 162752
rect 445906 162696 445956 162752
rect 445892 162692 445956 162696
rect 448284 162752 448348 162756
rect 448284 162696 448298 162752
rect 448298 162696 448348 162752
rect 448284 162692 448348 162696
rect 453436 162752 453500 162756
rect 453436 162696 453450 162752
rect 453450 162696 453500 162752
rect 453436 162692 453500 162696
rect 458404 162752 458468 162756
rect 458404 162696 458418 162752
rect 458418 162696 458468 162752
rect 458404 162692 458468 162696
rect 503116 162692 503180 162756
rect 158484 162556 158548 162620
rect 183140 162616 183204 162620
rect 183140 162560 183190 162616
rect 183190 162560 183204 162616
rect 183140 162556 183204 162560
rect 207980 162556 208044 162620
rect 323348 162556 323412 162620
rect 343220 162556 343284 162620
rect 468524 162556 468588 162620
rect 503484 162556 503548 162620
rect 47900 162420 47964 162484
rect 91508 162420 91572 162484
rect 107516 162420 107580 162484
rect 115980 162480 116044 162484
rect 115980 162424 116030 162480
rect 116030 162424 116044 162480
rect 115980 162420 116044 162424
rect 203196 162420 203260 162484
rect 311020 162420 311084 162484
rect 462636 162420 462700 162484
rect 47716 162284 47780 162348
rect 160876 162284 160940 162348
rect 213316 162284 213380 162348
rect 315068 162284 315132 162348
rect 460980 162284 461044 162348
rect 77156 162148 77220 162212
rect 88380 162208 88444 162212
rect 88380 162152 88394 162208
rect 88394 162152 88444 162208
rect 88380 162148 88444 162152
rect 93716 162148 93780 162212
rect 112300 162148 112364 162212
rect 215892 162148 215956 162212
rect 278452 162148 278516 162212
rect 397132 162148 397196 162212
rect 404124 162148 404188 162212
rect 412404 162148 412468 162212
rect 418108 162148 418172 162212
rect 427676 162148 427740 162212
rect 433380 162148 433444 162212
rect 101812 162012 101876 162076
rect 245332 162012 245396 162076
rect 252324 162012 252388 162076
rect 260604 162012 260668 162076
rect 273300 162012 273364 162076
rect 433564 162072 433628 162076
rect 433564 162016 433578 162072
rect 433578 162016 433628 162072
rect 433564 162012 433628 162016
rect 206324 161740 206388 161804
rect 326660 161740 326724 161804
rect 465948 161740 466012 161804
rect 238708 161528 238772 161532
rect 238708 161472 238758 161528
rect 238758 161472 238772 161528
rect 238708 161468 238772 161472
rect 258396 161468 258460 161532
rect 277348 161468 277412 161532
rect 217548 161060 217612 161124
rect 57836 160108 57900 160172
rect 360884 149092 360948 149156
rect 379468 148412 379532 148476
rect 217364 148276 217428 148340
rect 377628 148276 377692 148340
rect 57284 147460 57348 147524
rect 217180 146372 217244 146436
rect 377996 146236 378060 146300
rect 57652 145692 57716 145756
rect 190868 145420 190932 145484
rect 377812 145556 377876 145620
rect 510844 145420 510908 145484
rect 178540 144876 178604 144940
rect 179644 144936 179708 144940
rect 179644 144880 179694 144936
rect 179694 144880 179708 144936
rect 179644 144876 179708 144880
rect 338436 144936 338500 144940
rect 338436 144880 338486 144936
rect 338486 144880 338500 144936
rect 338436 144876 338500 144880
rect 339724 144876 339788 144940
rect 350948 144876 351012 144940
rect 498516 144876 498580 144940
rect 499804 144876 499868 144940
rect 57100 144740 57164 144804
rect 57652 144740 57716 144804
rect 57468 140796 57532 140860
rect 46796 68988 46860 69052
rect 205036 68036 205100 68100
rect 367876 68036 367940 68100
rect 218652 60616 218716 60620
rect 218652 60560 218702 60616
rect 218702 60560 218716 60616
rect 218652 60556 218716 60560
rect 219204 60616 219268 60620
rect 219204 60560 219254 60616
rect 219254 60560 219268 60616
rect 219204 60556 219268 60560
rect 77142 59800 77206 59804
rect 77142 59744 77170 59800
rect 77170 59744 77206 59800
rect 77142 59740 77206 59744
rect 83126 59800 83190 59804
rect 83126 59744 83150 59800
rect 83150 59744 83190 59800
rect 83126 59740 83190 59744
rect 99446 59800 99510 59804
rect 99446 59744 99470 59800
rect 99470 59744 99510 59800
rect 99446 59740 99510 59744
rect 113590 59800 113654 59804
rect 113590 59744 113602 59800
rect 113602 59744 113654 59800
rect 113590 59740 113654 59744
rect 237142 59800 237206 59804
rect 237142 59744 237158 59800
rect 237158 59744 237206 59800
rect 237142 59740 237206 59744
rect 255910 59800 255974 59804
rect 255910 59744 255926 59800
rect 255926 59744 255974 59800
rect 255910 59740 255974 59744
rect 256998 59800 257062 59804
rect 256998 59744 257030 59800
rect 257030 59744 257062 59800
rect 256998 59740 257062 59744
rect 261758 59800 261822 59804
rect 261758 59744 261814 59800
rect 261814 59744 261822 59800
rect 261758 59740 261822 59744
rect 263934 59740 263998 59804
rect 396054 59800 396118 59804
rect 396054 59744 396078 59800
rect 396078 59744 396118 59800
rect 396054 59740 396118 59744
rect 397142 59800 397206 59804
rect 397142 59744 397146 59800
rect 397146 59744 397206 59800
rect 397142 59740 397206 59744
rect 416998 59800 417062 59804
rect 416998 59744 417018 59800
rect 417018 59744 417062 59800
rect 416998 59740 417062 59744
rect 418494 59740 418558 59804
rect 423934 59800 423998 59804
rect 423934 59744 423954 59800
rect 423954 59744 423998 59800
rect 423934 59740 423998 59744
rect 94550 59664 94614 59668
rect 94550 59608 94558 59664
rect 94558 59608 94614 59664
rect 94550 59604 94614 59608
rect 101078 59604 101142 59668
rect 102846 59604 102910 59668
rect 103934 59664 103998 59668
rect 103934 59608 103942 59664
rect 103942 59608 103998 59664
rect 103934 59604 103998 59608
rect 260670 59664 260734 59668
rect 260670 59608 260710 59664
rect 260710 59608 260734 59664
rect 260670 59604 260734 59608
rect 305958 59664 306022 59668
rect 305958 59608 305974 59664
rect 305974 59608 306022 59664
rect 305958 59604 306022 59608
rect 318470 59664 318534 59668
rect 318470 59608 318486 59664
rect 318486 59608 318534 59664
rect 318470 59604 318534 59608
rect 403126 59604 403190 59668
rect 404214 59664 404278 59668
rect 404214 59608 404230 59664
rect 404230 59608 404278 59664
rect 404214 59604 404278 59608
rect 413462 59604 413526 59668
rect 419446 59664 419510 59668
rect 419446 59608 419502 59664
rect 419502 59608 419510 59664
rect 419446 59604 419510 59608
rect 421758 59664 421822 59668
rect 421758 59608 421802 59664
rect 421802 59608 421822 59664
rect 421758 59604 421822 59608
rect 423526 59664 423590 59668
rect 423526 59608 423550 59664
rect 423550 59608 423590 59664
rect 423526 59604 423590 59608
rect 503222 59664 503286 59668
rect 503222 59608 503258 59664
rect 503258 59608 503286 59664
rect 503222 59604 503286 59608
rect 57100 59468 57164 59532
rect 100708 59468 100772 59532
rect 262812 59528 262876 59532
rect 262812 59472 262826 59528
rect 262826 59472 262876 59528
rect 262812 59468 262876 59472
rect 418108 59528 418172 59532
rect 418108 59472 418158 59528
rect 418158 59472 418172 59528
rect 418108 59468 418172 59472
rect 420684 59528 420748 59532
rect 420684 59472 420698 59528
rect 420698 59472 420748 59528
rect 420684 59468 420748 59472
rect 46612 59332 46676 59396
rect 95924 59392 95988 59396
rect 95924 59336 95938 59392
rect 95938 59336 95988 59392
rect 95924 59332 95988 59336
rect 97028 59392 97092 59396
rect 97028 59336 97042 59392
rect 97042 59336 97092 59392
rect 97028 59332 97092 59336
rect 101812 59392 101876 59396
rect 101812 59336 101826 59392
rect 101826 59336 101876 59392
rect 101812 59332 101876 59336
rect 111196 59392 111260 59396
rect 111196 59336 111210 59392
rect 111210 59336 111260 59392
rect 111196 59332 111260 59336
rect 115980 59392 116044 59396
rect 115980 59336 115994 59392
rect 115994 59336 116044 59392
rect 115980 59332 116044 59336
rect 198044 59332 198108 59396
rect 263548 59332 263612 59396
rect 377812 59332 377876 59396
rect 422892 59332 422956 59396
rect 425284 59392 425348 59396
rect 425284 59336 425298 59392
rect 425298 59336 425348 59392
rect 425284 59332 425348 59336
rect 426020 59392 426084 59396
rect 426020 59336 426034 59392
rect 426034 59336 426084 59392
rect 426020 59332 426084 59336
rect 428228 59392 428292 59396
rect 428228 59336 428242 59392
rect 428242 59336 428292 59392
rect 428228 59332 428292 59336
rect 465948 59392 466012 59396
rect 465948 59336 465962 59392
rect 465962 59336 466012 59392
rect 465948 59332 466012 59336
rect 52316 59196 52380 59260
rect 143580 59196 143644 59260
rect 148548 59256 148612 59260
rect 148548 59200 148562 59256
rect 148562 59200 148612 59256
rect 148548 59196 148612 59200
rect 150940 59256 151004 59260
rect 150940 59200 150954 59256
rect 150954 59200 151004 59256
rect 150940 59196 151004 59200
rect 201356 59196 201420 59260
rect 279188 59256 279252 59260
rect 279188 59200 279238 59256
rect 279238 59200 279252 59256
rect 54708 59060 54772 59124
rect 140820 59060 140884 59124
rect 198596 59060 198660 59124
rect 273484 59060 273548 59124
rect 279188 59196 279252 59200
rect 290964 59256 291028 59260
rect 290964 59200 290978 59256
rect 290978 59200 291028 59256
rect 290964 59196 291028 59200
rect 298508 59256 298572 59260
rect 298508 59200 298522 59256
rect 298522 59200 298572 59256
rect 298508 59196 298572 59200
rect 313412 59256 313476 59260
rect 313412 59200 313426 59256
rect 313426 59200 313476 59256
rect 313412 59196 313476 59200
rect 325924 59256 325988 59260
rect 325924 59200 325938 59256
rect 325938 59200 325988 59256
rect 325924 59196 325988 59200
rect 360700 59196 360764 59260
rect 483428 59196 483492 59260
rect 486004 59256 486068 59260
rect 486004 59200 486018 59256
rect 486018 59200 486068 59256
rect 486004 59196 486068 59200
rect 285996 59060 286060 59124
rect 357940 59060 358004 59124
rect 475884 59060 475948 59124
rect 53420 58924 53484 58988
rect 138428 58924 138492 58988
rect 206876 58924 206940 58988
rect 276060 58924 276124 58988
rect 371740 58924 371804 58988
rect 480852 58924 480916 58988
rect 51948 58788 52012 58852
rect 135852 58788 135916 58852
rect 213684 58788 213748 58852
rect 278452 58788 278516 58852
rect 375972 58788 376036 58852
rect 470916 58788 470980 58852
rect 59308 58652 59372 58716
rect 120948 58652 121012 58716
rect 197860 58652 197924 58716
rect 253612 58652 253676 58716
rect 259500 58712 259564 58716
rect 259500 58656 259514 58712
rect 259514 58656 259564 58712
rect 259500 58652 259564 58656
rect 370452 58652 370516 58716
rect 458404 58652 458468 58716
rect 48084 58516 48148 58580
rect 108252 58516 108316 58580
rect 202092 58516 202156 58580
rect 250668 58516 250732 58580
rect 374684 58516 374748 58580
rect 463556 58516 463620 58580
rect 52132 58380 52196 58444
rect 111012 58380 111076 58444
rect 217548 58380 217612 58444
rect 257844 58380 257908 58444
rect 367692 58380 367756 58444
rect 453436 58380 453500 58444
rect 85436 58108 85500 58172
rect 92244 58108 92308 58172
rect 153332 58108 153396 58172
rect 235948 58108 236012 58172
rect 265204 58108 265268 58172
rect 272196 58108 272260 58172
rect 275692 58108 275756 58172
rect 300900 58108 300964 58172
rect 315804 58108 315868 58172
rect 398236 58108 398300 58172
rect 401732 58108 401796 58172
rect 405412 58108 405476 58172
rect 416084 58108 416148 58172
rect 83964 57972 84028 58036
rect 76052 57896 76116 57900
rect 76052 57840 76066 57896
rect 76066 57840 76116 57896
rect 76052 57836 76116 57840
rect 78260 57896 78324 57900
rect 78260 57840 78274 57896
rect 78274 57840 78324 57896
rect 78260 57836 78324 57840
rect 79548 57896 79612 57900
rect 79548 57840 79562 57896
rect 79562 57840 79612 57896
rect 79548 57836 79612 57840
rect 80468 57836 80532 57900
rect 81940 57836 82004 57900
rect 86540 57896 86604 57900
rect 86540 57840 86554 57896
rect 86554 57840 86604 57896
rect 86540 57836 86604 57840
rect 87644 57836 87708 57900
rect 88380 57896 88444 57900
rect 88380 57840 88394 57896
rect 88394 57840 88444 57896
rect 88380 57836 88444 57840
rect 88748 57896 88812 57900
rect 88748 57840 88762 57896
rect 88762 57840 88812 57896
rect 88748 57836 88812 57840
rect 90036 57836 90100 57900
rect 90772 57896 90836 57900
rect 90772 57840 90786 57896
rect 90786 57840 90836 57896
rect 90772 57836 90836 57840
rect 91324 57836 91388 57900
rect 93348 57836 93412 57900
rect 93716 57896 93780 57900
rect 93716 57840 93730 57896
rect 93730 57840 93780 57896
rect 93716 57836 93780 57840
rect 98132 57896 98196 57900
rect 98132 57840 98146 57896
rect 98146 57840 98196 57896
rect 98132 57836 98196 57840
rect 106412 57896 106476 57900
rect 106412 57840 106426 57896
rect 106426 57840 106476 57896
rect 106412 57836 106476 57840
rect 107516 57836 107580 57900
rect 108620 57836 108684 57900
rect 112116 57896 112180 57900
rect 112116 57840 112130 57896
rect 112130 57840 112180 57896
rect 112116 57836 112180 57840
rect 113220 57896 113284 57900
rect 113220 57840 113234 57896
rect 113234 57840 113284 57896
rect 113220 57836 113284 57840
rect 123524 57896 123588 57900
rect 123524 57840 123538 57896
rect 123538 57840 123588 57896
rect 123524 57836 123588 57840
rect 130884 57896 130948 57900
rect 130884 57840 130898 57896
rect 130898 57840 130948 57896
rect 130884 57836 130948 57840
rect 133460 57836 133524 57900
rect 145604 57896 145668 57900
rect 145604 57840 145618 57896
rect 145618 57840 145668 57896
rect 145604 57836 145668 57840
rect 158484 57836 158548 57900
rect 183140 57836 183204 57900
rect 238156 57836 238220 57900
rect 239260 57896 239324 57900
rect 239260 57840 239274 57896
rect 239274 57840 239324 57896
rect 239260 57836 239324 57840
rect 240548 57836 240612 57900
rect 241652 57896 241716 57900
rect 241652 57840 241666 57896
rect 241666 57840 241716 57896
rect 241652 57836 241716 57840
rect 242940 57896 243004 57900
rect 242940 57840 242954 57896
rect 242954 57840 243004 57896
rect 242940 57836 243004 57840
rect 244228 57836 244292 57900
rect 245332 57896 245396 57900
rect 245332 57840 245346 57896
rect 245346 57840 245396 57896
rect 245332 57836 245396 57840
rect 246436 57836 246500 57900
rect 247724 57836 247788 57900
rect 248644 57896 248708 57900
rect 248644 57840 248658 57896
rect 248658 57840 248708 57896
rect 248644 57836 248708 57840
rect 250116 57836 250180 57900
rect 251220 57896 251284 57900
rect 251220 57840 251234 57896
rect 251234 57840 251284 57896
rect 251220 57836 251284 57840
rect 252324 57836 252388 57900
rect 253428 57896 253492 57900
rect 253428 57840 253442 57896
rect 253442 57840 253492 57896
rect 253428 57836 253492 57840
rect 254532 57836 254596 57900
rect 265940 57896 266004 57900
rect 265940 57840 265954 57896
rect 265954 57840 266004 57896
rect 265940 57836 266004 57840
rect 266308 57896 266372 57900
rect 266308 57840 266358 57896
rect 266358 57840 266372 57896
rect 266308 57836 266372 57840
rect 268700 57836 268764 57900
rect 271276 57896 271340 57900
rect 271276 57840 271290 57896
rect 271290 57840 271340 57896
rect 271276 57836 271340 57840
rect 273300 57896 273364 57900
rect 273300 57840 273314 57896
rect 273314 57840 273364 57896
rect 273300 57836 273364 57840
rect 288204 57836 288268 57900
rect 293356 57896 293420 57900
rect 293356 57840 293370 57896
rect 293370 57840 293420 57896
rect 293356 57836 293420 57840
rect 295932 57896 295996 57900
rect 295932 57840 295946 57896
rect 295946 57840 295996 57896
rect 295932 57836 295996 57840
rect 303476 57896 303540 57900
rect 303476 57840 303490 57896
rect 303490 57840 303540 57896
rect 303476 57836 303540 57840
rect 308628 57836 308692 57900
rect 311020 57896 311084 57900
rect 311020 57840 311034 57896
rect 311034 57840 311084 57896
rect 311020 57836 311084 57840
rect 320956 57896 321020 57900
rect 320956 57840 320970 57896
rect 320970 57840 321020 57896
rect 320956 57836 321020 57840
rect 323348 57896 323412 57900
rect 323348 57840 323362 57896
rect 323362 57840 323412 57896
rect 323348 57836 323412 57840
rect 343220 57896 343284 57900
rect 343220 57840 343234 57896
rect 343234 57840 343284 57896
rect 343220 57836 343284 57840
rect 343404 57896 343468 57900
rect 343404 57840 343454 57896
rect 343454 57840 343468 57896
rect 343404 57836 343468 57840
rect 399524 57896 399588 57900
rect 399524 57840 399538 57896
rect 399538 57840 399588 57896
rect 399524 57836 399588 57840
rect 400444 57836 400508 57900
rect 406516 57836 406580 57900
rect 407620 57836 407684 57900
rect 408356 57896 408420 57900
rect 408356 57840 408370 57896
rect 408370 57840 408420 57896
rect 408356 57836 408420 57840
rect 408724 57896 408788 57900
rect 408724 57840 408738 57896
rect 408738 57840 408788 57896
rect 408724 57836 408788 57840
rect 410012 57836 410076 57900
rect 412404 57836 412468 57900
rect 414612 57896 414676 57900
rect 414612 57840 414626 57896
rect 414626 57840 414676 57896
rect 414612 57836 414676 57840
rect 415532 57896 415596 57900
rect 415532 57840 415546 57896
rect 415546 57840 415596 57896
rect 415532 57836 415596 57840
rect 426388 57896 426452 57900
rect 426388 57840 426438 57896
rect 426438 57840 426452 57896
rect 426388 57836 426452 57840
rect 427676 57896 427740 57900
rect 427676 57840 427690 57896
rect 427690 57840 427740 57896
rect 427676 57836 427740 57840
rect 428596 57836 428660 57900
rect 429700 57836 429764 57900
rect 431172 57836 431236 57900
rect 432276 57836 432340 57900
rect 434668 57836 434732 57900
rect 435956 57896 436020 57900
rect 435956 57840 435970 57896
rect 435970 57840 436020 57896
rect 435956 57836 436020 57840
rect 436876 57836 436940 57900
rect 438348 57896 438412 57900
rect 438348 57840 438362 57896
rect 438362 57840 438412 57896
rect 438348 57836 438412 57840
rect 438532 57896 438596 57900
rect 438532 57840 438546 57896
rect 438546 57840 438596 57896
rect 438532 57836 438596 57840
rect 439084 57836 439148 57900
rect 440924 57896 440988 57900
rect 440924 57840 440938 57896
rect 440938 57840 440988 57896
rect 440924 57836 440988 57840
rect 443500 57896 443564 57900
rect 443500 57840 443514 57896
rect 443514 57840 443564 57896
rect 443500 57836 443564 57840
rect 445892 57896 445956 57900
rect 445892 57840 445906 57896
rect 445906 57840 445956 57896
rect 445892 57836 445956 57840
rect 451044 57896 451108 57900
rect 451044 57840 451058 57896
rect 451058 57840 451108 57896
rect 451044 57836 451108 57840
rect 478460 57896 478524 57900
rect 478460 57840 478474 57896
rect 478474 57840 478524 57896
rect 478460 57836 478524 57840
rect 503300 57896 503364 57900
rect 503300 57840 503350 57896
rect 503350 57840 503364 57896
rect 503300 57836 503364 57840
rect 60228 57700 60292 57764
rect 125916 57700 125980 57764
rect 183508 57760 183572 57764
rect 183508 57704 183522 57760
rect 183522 57704 183572 57760
rect 183508 57700 183572 57704
rect 214420 57700 214484 57764
rect 280844 57700 280908 57764
rect 378732 57700 378796 57764
rect 473308 57700 473372 57764
rect 55076 57564 55140 57628
rect 58940 57428 59004 57492
rect 109540 57564 109604 57628
rect 114324 57564 114388 57628
rect 115796 57564 115860 57628
rect 116900 57564 116964 57628
rect 118004 57564 118068 57628
rect 119108 57564 119172 57628
rect 155908 57624 155972 57628
rect 155908 57568 155958 57624
rect 155958 57568 155972 57624
rect 155908 57564 155972 57568
rect 160876 57564 160940 57628
rect 165844 57564 165908 57628
rect 209084 57564 209148 57628
rect 118372 57428 118436 57492
rect 202276 57428 202340 57492
rect 258396 57428 258460 57492
rect 267596 57564 267660 57628
rect 269804 57564 269868 57628
rect 274404 57564 274468 57628
rect 276980 57564 277044 57628
rect 371924 57564 371988 57628
rect 460980 57564 461044 57628
rect 270908 57428 270972 57492
rect 378916 57428 378980 57492
rect 456380 57428 456444 57492
rect 58756 57292 58820 57356
rect 103836 57292 103900 57356
rect 204852 57292 204916 57356
rect 256004 57292 256068 57356
rect 376156 57292 376220 57356
rect 448284 57292 448348 57356
rect 59124 57156 59188 57220
rect 98500 57156 98564 57220
rect 213132 57156 213196 57220
rect 260972 57156 261036 57220
rect 379284 57156 379348 57220
rect 421052 57156 421116 57220
rect 430988 57216 431052 57220
rect 430988 57160 431002 57216
rect 431002 57160 431052 57216
rect 430988 57156 431052 57160
rect 433380 57216 433444 57220
rect 433380 57160 433394 57216
rect 433394 57160 433444 57216
rect 433380 57156 433444 57160
rect 433564 57216 433628 57220
rect 433564 57160 433578 57216
rect 433578 57160 433628 57216
rect 433564 57156 433628 57160
rect 435772 57216 435836 57220
rect 435772 57160 435786 57216
rect 435786 57160 435836 57216
rect 435772 57156 435836 57160
rect 58572 57020 58636 57084
rect 96292 57020 96356 57084
rect 105860 57020 105924 57084
rect 211660 57020 211724 57084
rect 248276 57020 248340 57084
rect 379100 57020 379164 57084
rect 413508 57020 413572 57084
rect 411300 56944 411364 56948
rect 411300 56888 411314 56944
rect 411314 56888 411364 56944
rect 411300 56884 411364 56888
rect 54892 56612 54956 56676
rect 128676 56612 128740 56676
rect 163268 56612 163332 56676
rect 214604 56612 214668 56676
rect 283788 56612 283852 56676
rect 363644 56612 363708 56676
rect 468524 56612 468588 56676
rect 53604 56476 53668 56540
rect 219940 56476 220004 56540
rect 410748 56476 410812 56540
rect 55628 56340 55692 56404
rect 200620 56340 200684 56404
rect 268332 56340 268396 56404
rect 57652 56204 57716 56268
rect 105308 56204 105372 56268
rect 217364 56204 217428 56268
rect 277164 56204 277228 56268
rect 50476 55116 50540 55180
rect 217180 55116 217244 55180
rect 377628 55116 377692 55180
rect 50844 54980 50908 55044
rect 379468 54980 379532 55044
rect 50660 54844 50724 54908
rect 57468 54708 57532 54772
rect 57836 54572 57900 54636
rect 208900 3980 208964 4044
rect 206140 3844 206204 3908
rect 365116 3708 365180 3772
rect 363460 3572 363524 3636
rect 374500 3436 374564 3500
rect 364932 3300 364996 3364
rect 210372 3164 210436 3228
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 44771 469980 44837 469981
rect 44771 469916 44772 469980
rect 44836 469916 44837 469980
rect 44771 469915 44837 469916
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 44774 249797 44834 469915
rect 44955 469844 45021 469845
rect 44955 469780 44956 469844
rect 45020 469780 45021 469844
rect 44955 469779 45021 469780
rect 44771 249796 44837 249797
rect 44771 249732 44772 249796
rect 44836 249732 44837 249796
rect 44771 249731 44837 249732
rect 44958 249117 45018 469779
rect 45234 442894 45854 478338
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 53051 630868 53117 630869
rect 53051 630804 53052 630868
rect 53116 630804 53117 630868
rect 53051 630803 53117 630804
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 46795 478140 46861 478141
rect 46795 478076 46796 478140
rect 46860 478076 46861 478140
rect 46795 478075 46861 478076
rect 46611 460732 46677 460733
rect 46611 460668 46612 460732
rect 46676 460668 46677 460732
rect 46611 460667 46677 460668
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 44955 249116 45021 249117
rect 44955 249052 44956 249116
rect 45020 249052 45021 249116
rect 44955 249051 45021 249052
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 46614 59397 46674 460667
rect 46798 69053 46858 478075
rect 47899 465900 47965 465901
rect 47899 465836 47900 465900
rect 47964 465836 47965 465900
rect 47899 465835 47965 465836
rect 47715 462908 47781 462909
rect 47715 462844 47716 462908
rect 47780 462844 47781 462908
rect 47715 462843 47781 462844
rect 47718 162349 47778 462843
rect 47902 162485 47962 465835
rect 48083 460868 48149 460869
rect 48083 460804 48084 460868
rect 48148 460804 48149 460868
rect 48083 460803 48149 460804
rect 47899 162484 47965 162485
rect 47899 162420 47900 162484
rect 47964 162420 47965 162484
rect 47899 162419 47965 162420
rect 47715 162348 47781 162349
rect 47715 162284 47716 162348
rect 47780 162284 47781 162348
rect 47715 162283 47781 162284
rect 46795 69052 46861 69053
rect 46795 68988 46796 69052
rect 46860 68988 46861 69052
rect 46795 68987 46861 68988
rect 46611 59396 46677 59397
rect 46611 59332 46612 59396
rect 46676 59332 46677 59396
rect 46611 59331 46677 59332
rect 48086 58581 48146 460803
rect 48954 446614 49574 482058
rect 52315 478276 52381 478277
rect 52315 478212 52316 478276
rect 52380 478212 52381 478276
rect 52315 478211 52381 478212
rect 50843 477596 50909 477597
rect 50843 477532 50844 477596
rect 50908 477532 50909 477596
rect 50843 477531 50909 477532
rect 50659 460188 50725 460189
rect 50659 460124 50660 460188
rect 50724 460124 50725 460188
rect 50659 460123 50725 460124
rect 50475 459644 50541 459645
rect 50475 459580 50476 459644
rect 50540 459580 50541 459644
rect 50475 459579 50541 459580
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48083 58580 48149 58581
rect 48083 58516 48084 58580
rect 48148 58516 48149 58580
rect 48083 58515 48149 58516
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 50614 49574 86058
rect 50478 55181 50538 459579
rect 50475 55180 50541 55181
rect 50475 55116 50476 55180
rect 50540 55116 50541 55180
rect 50475 55115 50541 55116
rect 50662 54909 50722 460123
rect 50846 55045 50906 477531
rect 52131 463452 52197 463453
rect 52131 463388 52132 463452
rect 52196 463388 52197 463452
rect 52131 463387 52197 463388
rect 51947 460460 52013 460461
rect 51947 460396 51948 460460
rect 52012 460396 52013 460460
rect 51947 460395 52013 460396
rect 51763 460324 51829 460325
rect 51763 460260 51764 460324
rect 51828 460260 51829 460324
rect 51763 460259 51829 460260
rect 51766 375325 51826 460259
rect 51763 375324 51829 375325
rect 51763 375260 51764 375324
rect 51828 375260 51829 375324
rect 51763 375259 51829 375260
rect 51950 58853 52010 460395
rect 51947 58852 52013 58853
rect 51947 58788 51948 58852
rect 52012 58788 52013 58852
rect 51947 58787 52013 58788
rect 52134 58445 52194 463387
rect 52318 59261 52378 478211
rect 53054 254013 53114 630803
rect 54339 630732 54405 630733
rect 54339 630668 54340 630732
rect 54404 630668 54405 630732
rect 54339 630667 54405 630668
rect 53235 477596 53301 477597
rect 53235 477532 53236 477596
rect 53300 477532 53301 477596
rect 53235 477531 53301 477532
rect 53238 375325 53298 477531
rect 53419 460052 53485 460053
rect 53419 459988 53420 460052
rect 53484 459988 53485 460052
rect 53419 459987 53485 459988
rect 53235 375324 53301 375325
rect 53235 375260 53236 375324
rect 53300 375260 53301 375324
rect 53235 375259 53301 375260
rect 53051 254012 53117 254013
rect 53051 253948 53052 254012
rect 53116 253948 53117 254012
rect 53051 253947 53117 253948
rect 52315 59260 52381 59261
rect 52315 59196 52316 59260
rect 52380 59196 52381 59260
rect 52315 59195 52381 59196
rect 53422 58989 53482 459987
rect 53603 459644 53669 459645
rect 53603 459580 53604 459644
rect 53668 459580 53669 459644
rect 53603 459579 53669 459580
rect 53419 58988 53485 58989
rect 53419 58924 53420 58988
rect 53484 58924 53485 58988
rect 53419 58923 53485 58924
rect 52131 58444 52197 58445
rect 52131 58380 52132 58444
rect 52196 58380 52197 58444
rect 52131 58379 52197 58380
rect 53606 56541 53666 459579
rect 54342 305013 54402 630667
rect 55794 597454 56414 632898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 625099 60134 636618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 625099 63854 640338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 625099 67574 644058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 625099 74414 650898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 625099 78134 654618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 625099 81854 658338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 625099 85574 626058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 625099 92414 632898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 625099 96134 636618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 625099 99854 640338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 625099 103574 644058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 625099 110414 650898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 625099 114134 654618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 625099 117854 658338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 625099 121574 626058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 64208 615454 64528 615486
rect 64208 615218 64250 615454
rect 64486 615218 64528 615454
rect 64208 615134 64528 615218
rect 64208 614898 64250 615134
rect 64486 614898 64528 615134
rect 64208 614866 64528 614898
rect 94928 615454 95248 615486
rect 94928 615218 94970 615454
rect 95206 615218 95248 615454
rect 94928 615134 95248 615218
rect 94928 614898 94970 615134
rect 95206 614898 95248 615134
rect 94928 614866 95248 614898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 79568 597454 79888 597486
rect 79568 597218 79610 597454
rect 79846 597218 79888 597454
rect 79568 597134 79888 597218
rect 79568 596898 79610 597134
rect 79846 596898 79888 597134
rect 79568 596866 79888 596898
rect 110288 597454 110608 597486
rect 110288 597218 110330 597454
rect 110566 597218 110608 597454
rect 110288 597134 110608 597218
rect 110288 596898 110330 597134
rect 110566 596898 110608 597134
rect 110288 596866 110608 596898
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 64208 579454 64528 579486
rect 64208 579218 64250 579454
rect 64486 579218 64528 579454
rect 64208 579134 64528 579218
rect 64208 578898 64250 579134
rect 64486 578898 64528 579134
rect 64208 578866 64528 578898
rect 94928 579454 95248 579486
rect 94928 579218 94970 579454
rect 95206 579218 95248 579454
rect 94928 579134 95248 579218
rect 94928 578898 94970 579134
rect 95206 578898 95248 579134
rect 94928 578866 95248 578898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 59514 548114 60134 558000
rect 59514 547878 59546 548114
rect 59782 547878 59866 548114
rect 60102 547878 60134 548114
rect 59514 547794 60134 547878
rect 59514 547558 59546 547794
rect 59782 547558 59866 547794
rect 60102 547558 60134 547794
rect 59514 542000 60134 547558
rect 63234 549954 63854 558000
rect 63234 549718 63266 549954
rect 63502 549718 63586 549954
rect 63822 549718 63854 549954
rect 63234 549634 63854 549718
rect 63234 549398 63266 549634
rect 63502 549398 63586 549634
rect 63822 549398 63854 549634
rect 63234 542000 63854 549398
rect 66954 553674 67574 558000
rect 66954 553438 66986 553674
rect 67222 553438 67306 553674
rect 67542 553438 67574 553674
rect 66954 553354 67574 553438
rect 66954 553118 66986 553354
rect 67222 553118 67306 553354
rect 67542 553118 67574 553354
rect 66954 542000 67574 553118
rect 73794 543454 74414 558000
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 542000 74414 542898
rect 77514 547174 78134 558000
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 542000 78134 546618
rect 81234 550894 81854 558000
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 542000 81854 550338
rect 84954 554614 85574 558000
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 542000 85574 554058
rect 91794 544394 92414 558000
rect 91794 544158 91826 544394
rect 92062 544158 92146 544394
rect 92382 544158 92414 544394
rect 91794 544074 92414 544158
rect 91794 543838 91826 544074
rect 92062 543838 92146 544074
rect 92382 543838 92414 544074
rect 91794 542000 92414 543838
rect 95514 548114 96134 558000
rect 95514 547878 95546 548114
rect 95782 547878 95866 548114
rect 96102 547878 96134 548114
rect 95514 547794 96134 547878
rect 95514 547558 95546 547794
rect 95782 547558 95866 547794
rect 96102 547558 96134 547794
rect 95514 542000 96134 547558
rect 99234 549954 99854 558000
rect 99234 549718 99266 549954
rect 99502 549718 99586 549954
rect 99822 549718 99854 549954
rect 99234 549634 99854 549718
rect 99234 549398 99266 549634
rect 99502 549398 99586 549634
rect 99822 549398 99854 549634
rect 99234 542000 99854 549398
rect 102954 553674 103574 558000
rect 102954 553438 102986 553674
rect 103222 553438 103306 553674
rect 103542 553438 103574 553674
rect 102954 553354 103574 553438
rect 102954 553118 102986 553354
rect 103222 553118 103306 553354
rect 103542 553118 103574 553354
rect 102954 542000 103574 553118
rect 109794 543454 110414 558000
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 542000 110414 542898
rect 113514 547174 114134 558000
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 542000 114134 546618
rect 117234 550894 117854 558000
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 542000 117854 550338
rect 120954 554614 121574 558000
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 542000 121574 554058
rect 127794 544394 128414 560898
rect 127794 544158 127826 544394
rect 128062 544158 128146 544394
rect 128382 544158 128414 544394
rect 127794 544074 128414 544158
rect 127794 543838 127826 544074
rect 128062 543838 128146 544074
rect 128382 543838 128414 544074
rect 127794 542000 128414 543838
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 548114 132134 564618
rect 131514 547878 131546 548114
rect 131782 547878 131866 548114
rect 132102 547878 132134 548114
rect 131514 547794 132134 547878
rect 131514 547558 131546 547794
rect 131782 547558 131866 547794
rect 132102 547558 132134 547794
rect 131514 542000 132134 547558
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 625099 139574 644058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 625099 146414 650898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 625099 150134 654618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 625099 153854 658338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 625099 157574 626058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 625099 164414 632898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 625099 168134 636618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 625099 171854 640338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 625099 175574 644058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 625099 182414 650898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 625099 186134 654618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 625099 189854 658338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 625099 193574 626058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 625099 200414 632898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 144208 615454 144528 615486
rect 144208 615218 144250 615454
rect 144486 615218 144528 615454
rect 144208 615134 144528 615218
rect 144208 614898 144250 615134
rect 144486 614898 144528 615134
rect 144208 614866 144528 614898
rect 174928 615454 175248 615486
rect 174928 615218 174970 615454
rect 175206 615218 175248 615454
rect 174928 615134 175248 615218
rect 174928 614898 174970 615134
rect 175206 614898 175248 615134
rect 174928 614866 175248 614898
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 159568 597454 159888 597486
rect 159568 597218 159610 597454
rect 159846 597218 159888 597454
rect 159568 597134 159888 597218
rect 159568 596898 159610 597134
rect 159846 596898 159888 597134
rect 159568 596866 159888 596898
rect 190288 597454 190608 597486
rect 190288 597218 190330 597454
rect 190566 597218 190608 597454
rect 190288 597134 190608 597218
rect 190288 596898 190330 597134
rect 190566 596898 190608 597134
rect 190288 596866 190608 596898
rect 144208 579454 144528 579486
rect 144208 579218 144250 579454
rect 144486 579218 144528 579454
rect 144208 579134 144528 579218
rect 144208 578898 144250 579134
rect 144486 578898 144528 579134
rect 144208 578866 144528 578898
rect 174928 579454 175248 579486
rect 174928 579218 174970 579454
rect 175206 579218 175248 579454
rect 174928 579134 175248 579218
rect 174928 578898 174970 579134
rect 175206 578898 175248 579134
rect 174928 578866 175248 578898
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 549954 135854 568338
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 135234 549718 135266 549954
rect 135502 549718 135586 549954
rect 135822 549718 135854 549954
rect 135234 549634 135854 549718
rect 135234 549398 135266 549634
rect 135502 549398 135586 549634
rect 135822 549398 135854 549634
rect 135234 542000 135854 549398
rect 138954 553674 139574 558000
rect 138954 553438 138986 553674
rect 139222 553438 139306 553674
rect 139542 553438 139574 553674
rect 138954 553354 139574 553438
rect 138954 553118 138986 553354
rect 139222 553118 139306 553354
rect 139542 553118 139574 553354
rect 138954 542000 139574 553118
rect 145794 543454 146414 558000
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 542000 146414 542898
rect 149514 547174 150134 558000
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 542000 150134 546618
rect 153234 550894 153854 558000
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 542000 153854 550338
rect 156954 554614 157574 558000
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 542000 157574 554058
rect 163794 544394 164414 558000
rect 163794 544158 163826 544394
rect 164062 544158 164146 544394
rect 164382 544158 164414 544394
rect 163794 544074 164414 544158
rect 163794 543838 163826 544074
rect 164062 543838 164146 544074
rect 164382 543838 164414 544074
rect 163794 542000 164414 543838
rect 167514 548114 168134 558000
rect 167514 547878 167546 548114
rect 167782 547878 167866 548114
rect 168102 547878 168134 548114
rect 167514 547794 168134 547878
rect 167514 547558 167546 547794
rect 167782 547558 167866 547794
rect 168102 547558 168134 547794
rect 167514 542000 168134 547558
rect 171234 549954 171854 558000
rect 171234 549718 171266 549954
rect 171502 549718 171586 549954
rect 171822 549718 171854 549954
rect 171234 549634 171854 549718
rect 171234 549398 171266 549634
rect 171502 549398 171586 549634
rect 171822 549398 171854 549634
rect 171234 542000 171854 549398
rect 174954 553674 175574 558000
rect 174954 553438 174986 553674
rect 175222 553438 175306 553674
rect 175542 553438 175574 553674
rect 174954 553354 175574 553438
rect 174954 553118 174986 553354
rect 175222 553118 175306 553354
rect 175542 553118 175574 553354
rect 174954 542000 175574 553118
rect 181794 543454 182414 558000
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 542000 182414 542898
rect 185514 547174 186134 558000
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 542000 186134 546618
rect 189234 550894 189854 558000
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 542000 189854 550338
rect 192954 554614 193574 558000
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 542000 193574 554058
rect 199794 544394 200414 558000
rect 199794 544158 199826 544394
rect 200062 544158 200146 544394
rect 200382 544158 200414 544394
rect 199794 544074 200414 544158
rect 199794 543838 199826 544074
rect 200062 543838 200146 544074
rect 200382 543838 200414 544074
rect 199794 542000 200414 543838
rect 203514 548114 204134 564618
rect 203514 547878 203546 548114
rect 203782 547878 203866 548114
rect 204102 547878 204134 548114
rect 203514 547794 204134 547878
rect 203514 547558 203546 547794
rect 203782 547558 203866 547794
rect 204102 547558 204134 547794
rect 203514 542000 204134 547558
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 549954 207854 568338
rect 207234 549718 207266 549954
rect 207502 549718 207586 549954
rect 207822 549718 207854 549954
rect 207234 549634 207854 549718
rect 207234 549398 207266 549634
rect 207502 549398 207586 549634
rect 207822 549398 207854 549634
rect 207234 542000 207854 549398
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 625099 218414 650898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 625099 222134 654618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 625099 225854 658338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 625099 229574 626058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 625099 236414 632898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 625099 240134 636618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 625099 243854 640338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 625099 247574 644058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 625099 254414 650898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 625099 258134 654618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 625099 261854 658338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 625099 265574 626058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 625099 272414 632898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 625099 276134 636618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 625099 279854 640338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 280659 633452 280725 633453
rect 280659 633388 280660 633452
rect 280724 633388 280725 633452
rect 280659 633387 280725 633388
rect 224208 615454 224528 615486
rect 224208 615218 224250 615454
rect 224486 615218 224528 615454
rect 224208 615134 224528 615218
rect 224208 614898 224250 615134
rect 224486 614898 224528 615134
rect 224208 614866 224528 614898
rect 254928 615454 255248 615486
rect 254928 615218 254970 615454
rect 255206 615218 255248 615454
rect 254928 615134 255248 615218
rect 254928 614898 254970 615134
rect 255206 614898 255248 615134
rect 254928 614866 255248 614898
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 239568 597454 239888 597486
rect 239568 597218 239610 597454
rect 239846 597218 239888 597454
rect 239568 597134 239888 597218
rect 239568 596898 239610 597134
rect 239846 596898 239888 597134
rect 239568 596866 239888 596898
rect 270288 597454 270608 597486
rect 270288 597218 270330 597454
rect 270566 597218 270608 597454
rect 270288 597134 270608 597218
rect 270288 596898 270330 597134
rect 270566 596898 270608 597134
rect 270288 596866 270608 596898
rect 224208 579454 224528 579486
rect 224208 579218 224250 579454
rect 224486 579218 224528 579454
rect 224208 579134 224528 579218
rect 224208 578898 224250 579134
rect 224486 578898 224528 579134
rect 224208 578866 224528 578898
rect 254928 579454 255248 579486
rect 254928 579218 254970 579454
rect 255206 579218 255248 579454
rect 254928 579134 255248 579218
rect 254928 578898 254970 579134
rect 255206 578898 255248 579134
rect 254928 578866 255248 578898
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 553674 211574 572058
rect 210954 553438 210986 553674
rect 211222 553438 211306 553674
rect 211542 553438 211574 553674
rect 210954 553354 211574 553438
rect 210954 553118 210986 553354
rect 211222 553118 211306 553354
rect 211542 553118 211574 553354
rect 210954 542000 211574 553118
rect 217794 543454 218414 558000
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 542000 218414 542898
rect 221514 547174 222134 558000
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 542000 222134 546618
rect 225234 550894 225854 558000
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 542000 225854 550338
rect 228954 554614 229574 558000
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 542000 229574 554058
rect 235794 544394 236414 558000
rect 235794 544158 235826 544394
rect 236062 544158 236146 544394
rect 236382 544158 236414 544394
rect 235794 544074 236414 544158
rect 235794 543838 235826 544074
rect 236062 543838 236146 544074
rect 236382 543838 236414 544074
rect 235794 542000 236414 543838
rect 239514 548114 240134 558000
rect 239514 547878 239546 548114
rect 239782 547878 239866 548114
rect 240102 547878 240134 548114
rect 239514 547794 240134 547878
rect 239514 547558 239546 547794
rect 239782 547558 239866 547794
rect 240102 547558 240134 547794
rect 239514 542000 240134 547558
rect 243234 549954 243854 558000
rect 243234 549718 243266 549954
rect 243502 549718 243586 549954
rect 243822 549718 243854 549954
rect 243234 549634 243854 549718
rect 243234 549398 243266 549634
rect 243502 549398 243586 549634
rect 243822 549398 243854 549634
rect 243234 542000 243854 549398
rect 246954 553674 247574 558000
rect 246954 553438 246986 553674
rect 247222 553438 247306 553674
rect 247542 553438 247574 553674
rect 246954 553354 247574 553438
rect 246954 553118 246986 553354
rect 247222 553118 247306 553354
rect 247542 553118 247574 553354
rect 246954 542000 247574 553118
rect 253794 543454 254414 558000
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 542000 254414 542898
rect 257514 547174 258134 558000
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 542000 258134 546618
rect 261234 550894 261854 558000
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 542000 261854 550338
rect 264954 554614 265574 558000
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 542000 265574 554058
rect 271794 544394 272414 558000
rect 271794 544158 271826 544394
rect 272062 544158 272146 544394
rect 272382 544158 272414 544394
rect 271794 544074 272414 544158
rect 271794 543838 271826 544074
rect 272062 543838 272146 544074
rect 272382 543838 272414 544074
rect 271794 542000 272414 543838
rect 275514 548114 276134 558000
rect 275514 547878 275546 548114
rect 275782 547878 275866 548114
rect 276102 547878 276134 548114
rect 275514 547794 276134 547878
rect 275514 547558 275546 547794
rect 275782 547558 275866 547794
rect 276102 547558 276134 547794
rect 275514 542000 276134 547558
rect 279234 549954 279854 558000
rect 279234 549718 279266 549954
rect 279502 549718 279586 549954
rect 279822 549718 279854 549954
rect 279234 549634 279854 549718
rect 279234 549398 279266 549634
rect 279502 549398 279586 549634
rect 279822 549398 279854 549634
rect 279234 542000 279854 549398
rect 280662 543013 280722 633387
rect 282954 625099 283574 644058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 282954 553674 283574 558000
rect 282954 553438 282986 553674
rect 283222 553438 283306 553674
rect 283542 553438 283574 553674
rect 282954 553354 283574 553438
rect 282954 553118 282986 553354
rect 283222 553118 283306 553354
rect 283542 553118 283574 553354
rect 280659 543012 280725 543013
rect 280659 542948 280660 543012
rect 280724 542948 280725 543012
rect 280659 542947 280725 542948
rect 282954 542000 283574 553118
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 542000 290414 542898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 542000 294134 546618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 542000 297854 550338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 299979 542604 300045 542605
rect 299979 542540 299980 542604
rect 300044 542540 300045 542604
rect 299979 542539 300045 542540
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 79568 525454 79888 525486
rect 79568 525218 79610 525454
rect 79846 525218 79888 525454
rect 79568 525134 79888 525218
rect 79568 524898 79610 525134
rect 79846 524898 79888 525134
rect 79568 524866 79888 524898
rect 110288 525454 110608 525486
rect 110288 525218 110330 525454
rect 110566 525218 110608 525454
rect 110288 525134 110608 525218
rect 110288 524898 110330 525134
rect 110566 524898 110608 525134
rect 110288 524866 110608 524898
rect 141008 525454 141328 525486
rect 141008 525218 141050 525454
rect 141286 525218 141328 525454
rect 141008 525134 141328 525218
rect 141008 524898 141050 525134
rect 141286 524898 141328 525134
rect 141008 524866 141328 524898
rect 171728 525454 172048 525486
rect 171728 525218 171770 525454
rect 172006 525218 172048 525454
rect 171728 525134 172048 525218
rect 171728 524898 171770 525134
rect 172006 524898 172048 525134
rect 171728 524866 172048 524898
rect 202448 525454 202768 525486
rect 202448 525218 202490 525454
rect 202726 525218 202768 525454
rect 202448 525134 202768 525218
rect 202448 524898 202490 525134
rect 202726 524898 202768 525134
rect 202448 524866 202768 524898
rect 233168 525454 233488 525486
rect 233168 525218 233210 525454
rect 233446 525218 233488 525454
rect 233168 525134 233488 525218
rect 233168 524898 233210 525134
rect 233446 524898 233488 525134
rect 233168 524866 233488 524898
rect 263888 525454 264208 525486
rect 263888 525218 263930 525454
rect 264166 525218 264208 525454
rect 263888 525134 264208 525218
rect 263888 524898 263930 525134
rect 264166 524898 264208 525134
rect 263888 524866 264208 524898
rect 294608 525454 294928 525486
rect 294608 525218 294650 525454
rect 294886 525218 294928 525454
rect 294608 525134 294928 525218
rect 294608 524898 294650 525134
rect 294886 524898 294928 525134
rect 294608 524866 294928 524898
rect 299982 517309 300042 542539
rect 300954 542000 301574 554058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 299979 517308 300045 517309
rect 299979 517244 299980 517308
rect 300044 517244 300045 517308
rect 299979 517243 300045 517244
rect 64208 507454 64528 507486
rect 64208 507218 64250 507454
rect 64486 507218 64528 507454
rect 64208 507134 64528 507218
rect 64208 506898 64250 507134
rect 64486 506898 64528 507134
rect 64208 506866 64528 506898
rect 94928 507454 95248 507486
rect 94928 507218 94970 507454
rect 95206 507218 95248 507454
rect 94928 507134 95248 507218
rect 94928 506898 94970 507134
rect 95206 506898 95248 507134
rect 94928 506866 95248 506898
rect 125648 507454 125968 507486
rect 125648 507218 125690 507454
rect 125926 507218 125968 507454
rect 125648 507134 125968 507218
rect 125648 506898 125690 507134
rect 125926 506898 125968 507134
rect 125648 506866 125968 506898
rect 156368 507454 156688 507486
rect 156368 507218 156410 507454
rect 156646 507218 156688 507454
rect 156368 507134 156688 507218
rect 156368 506898 156410 507134
rect 156646 506898 156688 507134
rect 156368 506866 156688 506898
rect 187088 507454 187408 507486
rect 187088 507218 187130 507454
rect 187366 507218 187408 507454
rect 187088 507134 187408 507218
rect 187088 506898 187130 507134
rect 187366 506898 187408 507134
rect 187088 506866 187408 506898
rect 217808 507454 218128 507486
rect 217808 507218 217850 507454
rect 218086 507218 218128 507454
rect 217808 507134 218128 507218
rect 217808 506898 217850 507134
rect 218086 506898 218128 507134
rect 217808 506866 218128 506898
rect 248528 507454 248848 507486
rect 248528 507218 248570 507454
rect 248806 507218 248848 507454
rect 248528 507134 248848 507218
rect 248528 506898 248570 507134
rect 248806 506898 248848 507134
rect 248528 506866 248848 506898
rect 279248 507454 279568 507486
rect 279248 507218 279290 507454
rect 279526 507218 279568 507454
rect 279248 507134 279568 507218
rect 279248 506898 279290 507134
rect 279526 506898 279568 507134
rect 279248 506866 279568 506898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55075 478820 55141 478821
rect 55075 478756 55076 478820
rect 55140 478756 55141 478820
rect 55075 478755 55141 478756
rect 54891 478684 54957 478685
rect 54891 478620 54892 478684
rect 54956 478620 54957 478684
rect 54891 478619 54957 478620
rect 54707 478412 54773 478413
rect 54707 478348 54708 478412
rect 54772 478348 54773 478412
rect 54707 478347 54773 478348
rect 54339 305012 54405 305013
rect 54339 304948 54340 305012
rect 54404 304948 54405 305012
rect 54339 304947 54405 304948
rect 54710 59125 54770 478347
rect 54707 59124 54773 59125
rect 54707 59060 54708 59124
rect 54772 59060 54773 59124
rect 54707 59059 54773 59060
rect 54894 56677 54954 478619
rect 55078 57629 55138 478755
rect 55443 478548 55509 478549
rect 55443 478484 55444 478548
rect 55508 478484 55509 478548
rect 55443 478483 55509 478484
rect 55446 375325 55506 478483
rect 55627 460596 55693 460597
rect 55627 460532 55628 460596
rect 55692 460532 55693 460596
rect 55627 460531 55693 460532
rect 55443 375324 55509 375325
rect 55443 375260 55444 375324
rect 55508 375260 55509 375324
rect 55443 375259 55509 375260
rect 55075 57628 55141 57629
rect 55075 57564 55076 57628
rect 55140 57564 55141 57628
rect 55075 57563 55141 57564
rect 54891 56676 54957 56677
rect 54891 56612 54892 56676
rect 54956 56612 54957 56676
rect 54891 56611 54957 56612
rect 53603 56540 53669 56541
rect 53603 56476 53604 56540
rect 53668 56476 53669 56540
rect 53603 56475 53669 56476
rect 55630 56405 55690 460531
rect 55794 453454 56414 488898
rect 79568 489454 79888 489486
rect 79568 489218 79610 489454
rect 79846 489218 79888 489454
rect 79568 489134 79888 489218
rect 79568 488898 79610 489134
rect 79846 488898 79888 489134
rect 79568 488866 79888 488898
rect 110288 489454 110608 489486
rect 110288 489218 110330 489454
rect 110566 489218 110608 489454
rect 110288 489134 110608 489218
rect 110288 488898 110330 489134
rect 110566 488898 110608 489134
rect 110288 488866 110608 488898
rect 141008 489454 141328 489486
rect 141008 489218 141050 489454
rect 141286 489218 141328 489454
rect 141008 489134 141328 489218
rect 141008 488898 141050 489134
rect 141286 488898 141328 489134
rect 141008 488866 141328 488898
rect 171728 489454 172048 489486
rect 171728 489218 171770 489454
rect 172006 489218 172048 489454
rect 171728 489134 172048 489218
rect 171728 488898 171770 489134
rect 172006 488898 172048 489134
rect 171728 488866 172048 488898
rect 202448 489454 202768 489486
rect 202448 489218 202490 489454
rect 202726 489218 202768 489454
rect 202448 489134 202768 489218
rect 202448 488898 202490 489134
rect 202726 488898 202768 489134
rect 202448 488866 202768 488898
rect 233168 489454 233488 489486
rect 233168 489218 233210 489454
rect 233446 489218 233488 489454
rect 233168 489134 233488 489218
rect 233168 488898 233210 489134
rect 233446 488898 233488 489134
rect 233168 488866 233488 488898
rect 263888 489454 264208 489486
rect 263888 489218 263930 489454
rect 264166 489218 264208 489454
rect 263888 489134 264208 489218
rect 263888 488898 263930 489134
rect 264166 488898 264208 489134
rect 263888 488866 264208 488898
rect 294608 489454 294928 489486
rect 294608 489218 294650 489454
rect 294886 489218 294928 489454
rect 294608 489134 294928 489218
rect 294608 488898 294650 489134
rect 294886 488898 294928 489134
rect 294608 488866 294928 488898
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 208899 479636 208965 479637
rect 208899 479572 208900 479636
rect 208964 479572 208965 479636
rect 208899 479571 208965 479572
rect 206139 479500 206205 479501
rect 206139 479436 206140 479500
rect 206204 479436 206205 479500
rect 206139 479435 206205 479436
rect 198779 478956 198845 478957
rect 198779 478892 198780 478956
rect 198844 478892 198845 478956
rect 198779 478891 198845 478892
rect 198227 478820 198293 478821
rect 198227 478756 198228 478820
rect 198292 478756 198293 478820
rect 198227 478755 198293 478756
rect 196571 478684 196637 478685
rect 196571 478620 196572 478684
rect 196636 478620 196637 478684
rect 196571 478619 196637 478620
rect 59307 478004 59373 478005
rect 59307 477940 59308 478004
rect 59372 477940 59373 478004
rect 59307 477939 59373 477940
rect 57099 475828 57165 475829
rect 57099 475764 57100 475828
rect 57164 475764 57165 475828
rect 57099 475763 57165 475764
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 56547 415308 56613 415309
rect 56547 415244 56548 415308
rect 56612 415244 56613 415308
rect 56547 415243 56613 415244
rect 56550 407829 56610 415243
rect 56547 407828 56613 407829
rect 56547 407764 56548 407828
rect 56612 407764 56613 407828
rect 56547 407763 56613 407764
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 57102 372877 57162 475763
rect 57283 472700 57349 472701
rect 57283 472636 57284 472700
rect 57348 472636 57349 472700
rect 57283 472635 57349 472636
rect 57099 372876 57165 372877
rect 57099 372812 57100 372876
rect 57164 372812 57165 372876
rect 57099 372811 57165 372812
rect 57286 372741 57346 472635
rect 57835 465764 57901 465765
rect 57835 465700 57836 465764
rect 57900 465700 57901 465764
rect 57835 465699 57901 465700
rect 57283 372740 57349 372741
rect 57283 372676 57284 372740
rect 57348 372676 57349 372740
rect 57283 372675 57349 372676
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 57838 267613 57898 465699
rect 59123 461684 59189 461685
rect 59123 461620 59124 461684
rect 59188 461620 59189 461684
rect 59123 461619 59189 461620
rect 58571 459100 58637 459101
rect 58571 459036 58572 459100
rect 58636 459036 58637 459100
rect 58571 459035 58637 459036
rect 57835 267612 57901 267613
rect 57835 267548 57836 267612
rect 57900 267548 57901 267612
rect 57835 267547 57901 267548
rect 57099 262308 57165 262309
rect 57099 262244 57100 262308
rect 57164 262244 57165 262308
rect 57099 262243 57165 262244
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 57102 151830 57162 262243
rect 57835 160172 57901 160173
rect 57835 160108 57836 160172
rect 57900 160108 57901 160172
rect 57835 160107 57901 160108
rect 57102 151770 57346 151830
rect 57286 147525 57346 151770
rect 57283 147524 57349 147525
rect 57283 147460 57284 147524
rect 57348 147460 57349 147524
rect 57283 147459 57349 147460
rect 57099 144804 57165 144805
rect 57099 144740 57100 144804
rect 57164 144740 57165 144804
rect 57099 144739 57165 144740
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 57102 59533 57162 144739
rect 57286 142170 57346 147459
rect 57651 145756 57717 145757
rect 57651 145692 57652 145756
rect 57716 145692 57717 145756
rect 57651 145691 57717 145692
rect 57654 144805 57714 145691
rect 57651 144804 57717 144805
rect 57651 144740 57652 144804
rect 57716 144740 57717 144804
rect 57651 144739 57717 144740
rect 57286 142110 57714 142170
rect 57467 140860 57533 140861
rect 57467 140796 57468 140860
rect 57532 140796 57533 140860
rect 57467 140795 57533 140796
rect 57099 59532 57165 59533
rect 57099 59468 57100 59532
rect 57164 59468 57165 59532
rect 57099 59467 57165 59468
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55627 56404 55693 56405
rect 55627 56340 55628 56404
rect 55692 56340 55693 56404
rect 55627 56339 55693 56340
rect 50843 55044 50909 55045
rect 50843 54980 50844 55044
rect 50908 54980 50909 55044
rect 50843 54979 50909 54980
rect 50659 54908 50725 54909
rect 50659 54844 50660 54908
rect 50724 54844 50725 54908
rect 50659 54843 50725 54844
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 21454 56414 56898
rect 57470 54773 57530 140795
rect 57654 56269 57714 142110
rect 57651 56268 57717 56269
rect 57651 56204 57652 56268
rect 57716 56204 57717 56268
rect 57651 56203 57717 56204
rect 57467 54772 57533 54773
rect 57467 54708 57468 54772
rect 57532 54708 57533 54772
rect 57467 54707 57533 54708
rect 57838 54637 57898 160107
rect 58574 57085 58634 459035
rect 58939 458964 59005 458965
rect 58939 458900 58940 458964
rect 59004 458900 59005 458964
rect 58939 458899 59005 458900
rect 58755 458828 58821 458829
rect 58755 458764 58756 458828
rect 58820 458764 58821 458828
rect 58755 458763 58821 458764
rect 58758 57357 58818 458763
rect 58942 57493 59002 458899
rect 58939 57492 59005 57493
rect 58939 57428 58940 57492
rect 59004 57428 59005 57492
rect 58939 57427 59005 57428
rect 58755 57356 58821 57357
rect 58755 57292 58756 57356
rect 58820 57292 58821 57356
rect 58755 57291 58821 57292
rect 59126 57221 59186 461619
rect 59310 58717 59370 477939
rect 59514 474234 60134 478000
rect 59514 473998 59546 474234
rect 59782 473998 59866 474234
rect 60102 473998 60134 474234
rect 59514 473914 60134 473998
rect 59514 473678 59546 473914
rect 59782 473678 59866 473914
rect 60102 473678 60134 473914
rect 59514 460308 60134 473678
rect 63234 470078 63854 478000
rect 63234 469842 63266 470078
rect 63502 469842 63586 470078
rect 63822 469842 63854 470078
rect 63234 469758 63854 469842
rect 63234 469522 63266 469758
rect 63502 469522 63586 469758
rect 63822 469522 63854 469758
rect 60227 461548 60293 461549
rect 60227 461484 60228 461548
rect 60292 461484 60293 461548
rect 60227 461483 60293 461484
rect 60230 458690 60290 461483
rect 63234 460308 63854 469522
rect 66954 464614 67574 478000
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 460308 67574 464058
rect 73794 471454 74414 478000
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 460308 74414 470898
rect 77514 475174 78134 478000
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 460308 78134 474618
rect 81234 469138 81854 478000
rect 81234 468902 81266 469138
rect 81502 468902 81586 469138
rect 81822 468902 81854 469138
rect 81234 468818 81854 468902
rect 81234 468582 81266 468818
rect 81502 468582 81586 468818
rect 81822 468582 81854 468818
rect 81234 460308 81854 468582
rect 84954 465554 85574 478000
rect 84954 465318 84986 465554
rect 85222 465318 85306 465554
rect 85542 465318 85574 465554
rect 84954 465234 85574 465318
rect 84954 464998 84986 465234
rect 85222 464998 85306 465234
rect 85542 464998 85574 465234
rect 84954 460308 85574 464998
rect 91794 470514 92414 478000
rect 91794 470278 91826 470514
rect 92062 470278 92146 470514
rect 92382 470278 92414 470514
rect 91794 470194 92414 470278
rect 91794 469958 91826 470194
rect 92062 469958 92146 470194
rect 92382 469958 92414 470194
rect 91794 460308 92414 469958
rect 95514 474234 96134 478000
rect 95514 473998 95546 474234
rect 95782 473998 95866 474234
rect 96102 473998 96134 474234
rect 95514 473914 96134 473998
rect 95514 473678 95546 473914
rect 95782 473678 95866 473914
rect 96102 473678 96134 473914
rect 95514 460308 96134 473678
rect 99234 470078 99854 478000
rect 99234 469842 99266 470078
rect 99502 469842 99586 470078
rect 99822 469842 99854 470078
rect 99234 469758 99854 469842
rect 99234 469522 99266 469758
rect 99502 469522 99586 469758
rect 99822 469522 99854 469758
rect 99234 460308 99854 469522
rect 102954 464614 103574 478000
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 460308 103574 464058
rect 109794 471454 110414 478000
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 460308 110414 470898
rect 113514 475174 114134 478000
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 460308 114134 474618
rect 117234 469138 117854 478000
rect 117234 468902 117266 469138
rect 117502 468902 117586 469138
rect 117822 468902 117854 469138
rect 117234 468818 117854 468902
rect 117234 468582 117266 468818
rect 117502 468582 117586 468818
rect 117822 468582 117854 468818
rect 117234 460308 117854 468582
rect 120954 465554 121574 478000
rect 120954 465318 120986 465554
rect 121222 465318 121306 465554
rect 121542 465318 121574 465554
rect 120954 465234 121574 465318
rect 120954 464998 120986 465234
rect 121222 464998 121306 465234
rect 121542 464998 121574 465234
rect 120954 460308 121574 464998
rect 127794 470514 128414 478000
rect 127794 470278 127826 470514
rect 128062 470278 128146 470514
rect 128382 470278 128414 470514
rect 127794 470194 128414 470278
rect 127794 469958 127826 470194
rect 128062 469958 128146 470194
rect 128382 469958 128414 470194
rect 127794 460308 128414 469958
rect 131514 474234 132134 478000
rect 131514 473998 131546 474234
rect 131782 473998 131866 474234
rect 132102 473998 132134 474234
rect 131514 473914 132134 473998
rect 131514 473678 131546 473914
rect 131782 473678 131866 473914
rect 132102 473678 132134 473914
rect 131514 460308 132134 473678
rect 135234 470078 135854 478000
rect 135234 469842 135266 470078
rect 135502 469842 135586 470078
rect 135822 469842 135854 470078
rect 135234 469758 135854 469842
rect 135234 469522 135266 469758
rect 135502 469522 135586 469758
rect 135822 469522 135854 469758
rect 135234 460308 135854 469522
rect 138954 464614 139574 478000
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 460308 139574 464058
rect 145794 471454 146414 478000
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 460308 146414 470898
rect 149514 475174 150134 478000
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 460308 150134 474618
rect 153234 469138 153854 478000
rect 153234 468902 153266 469138
rect 153502 468902 153586 469138
rect 153822 468902 153854 469138
rect 153234 468818 153854 468902
rect 153234 468582 153266 468818
rect 153502 468582 153586 468818
rect 153822 468582 153854 468818
rect 153234 460308 153854 468582
rect 156954 465554 157574 478000
rect 156954 465318 156986 465554
rect 157222 465318 157306 465554
rect 157542 465318 157574 465554
rect 156954 465234 157574 465318
rect 156954 464998 156986 465234
rect 157222 464998 157306 465234
rect 157542 464998 157574 465234
rect 156954 460308 157574 464998
rect 163794 470514 164414 478000
rect 163794 470278 163826 470514
rect 164062 470278 164146 470514
rect 164382 470278 164414 470514
rect 163794 470194 164414 470278
rect 163794 469958 163826 470194
rect 164062 469958 164146 470194
rect 164382 469958 164414 470194
rect 163794 460308 164414 469958
rect 167514 474234 168134 478000
rect 167514 473998 167546 474234
rect 167782 473998 167866 474234
rect 168102 473998 168134 474234
rect 167514 473914 168134 473998
rect 167514 473678 167546 473914
rect 167782 473678 167866 473914
rect 168102 473678 168134 473914
rect 167514 460308 168134 473678
rect 171234 470078 171854 478000
rect 171234 469842 171266 470078
rect 171502 469842 171586 470078
rect 171822 469842 171854 470078
rect 171234 469758 171854 469842
rect 171234 469522 171266 469758
rect 171502 469522 171586 469758
rect 171822 469522 171854 469758
rect 171234 460308 171854 469522
rect 174954 464614 175574 478000
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 460308 175574 464058
rect 181794 471454 182414 478000
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 179643 461684 179709 461685
rect 179643 461620 179644 461684
rect 179708 461620 179709 461684
rect 179643 461619 179709 461620
rect 178355 461412 178421 461413
rect 178355 461348 178356 461412
rect 178420 461348 178421 461412
rect 178355 461347 178421 461348
rect 59862 458630 60290 458690
rect 178358 458690 178418 461347
rect 179646 458690 179706 461619
rect 181794 460308 182414 470898
rect 185514 475174 186134 478000
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 460308 186134 474618
rect 189234 469138 189854 478000
rect 189234 468902 189266 469138
rect 189502 468902 189586 469138
rect 189822 468902 189854 469138
rect 189234 468818 189854 468902
rect 189234 468582 189266 468818
rect 189502 468582 189586 468818
rect 189822 468582 189854 468818
rect 189234 460308 189854 468582
rect 192954 465554 193574 478000
rect 192954 465318 192986 465554
rect 193222 465318 193306 465554
rect 193542 465318 193574 465554
rect 192954 465234 193574 465318
rect 192954 464998 192986 465234
rect 193222 464998 193306 465234
rect 193542 464998 193574 465234
rect 190867 461004 190933 461005
rect 190867 460940 190868 461004
rect 190932 460940 190933 461004
rect 190867 460939 190933 460940
rect 190870 458690 190930 460939
rect 192954 460308 193574 464998
rect 178358 458630 178524 458690
rect 179646 458630 179748 458690
rect 59862 374010 59922 458630
rect 178464 458202 178524 458630
rect 179688 458202 179748 458630
rect 190840 458630 190930 458690
rect 190840 458202 190900 458630
rect 60272 453454 60620 453486
rect 60272 453218 60328 453454
rect 60564 453218 60620 453454
rect 60272 453134 60620 453218
rect 60272 452898 60328 453134
rect 60564 452898 60620 453134
rect 60272 452866 60620 452898
rect 196000 453454 196348 453486
rect 196000 453218 196056 453454
rect 196292 453218 196348 453454
rect 196000 453134 196348 453218
rect 196000 452898 196056 453134
rect 196292 452898 196348 453134
rect 196000 452866 196348 452898
rect 60952 435454 61300 435486
rect 60952 435218 61008 435454
rect 61244 435218 61300 435454
rect 60952 435134 61300 435218
rect 60952 434898 61008 435134
rect 61244 434898 61300 435134
rect 60952 434866 61300 434898
rect 195320 435454 195668 435486
rect 195320 435218 195376 435454
rect 195612 435218 195668 435454
rect 195320 435134 195668 435218
rect 195320 434898 195376 435134
rect 195612 434898 195668 435134
rect 195320 434866 195668 434898
rect 60272 417454 60620 417486
rect 60272 417218 60328 417454
rect 60564 417218 60620 417454
rect 60272 417134 60620 417218
rect 60272 416898 60328 417134
rect 60564 416898 60620 417134
rect 60272 416866 60620 416898
rect 196000 417454 196348 417486
rect 196000 417218 196056 417454
rect 196292 417218 196348 417454
rect 196000 417134 196348 417218
rect 196000 416898 196056 417134
rect 196292 416898 196348 417134
rect 196000 416866 196348 416898
rect 60952 399454 61300 399486
rect 60952 399218 61008 399454
rect 61244 399218 61300 399454
rect 60952 399134 61300 399218
rect 60952 398898 61008 399134
rect 61244 398898 61300 399134
rect 60952 398866 61300 398898
rect 195320 399454 195668 399486
rect 195320 399218 195376 399454
rect 195612 399218 195668 399454
rect 195320 399134 195668 399218
rect 195320 398898 195376 399134
rect 195612 398898 195668 399134
rect 195320 398866 195668 398898
rect 60272 381454 60620 381486
rect 60272 381218 60328 381454
rect 60564 381218 60620 381454
rect 60272 381134 60620 381218
rect 60272 380898 60328 381134
rect 60564 380898 60620 381134
rect 60272 380866 60620 380898
rect 196000 381454 196348 381486
rect 196000 381218 196056 381454
rect 196292 381218 196348 381454
rect 196000 381134 196348 381218
rect 196000 380898 196056 381134
rect 196292 380898 196348 381134
rect 196000 380866 196348 380898
rect 76086 374990 76666 375050
rect 59862 373950 60290 374010
rect 59514 366234 60134 373000
rect 59514 365998 59546 366234
rect 59782 365998 59866 366234
rect 60102 365998 60134 366234
rect 59514 365914 60134 365998
rect 59514 365678 59546 365914
rect 59782 365678 59866 365914
rect 60102 365678 60134 365914
rect 59514 355308 60134 365678
rect 60230 354690 60290 373950
rect 63234 369954 63854 373000
rect 63234 369718 63266 369954
rect 63502 369718 63586 369954
rect 63822 369718 63854 369954
rect 63234 369634 63854 369718
rect 63234 369398 63266 369634
rect 63502 369398 63586 369634
rect 63822 369398 63854 369634
rect 63234 355308 63854 369398
rect 66954 356614 67574 373000
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 355308 67574 356058
rect 73794 363454 74414 373000
rect 76606 372197 76666 374990
rect 77158 372605 77218 375050
rect 78262 374990 78506 375050
rect 79622 374990 79978 375050
rect 77155 372604 77221 372605
rect 77155 372540 77156 372604
rect 77220 372540 77221 372604
rect 77155 372539 77221 372540
rect 76603 372196 76669 372197
rect 76603 372132 76604 372196
rect 76668 372132 76669 372196
rect 76603 372131 76669 372132
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 355308 74414 362898
rect 77514 367174 78134 373000
rect 78446 372469 78506 374990
rect 79918 372469 79978 374990
rect 80470 374990 80574 375050
rect 81798 374990 82002 375050
rect 83158 374990 83842 375050
rect 84246 374990 84578 375050
rect 78443 372468 78509 372469
rect 78443 372404 78444 372468
rect 78508 372404 78509 372468
rect 78443 372403 78509 372404
rect 79915 372468 79981 372469
rect 79915 372404 79916 372468
rect 79980 372404 79981 372468
rect 79915 372403 79981 372404
rect 80470 372333 80530 374990
rect 80467 372332 80533 372333
rect 80467 372268 80468 372332
rect 80532 372268 80533 372332
rect 80467 372267 80533 372268
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 355308 78134 366618
rect 81234 370894 81854 373000
rect 81942 372333 82002 374990
rect 81939 372332 82005 372333
rect 81939 372268 81940 372332
rect 82004 372268 82005 372332
rect 81939 372267 82005 372268
rect 83782 371925 83842 374990
rect 84518 372605 84578 374990
rect 84702 374990 85470 375050
rect 84515 372604 84581 372605
rect 84515 372540 84516 372604
rect 84580 372540 84581 372604
rect 84515 372539 84581 372540
rect 84702 372469 84762 374990
rect 84699 372468 84765 372469
rect 84699 372404 84700 372468
rect 84764 372404 84765 372468
rect 84699 372403 84765 372404
rect 83779 371924 83845 371925
rect 83779 371860 83780 371924
rect 83844 371860 83845 371924
rect 83779 371859 83845 371860
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 355308 81854 370338
rect 84954 357554 85574 373000
rect 86542 372605 86602 375050
rect 87646 374990 88074 375050
rect 88326 374990 88442 375050
rect 88734 374990 89362 375050
rect 88014 372605 88074 374990
rect 88382 373285 88442 374990
rect 88379 373284 88445 373285
rect 88379 373220 88380 373284
rect 88444 373220 88445 373284
rect 88379 373219 88445 373220
rect 89302 372605 89362 374990
rect 90038 372605 90098 375050
rect 90222 374990 90774 375050
rect 91318 374990 91570 375050
rect 92406 374990 92490 375050
rect 90222 373149 90282 374990
rect 90219 373148 90285 373149
rect 90219 373084 90220 373148
rect 90284 373084 90285 373148
rect 90219 373083 90285 373084
rect 91510 372605 91570 374990
rect 92430 373149 92490 374990
rect 93350 374990 93494 375050
rect 93630 374990 93778 375050
rect 94582 374990 95066 375050
rect 92427 373148 92493 373149
rect 92427 373084 92428 373148
rect 92492 373084 92493 373148
rect 92427 373083 92493 373084
rect 86539 372604 86605 372605
rect 86539 372540 86540 372604
rect 86604 372540 86605 372604
rect 86539 372539 86605 372540
rect 88011 372604 88077 372605
rect 88011 372540 88012 372604
rect 88076 372540 88077 372604
rect 88011 372539 88077 372540
rect 89299 372604 89365 372605
rect 89299 372540 89300 372604
rect 89364 372540 89365 372604
rect 89299 372539 89365 372540
rect 90035 372604 90101 372605
rect 90035 372540 90036 372604
rect 90100 372540 90101 372604
rect 90035 372539 90101 372540
rect 91507 372604 91573 372605
rect 91507 372540 91508 372604
rect 91572 372540 91573 372604
rect 91507 372539 91573 372540
rect 84954 357318 84986 357554
rect 85222 357318 85306 357554
rect 85542 357318 85574 357554
rect 84954 357234 85574 357318
rect 84954 356998 84986 357234
rect 85222 356998 85306 357234
rect 85542 356998 85574 357234
rect 84954 355308 85574 356998
rect 91794 364394 92414 373000
rect 93350 372605 93410 374990
rect 93718 373421 93778 374990
rect 95006 373693 95066 374990
rect 95912 374370 95972 375020
rect 96078 374990 96170 375050
rect 97030 374990 97642 375050
rect 98118 374990 98194 375050
rect 95912 374310 95986 374370
rect 95003 373692 95069 373693
rect 95003 373628 95004 373692
rect 95068 373628 95069 373692
rect 95003 373627 95069 373628
rect 93715 373420 93781 373421
rect 93715 373356 93716 373420
rect 93780 373356 93781 373420
rect 93715 373355 93781 373356
rect 95926 373285 95986 374310
rect 96110 373693 96170 374990
rect 96107 373692 96173 373693
rect 96107 373628 96108 373692
rect 96172 373628 96173 373692
rect 96107 373627 96173 373628
rect 95923 373284 95989 373285
rect 95923 373220 95924 373284
rect 95988 373220 95989 373284
rect 95923 373219 95989 373220
rect 93347 372604 93413 372605
rect 93347 372540 93348 372604
rect 93412 372540 93413 372604
rect 93347 372539 93413 372540
rect 91794 364158 91826 364394
rect 92062 364158 92146 364394
rect 92382 364158 92414 364394
rect 91794 364074 92414 364158
rect 91794 363838 91826 364074
rect 92062 363838 92146 364074
rect 92382 363838 92414 364074
rect 91794 355308 92414 363838
rect 95514 366234 96134 373000
rect 97582 371653 97642 374990
rect 98134 371653 98194 374990
rect 98318 374990 98526 375050
rect 99478 374990 100034 375050
rect 100702 374990 100770 375050
rect 98318 373421 98378 374990
rect 98315 373420 98381 373421
rect 98315 373356 98316 373420
rect 98380 373356 98381 373420
rect 98315 373355 98381 373356
rect 97579 371652 97645 371653
rect 97579 371588 97580 371652
rect 97644 371588 97645 371652
rect 97579 371587 97645 371588
rect 98131 371652 98197 371653
rect 98131 371588 98132 371652
rect 98196 371588 98197 371652
rect 98131 371587 98197 371588
rect 95514 365998 95546 366234
rect 95782 365998 95866 366234
rect 96102 365998 96134 366234
rect 95514 365914 96134 365998
rect 95514 365678 95546 365914
rect 95782 365678 95866 365914
rect 96102 365678 96134 365914
rect 95514 355308 96134 365678
rect 99234 369954 99854 373000
rect 99974 371653 100034 374990
rect 99971 371652 100037 371653
rect 99971 371588 99972 371652
rect 100036 371588 100037 371652
rect 99971 371587 100037 371588
rect 100710 371517 100770 374990
rect 100894 374990 101110 375050
rect 101790 374990 102058 375050
rect 100894 373285 100954 374990
rect 100891 373284 100957 373285
rect 100891 373220 100892 373284
rect 100956 373220 100957 373284
rect 100891 373219 100957 373220
rect 101998 372333 102058 374990
rect 102734 374990 102878 375050
rect 103286 374990 103558 375050
rect 103966 374990 104634 375050
rect 102734 372469 102794 374990
rect 103286 373693 103346 374990
rect 103283 373692 103349 373693
rect 103283 373628 103284 373692
rect 103348 373628 103349 373692
rect 103283 373627 103349 373628
rect 102731 372468 102797 372469
rect 102731 372404 102732 372468
rect 102796 372404 102797 372468
rect 102731 372403 102797 372404
rect 101995 372332 102061 372333
rect 101995 372268 101996 372332
rect 102060 372268 102061 372332
rect 101995 372267 102061 372268
rect 100707 371516 100773 371517
rect 100707 371452 100708 371516
rect 100772 371452 100773 371516
rect 100707 371451 100773 371452
rect 99234 369718 99266 369954
rect 99502 369718 99586 369954
rect 99822 369718 99854 369954
rect 99234 369634 99854 369718
rect 99234 369398 99266 369634
rect 99502 369398 99586 369634
rect 99822 369398 99854 369634
rect 99234 355308 99854 369398
rect 102954 356614 103574 373000
rect 104574 371925 104634 374990
rect 104571 371924 104637 371925
rect 104571 371860 104572 371924
rect 104636 371860 104637 371924
rect 104571 371859 104637 371860
rect 105310 371789 105370 375050
rect 105494 374990 106006 375050
rect 106414 374990 107026 375050
rect 105494 374509 105554 374990
rect 105491 374508 105557 374509
rect 105491 374444 105492 374508
rect 105556 374444 105557 374508
rect 105491 374443 105557 374444
rect 105307 371788 105373 371789
rect 105307 371724 105308 371788
rect 105372 371724 105373 371788
rect 105307 371723 105373 371724
rect 106966 371381 107026 374990
rect 107518 374990 107638 375050
rect 107886 374990 108318 375050
rect 108726 374990 108866 375050
rect 107518 371381 107578 374990
rect 107886 373693 107946 374990
rect 107883 373692 107949 373693
rect 107883 373628 107884 373692
rect 107948 373628 107949 373692
rect 107883 373627 107949 373628
rect 108806 372605 108866 374990
rect 109542 374990 109814 375050
rect 110462 374990 111038 375050
rect 111174 374990 111810 375050
rect 112262 374990 112914 375050
rect 108803 372604 108869 372605
rect 108803 372540 108804 372604
rect 108868 372540 108869 372604
rect 108803 372539 108869 372540
rect 109542 372333 109602 374990
rect 110462 373557 110522 374990
rect 110459 373556 110525 373557
rect 110459 373492 110460 373556
rect 110524 373492 110525 373556
rect 110459 373491 110525 373492
rect 109539 372332 109605 372333
rect 109539 372268 109540 372332
rect 109604 372268 109605 372332
rect 109539 372267 109605 372268
rect 106963 371380 107029 371381
rect 106963 371316 106964 371380
rect 107028 371316 107029 371380
rect 106963 371315 107029 371316
rect 107515 371380 107581 371381
rect 107515 371316 107516 371380
rect 107580 371316 107581 371380
rect 107515 371315 107581 371316
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 355308 103574 356058
rect 109794 363454 110414 373000
rect 111750 372197 111810 374990
rect 111747 372196 111813 372197
rect 111747 372132 111748 372196
rect 111812 372132 111813 372196
rect 111747 372131 111813 372132
rect 112854 371925 112914 374990
rect 113222 374990 113350 375050
rect 113222 372605 113282 374990
rect 113592 374370 113652 375020
rect 114438 374990 114570 375050
rect 113590 374310 113652 374370
rect 113590 373693 113650 374310
rect 113587 373692 113653 373693
rect 113587 373628 113588 373692
rect 113652 373628 113653 373692
rect 113587 373627 113653 373628
rect 113219 372604 113285 372605
rect 113219 372540 113220 372604
rect 113284 372540 113285 372604
rect 113219 372539 113285 372540
rect 112851 371924 112917 371925
rect 112851 371860 112852 371924
rect 112916 371860 112917 371924
rect 112851 371859 112917 371860
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 355308 110414 362898
rect 113514 367174 114134 373000
rect 114510 371789 114570 374990
rect 115768 374370 115828 375020
rect 116040 374509 116100 375020
rect 117022 374990 117146 375050
rect 118110 374990 118250 375050
rect 116037 374508 116103 374509
rect 116037 374444 116038 374508
rect 116102 374444 116103 374508
rect 116037 374443 116103 374444
rect 115768 374310 115858 374370
rect 114507 371788 114573 371789
rect 114507 371724 114508 371788
rect 114572 371724 114573 371788
rect 114507 371723 114573 371724
rect 115798 371381 115858 374310
rect 117086 372469 117146 374990
rect 117083 372468 117149 372469
rect 117083 372404 117084 372468
rect 117148 372404 117149 372468
rect 117083 372403 117149 372404
rect 115795 371380 115861 371381
rect 115795 371316 115796 371380
rect 115860 371316 115861 371380
rect 115795 371315 115861 371316
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 355308 114134 366618
rect 117234 370894 117854 373000
rect 118190 372333 118250 374990
rect 118374 374990 118518 375050
rect 119198 374990 119906 375050
rect 120966 374990 121378 375050
rect 123550 374990 124138 375050
rect 118374 373693 118434 374990
rect 118371 373692 118437 373693
rect 118371 373628 118372 373692
rect 118436 373628 118437 373692
rect 118371 373627 118437 373628
rect 119846 373557 119906 374990
rect 121318 373693 121378 374990
rect 121315 373692 121381 373693
rect 121315 373628 121316 373692
rect 121380 373628 121381 373692
rect 121315 373627 121381 373628
rect 124078 373557 124138 374990
rect 125734 374990 125998 375050
rect 128310 374990 128922 375050
rect 131030 374990 131130 375050
rect 133478 374990 133706 375050
rect 135926 374990 136466 375050
rect 138510 374990 139226 375050
rect 125734 373557 125794 374990
rect 128862 373557 128922 374990
rect 131070 373557 131130 374990
rect 133646 373557 133706 374990
rect 136406 373557 136466 374990
rect 139166 374101 139226 374990
rect 140928 374509 140988 375020
rect 143512 374509 143572 375020
rect 145990 374990 146218 375050
rect 148574 374990 148978 375050
rect 151022 374990 151738 375050
rect 153470 374990 154130 375050
rect 155918 374990 156522 375050
rect 140925 374508 140991 374509
rect 140925 374444 140926 374508
rect 140990 374444 140991 374508
rect 140925 374443 140991 374444
rect 143509 374508 143575 374509
rect 143509 374444 143510 374508
rect 143574 374444 143575 374508
rect 143509 374443 143575 374444
rect 146158 374373 146218 374990
rect 148918 374373 148978 374990
rect 146155 374372 146221 374373
rect 146155 374308 146156 374372
rect 146220 374308 146221 374372
rect 146155 374307 146221 374308
rect 148915 374372 148981 374373
rect 148915 374308 148916 374372
rect 148980 374308 148981 374372
rect 148915 374307 148981 374308
rect 139163 374100 139229 374101
rect 139163 374036 139164 374100
rect 139228 374036 139229 374100
rect 139163 374035 139229 374036
rect 151678 373557 151738 374990
rect 154070 373557 154130 374990
rect 156462 374509 156522 374990
rect 158486 374645 158546 375050
rect 158483 374644 158549 374645
rect 158483 374580 158484 374644
rect 158548 374580 158549 374644
rect 158483 374579 158549 374580
rect 160920 374509 160980 375020
rect 163368 374509 163428 375020
rect 165952 374645 166012 375020
rect 183142 374990 183254 375050
rect 165949 374644 166015 374645
rect 165949 374580 165950 374644
rect 166014 374580 166015 374644
rect 165949 374579 166015 374580
rect 156459 374508 156525 374509
rect 156459 374444 156460 374508
rect 156524 374444 156525 374508
rect 156459 374443 156525 374444
rect 160917 374508 160983 374509
rect 160917 374444 160918 374508
rect 160982 374444 160983 374508
rect 160917 374443 160983 374444
rect 163365 374508 163431 374509
rect 163365 374444 163366 374508
rect 163430 374444 163431 374508
rect 163365 374443 163431 374444
rect 119843 373556 119909 373557
rect 119843 373492 119844 373556
rect 119908 373492 119909 373556
rect 119843 373491 119909 373492
rect 124075 373556 124141 373557
rect 124075 373492 124076 373556
rect 124140 373492 124141 373556
rect 124075 373491 124141 373492
rect 125731 373556 125797 373557
rect 125731 373492 125732 373556
rect 125796 373492 125797 373556
rect 125731 373491 125797 373492
rect 128859 373556 128925 373557
rect 128859 373492 128860 373556
rect 128924 373492 128925 373556
rect 128859 373491 128925 373492
rect 131067 373556 131133 373557
rect 131067 373492 131068 373556
rect 131132 373492 131133 373556
rect 131067 373491 131133 373492
rect 133643 373556 133709 373557
rect 133643 373492 133644 373556
rect 133708 373492 133709 373556
rect 133643 373491 133709 373492
rect 136403 373556 136469 373557
rect 136403 373492 136404 373556
rect 136468 373492 136469 373556
rect 136403 373491 136469 373492
rect 151675 373556 151741 373557
rect 151675 373492 151676 373556
rect 151740 373492 151741 373556
rect 151675 373491 151741 373492
rect 154067 373556 154133 373557
rect 154067 373492 154068 373556
rect 154132 373492 154133 373556
rect 154067 373491 154133 373492
rect 118187 372332 118253 372333
rect 118187 372268 118188 372332
rect 118252 372268 118253 372332
rect 118187 372267 118253 372268
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 355308 117854 370338
rect 120954 357554 121574 373000
rect 120954 357318 120986 357554
rect 121222 357318 121306 357554
rect 121542 357318 121574 357554
rect 120954 357234 121574 357318
rect 120954 356998 120986 357234
rect 121222 356998 121306 357234
rect 121542 356998 121574 357234
rect 120954 355308 121574 356998
rect 127794 364394 128414 373000
rect 127794 364158 127826 364394
rect 128062 364158 128146 364394
rect 128382 364158 128414 364394
rect 127794 364074 128414 364158
rect 127794 363838 127826 364074
rect 128062 363838 128146 364074
rect 128382 363838 128414 364074
rect 127794 355308 128414 363838
rect 131514 366234 132134 373000
rect 131514 365998 131546 366234
rect 131782 365998 131866 366234
rect 132102 365998 132134 366234
rect 131514 365914 132134 365998
rect 131514 365678 131546 365914
rect 131782 365678 131866 365914
rect 132102 365678 132134 365914
rect 131514 355308 132134 365678
rect 135234 369954 135854 373000
rect 135234 369718 135266 369954
rect 135502 369718 135586 369954
rect 135822 369718 135854 369954
rect 135234 369634 135854 369718
rect 135234 369398 135266 369634
rect 135502 369398 135586 369634
rect 135822 369398 135854 369634
rect 135234 355308 135854 369398
rect 138954 356614 139574 373000
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 355308 139574 356058
rect 145794 363454 146414 373000
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 355308 146414 362898
rect 149514 367174 150134 373000
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 355308 150134 366618
rect 153234 370894 153854 373000
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 355308 153854 370338
rect 156954 357554 157574 373000
rect 156954 357318 156986 357554
rect 157222 357318 157306 357554
rect 157542 357318 157574 357554
rect 156954 357234 157574 357318
rect 156954 356998 156986 357234
rect 157222 356998 157306 357234
rect 157542 356998 157574 357234
rect 156954 355308 157574 356998
rect 163794 364394 164414 373000
rect 163794 364158 163826 364394
rect 164062 364158 164146 364394
rect 164382 364158 164414 364394
rect 163794 364074 164414 364158
rect 163794 363838 163826 364074
rect 164062 363838 164146 364074
rect 164382 363838 164414 364074
rect 163794 355308 164414 363838
rect 167514 366234 168134 373000
rect 167514 365998 167546 366234
rect 167782 365998 167866 366234
rect 168102 365998 168134 366234
rect 167514 365914 168134 365998
rect 167514 365678 167546 365914
rect 167782 365678 167866 365914
rect 168102 365678 168134 365914
rect 167514 355308 168134 365678
rect 171234 369954 171854 373000
rect 171234 369718 171266 369954
rect 171502 369718 171586 369954
rect 171822 369718 171854 369954
rect 171234 369634 171854 369718
rect 171234 369398 171266 369634
rect 171502 369398 171586 369634
rect 171822 369398 171854 369634
rect 171234 355308 171854 369398
rect 174954 356614 175574 373000
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 355308 175574 356058
rect 181794 363454 182414 373000
rect 183142 372605 183202 374990
rect 183360 374370 183420 375020
rect 183326 374310 183420 374370
rect 183139 372604 183205 372605
rect 183139 372540 183140 372604
rect 183204 372540 183205 372604
rect 183139 372539 183205 372540
rect 183326 371517 183386 374310
rect 183323 371516 183389 371517
rect 183323 371452 183324 371516
rect 183388 371452 183389 371516
rect 183323 371451 183389 371452
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 179643 355332 179709 355333
rect 179643 355268 179644 355332
rect 179708 355268 179709 355332
rect 181794 355308 182414 362898
rect 185514 367174 186134 373000
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 355308 186134 366618
rect 189234 370894 189854 373000
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 355308 189854 370338
rect 192954 357554 193574 373000
rect 192954 357318 192986 357554
rect 193222 357318 193306 357554
rect 193542 357318 193574 357554
rect 192954 357234 193574 357318
rect 192954 356998 192986 357234
rect 193222 356998 193306 357234
rect 193542 356998 193574 357234
rect 190867 355332 190933 355333
rect 179643 355267 179709 355268
rect 190867 355268 190868 355332
rect 190932 355268 190933 355332
rect 192954 355308 193574 356998
rect 190867 355267 190933 355268
rect 178539 354788 178605 354789
rect 178539 354724 178540 354788
rect 178604 354724 178605 354788
rect 178539 354723 178605 354724
rect 59862 354630 60290 354690
rect 59862 268290 59922 354630
rect 178542 353970 178602 354723
rect 178464 353910 178602 353970
rect 179646 353970 179706 355267
rect 190870 353970 190930 355267
rect 179646 353910 179748 353970
rect 178464 353260 178524 353910
rect 179688 353260 179748 353910
rect 190840 353910 190930 353970
rect 190840 353260 190900 353910
rect 60272 345454 60620 345486
rect 60272 345218 60328 345454
rect 60564 345218 60620 345454
rect 60272 345134 60620 345218
rect 60272 344898 60328 345134
rect 60564 344898 60620 345134
rect 60272 344866 60620 344898
rect 196000 345454 196348 345486
rect 196000 345218 196056 345454
rect 196292 345218 196348 345454
rect 196000 345134 196348 345218
rect 196000 344898 196056 345134
rect 196292 344898 196348 345134
rect 196000 344866 196348 344898
rect 60952 327454 61300 327486
rect 60952 327218 61008 327454
rect 61244 327218 61300 327454
rect 60952 327134 61300 327218
rect 60952 326898 61008 327134
rect 61244 326898 61300 327134
rect 60952 326866 61300 326898
rect 195320 327454 195668 327486
rect 195320 327218 195376 327454
rect 195612 327218 195668 327454
rect 195320 327134 195668 327218
rect 195320 326898 195376 327134
rect 195612 326898 195668 327134
rect 195320 326866 195668 326898
rect 60272 309454 60620 309486
rect 60272 309218 60328 309454
rect 60564 309218 60620 309454
rect 60272 309134 60620 309218
rect 60272 308898 60328 309134
rect 60564 308898 60620 309134
rect 60272 308866 60620 308898
rect 196000 309454 196348 309486
rect 196000 309218 196056 309454
rect 196292 309218 196348 309454
rect 196000 309134 196348 309218
rect 196000 308898 196056 309134
rect 196292 308898 196348 309134
rect 196000 308866 196348 308898
rect 60952 291454 61300 291486
rect 60952 291218 61008 291454
rect 61244 291218 61300 291454
rect 60952 291134 61300 291218
rect 60952 290898 61008 291134
rect 61244 290898 61300 291134
rect 60952 290866 61300 290898
rect 195320 291454 195668 291486
rect 195320 291218 195376 291454
rect 195612 291218 195668 291454
rect 195320 291134 195668 291218
rect 195320 290898 195376 291134
rect 195612 290898 195668 291134
rect 195320 290866 195668 290898
rect 60272 273454 60620 273486
rect 60272 273218 60328 273454
rect 60564 273218 60620 273454
rect 60272 273134 60620 273218
rect 60272 272898 60328 273134
rect 60564 272898 60620 273134
rect 60272 272866 60620 272898
rect 196000 273454 196348 273486
rect 196000 273218 196056 273454
rect 196292 273218 196348 273454
rect 196000 273134 196348 273218
rect 196000 272898 196056 273134
rect 196292 272898 196348 273134
rect 196000 272866 196348 272898
rect 76056 269650 76116 270106
rect 76054 269590 76116 269650
rect 77144 269650 77204 270106
rect 78232 269650 78292 270106
rect 79592 269650 79652 270106
rect 80544 269650 80604 270106
rect 77144 269590 77218 269650
rect 78232 269590 78322 269650
rect 76054 268837 76114 269590
rect 77158 268837 77218 269590
rect 76051 268836 76117 268837
rect 76051 268772 76052 268836
rect 76116 268772 76117 268836
rect 76051 268771 76117 268772
rect 77155 268836 77221 268837
rect 77155 268772 77156 268836
rect 77220 268772 77221 268836
rect 77155 268771 77221 268772
rect 59862 268230 60290 268290
rect 59514 260114 60134 268000
rect 59514 259878 59546 260114
rect 59782 259878 59866 260114
rect 60102 259878 60134 260114
rect 59514 259794 60134 259878
rect 59514 259558 59546 259794
rect 59782 259558 59866 259794
rect 60102 259558 60134 259794
rect 59514 250308 60134 259558
rect 60230 248430 60290 268230
rect 63234 261954 63854 268000
rect 63234 261718 63266 261954
rect 63502 261718 63586 261954
rect 63822 261718 63854 261954
rect 63234 261634 63854 261718
rect 63234 261398 63266 261634
rect 63502 261398 63586 261634
rect 63822 261398 63854 261634
rect 63234 250308 63854 261398
rect 66954 265674 67574 268000
rect 66954 265438 66986 265674
rect 67222 265438 67306 265674
rect 67542 265438 67574 265674
rect 66954 265354 67574 265438
rect 66954 265118 66986 265354
rect 67222 265118 67306 265354
rect 67542 265118 67574 265354
rect 66954 250308 67574 265118
rect 73794 255454 74414 268000
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 250308 74414 254898
rect 77514 259174 78134 268000
rect 78262 267069 78322 269590
rect 79550 269590 79652 269650
rect 80470 269590 80604 269650
rect 81768 269650 81828 270106
rect 83128 269653 83188 270106
rect 83125 269652 83191 269653
rect 81768 269590 82002 269650
rect 79550 267069 79610 269590
rect 80470 267477 80530 269590
rect 80467 267476 80533 267477
rect 80467 267412 80468 267476
rect 80532 267412 80533 267476
rect 80467 267411 80533 267412
rect 78259 267068 78325 267069
rect 78259 267004 78260 267068
rect 78324 267004 78325 267068
rect 78259 267003 78325 267004
rect 79547 267068 79613 267069
rect 79547 267004 79548 267068
rect 79612 267004 79613 267068
rect 79547 267003 79613 267004
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 250308 78134 258618
rect 81234 262894 81854 268000
rect 81942 267341 82002 269590
rect 83125 269588 83126 269652
rect 83190 269588 83191 269652
rect 84216 269650 84276 270106
rect 85440 269650 85500 270106
rect 83125 269587 83191 269588
rect 83966 269590 84276 269650
rect 85438 269590 85500 269650
rect 86528 269650 86588 270106
rect 87616 269650 87676 270106
rect 86528 269590 86602 269650
rect 83966 267749 84026 269590
rect 85438 268157 85498 269590
rect 85435 268156 85501 268157
rect 85435 268092 85436 268156
rect 85500 268092 85501 268156
rect 85435 268091 85501 268092
rect 83963 267748 84029 267749
rect 83963 267684 83964 267748
rect 84028 267684 84029 267748
rect 83963 267683 84029 267684
rect 81939 267340 82005 267341
rect 81939 267276 81940 267340
rect 82004 267276 82005 267340
rect 81939 267275 82005 267276
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 250308 81854 262338
rect 84954 266614 85574 268000
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 86542 266389 86602 269590
rect 87462 269590 87676 269650
rect 88296 269650 88356 270106
rect 88704 269650 88764 270106
rect 90064 269650 90124 270106
rect 88296 269590 88442 269650
rect 88704 269590 88810 269650
rect 87462 266389 87522 269590
rect 88382 267069 88442 269590
rect 88379 267068 88445 267069
rect 88379 267004 88380 267068
rect 88444 267004 88445 267068
rect 88379 267003 88445 267004
rect 88750 266389 88810 269590
rect 90038 269590 90124 269650
rect 90744 269650 90804 270106
rect 91288 269653 91348 270106
rect 91285 269652 91351 269653
rect 90744 269590 90834 269650
rect 90038 266389 90098 269590
rect 90774 268837 90834 269590
rect 91285 269588 91286 269652
rect 91350 269588 91351 269652
rect 92376 269650 92436 270106
rect 93464 269650 93524 270106
rect 93600 269653 93660 270106
rect 94552 269653 94612 270106
rect 92376 269590 92490 269650
rect 91285 269587 91351 269588
rect 90771 268836 90837 268837
rect 90771 268772 90772 268836
rect 90836 268772 90837 268836
rect 90771 268771 90837 268772
rect 92430 268157 92490 269590
rect 93350 269590 93524 269650
rect 93597 269652 93663 269653
rect 92427 268156 92493 268157
rect 92427 268092 92428 268156
rect 92492 268092 92493 268156
rect 92427 268091 92493 268092
rect 84954 266294 85574 266378
rect 86539 266388 86605 266389
rect 86539 266324 86540 266388
rect 86604 266324 86605 266388
rect 86539 266323 86605 266324
rect 87459 266388 87525 266389
rect 87459 266324 87460 266388
rect 87524 266324 87525 266388
rect 87459 266323 87525 266324
rect 88747 266388 88813 266389
rect 88747 266324 88748 266388
rect 88812 266324 88813 266388
rect 88747 266323 88813 266324
rect 90035 266388 90101 266389
rect 90035 266324 90036 266388
rect 90100 266324 90101 266388
rect 90035 266323 90101 266324
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 250308 85574 266058
rect 91794 256394 92414 268000
rect 93350 266389 93410 269590
rect 93597 269588 93598 269652
rect 93662 269588 93663 269652
rect 93597 269587 93663 269588
rect 94549 269652 94615 269653
rect 94549 269588 94550 269652
rect 94614 269588 94615 269652
rect 95912 269650 95972 270106
rect 96048 269650 96108 270106
rect 97000 269650 97060 270106
rect 98088 269650 98148 270106
rect 98496 269650 98556 270106
rect 99448 269650 99508 270106
rect 95912 269590 95986 269650
rect 96048 269590 96170 269650
rect 97000 269590 97090 269650
rect 98088 269590 98194 269650
rect 98496 269590 98562 269650
rect 94549 269587 94615 269588
rect 95926 268837 95986 269590
rect 96110 268837 96170 269590
rect 95923 268836 95989 268837
rect 95923 268772 95924 268836
rect 95988 268772 95989 268836
rect 95923 268771 95989 268772
rect 96107 268836 96173 268837
rect 96107 268772 96108 268836
rect 96172 268772 96173 268836
rect 96107 268771 96173 268772
rect 93347 266388 93413 266389
rect 93347 266324 93348 266388
rect 93412 266324 93413 266388
rect 93347 266323 93413 266324
rect 91794 256158 91826 256394
rect 92062 256158 92146 256394
rect 92382 256158 92414 256394
rect 91794 256074 92414 256158
rect 91794 255838 91826 256074
rect 92062 255838 92146 256074
rect 92382 255838 92414 256074
rect 91794 250308 92414 255838
rect 95514 260114 96134 268000
rect 97030 267749 97090 269590
rect 98134 267749 98194 269590
rect 98502 268837 98562 269590
rect 99422 269590 99508 269650
rect 100672 269650 100732 270106
rect 101080 269650 101140 270106
rect 100672 269590 100770 269650
rect 99422 268837 99482 269590
rect 100710 268837 100770 269590
rect 101078 269590 101140 269650
rect 101760 269650 101820 270106
rect 102848 269650 102908 270106
rect 103528 269650 103588 270106
rect 103936 269650 103996 270106
rect 101760 269590 101874 269650
rect 98499 268836 98565 268837
rect 98499 268772 98500 268836
rect 98564 268772 98565 268836
rect 98499 268771 98565 268772
rect 99419 268836 99485 268837
rect 99419 268772 99420 268836
rect 99484 268772 99485 268836
rect 99419 268771 99485 268772
rect 100707 268836 100773 268837
rect 100707 268772 100708 268836
rect 100772 268772 100773 268836
rect 100707 268771 100773 268772
rect 97027 267748 97093 267749
rect 97027 267684 97028 267748
rect 97092 267684 97093 267748
rect 97027 267683 97093 267684
rect 98131 267748 98197 267749
rect 98131 267684 98132 267748
rect 98196 267684 98197 267748
rect 98131 267683 98197 267684
rect 95514 259878 95546 260114
rect 95782 259878 95866 260114
rect 96102 259878 96134 260114
rect 95514 259794 96134 259878
rect 95514 259558 95546 259794
rect 95782 259558 95866 259794
rect 96102 259558 96134 259794
rect 95514 250308 96134 259558
rect 99234 261954 99854 268000
rect 101078 267069 101138 269590
rect 101814 268565 101874 269590
rect 102734 269590 102908 269650
rect 103286 269590 103588 269650
rect 103838 269590 103996 269650
rect 105296 269650 105356 270106
rect 105976 269650 106036 270106
rect 105296 269590 105370 269650
rect 101811 268564 101877 268565
rect 101811 268500 101812 268564
rect 101876 268500 101877 268564
rect 101811 268499 101877 268500
rect 102734 267749 102794 269590
rect 103286 268157 103346 269590
rect 103838 268429 103898 269590
rect 103835 268428 103901 268429
rect 103835 268364 103836 268428
rect 103900 268364 103901 268428
rect 103835 268363 103901 268364
rect 103283 268156 103349 268157
rect 103283 268092 103284 268156
rect 103348 268092 103349 268156
rect 103283 268091 103349 268092
rect 102731 267748 102797 267749
rect 102731 267684 102732 267748
rect 102796 267684 102797 267748
rect 102731 267683 102797 267684
rect 101075 267068 101141 267069
rect 101075 267004 101076 267068
rect 101140 267004 101141 267068
rect 101075 267003 101141 267004
rect 99234 261718 99266 261954
rect 99502 261718 99586 261954
rect 99822 261718 99854 261954
rect 99234 261634 99854 261718
rect 99234 261398 99266 261634
rect 99502 261398 99586 261634
rect 99822 261398 99854 261634
rect 99234 250308 99854 261398
rect 102954 265674 103574 268000
rect 105310 266525 105370 269590
rect 105862 269590 106036 269650
rect 106384 269650 106444 270106
rect 107608 269650 107668 270106
rect 108288 269650 108348 270106
rect 108696 269650 108756 270106
rect 109784 269650 109844 270106
rect 111008 269925 111068 270106
rect 111005 269924 111071 269925
rect 111005 269860 111006 269924
rect 111070 269860 111071 269924
rect 111005 269859 111071 269860
rect 106384 269590 106474 269650
rect 105862 267205 105922 269590
rect 106414 268837 106474 269590
rect 107518 269590 107668 269650
rect 108254 269590 108348 269650
rect 108622 269590 108756 269650
rect 109542 269590 109844 269650
rect 111144 269650 111204 270106
rect 112232 269650 112292 270106
rect 113320 269650 113380 270106
rect 113592 269650 113652 270106
rect 114408 269650 114468 270106
rect 111144 269590 111258 269650
rect 112232 269590 112362 269650
rect 106411 268836 106477 268837
rect 106411 268772 106412 268836
rect 106476 268772 106477 268836
rect 106411 268771 106477 268772
rect 105859 267204 105925 267205
rect 105859 267140 105860 267204
rect 105924 267140 105925 267204
rect 105859 267139 105925 267140
rect 105307 266524 105373 266525
rect 105307 266460 105308 266524
rect 105372 266460 105373 266524
rect 105307 266459 105373 266460
rect 107518 266389 107578 269590
rect 108254 267341 108314 269590
rect 108251 267340 108317 267341
rect 108251 267276 108252 267340
rect 108316 267276 108317 267340
rect 108251 267275 108317 267276
rect 108622 266389 108682 269590
rect 109542 267069 109602 269590
rect 109539 267068 109605 267069
rect 109539 267004 109540 267068
rect 109604 267004 109605 267068
rect 109539 267003 109605 267004
rect 107515 266388 107581 266389
rect 107515 266324 107516 266388
rect 107580 266324 107581 266388
rect 107515 266323 107581 266324
rect 108619 266388 108685 266389
rect 108619 266324 108620 266388
rect 108684 266324 108685 266388
rect 108619 266323 108685 266324
rect 102954 265438 102986 265674
rect 103222 265438 103306 265674
rect 103542 265438 103574 265674
rect 102954 265354 103574 265438
rect 102954 265118 102986 265354
rect 103222 265118 103306 265354
rect 103542 265118 103574 265354
rect 102954 250308 103574 265118
rect 109794 255454 110414 268000
rect 111198 267749 111258 269590
rect 112302 267749 112362 269590
rect 113222 269590 113380 269650
rect 113590 269590 113652 269650
rect 114326 269590 114468 269650
rect 115768 269650 115828 270106
rect 116040 269650 116100 270106
rect 116992 269650 117052 270106
rect 118080 269650 118140 270106
rect 118488 269650 118548 270106
rect 119168 269650 119228 270106
rect 120936 269650 120996 270106
rect 115768 269590 115858 269650
rect 111195 267748 111261 267749
rect 111195 267684 111196 267748
rect 111260 267684 111261 267748
rect 111195 267683 111261 267684
rect 112299 267748 112365 267749
rect 112299 267684 112300 267748
rect 112364 267684 112365 267748
rect 112299 267683 112365 267684
rect 113222 266661 113282 269590
rect 113590 268157 113650 269590
rect 113587 268156 113653 268157
rect 113587 268092 113588 268156
rect 113652 268092 113653 268156
rect 113587 268091 113653 268092
rect 113219 266660 113285 266661
rect 113219 266596 113220 266660
rect 113284 266596 113285 266660
rect 113219 266595 113285 266596
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 250308 110414 254898
rect 113514 259174 114134 268000
rect 114326 266389 114386 269590
rect 115798 269109 115858 269590
rect 115982 269590 116100 269650
rect 116902 269590 117052 269650
rect 118006 269590 118140 269650
rect 118374 269590 118548 269650
rect 119110 269590 119228 269650
rect 120766 269590 120996 269650
rect 123520 269650 123580 270106
rect 125968 269650 126028 270106
rect 123520 269590 123586 269650
rect 115795 269108 115861 269109
rect 115795 269044 115796 269108
rect 115860 269044 115861 269108
rect 115795 269043 115861 269044
rect 115982 267477 116042 269590
rect 116902 268973 116962 269590
rect 116899 268972 116965 268973
rect 116899 268908 116900 268972
rect 116964 268908 116965 268972
rect 116899 268907 116965 268908
rect 115979 267476 116045 267477
rect 115979 267412 115980 267476
rect 116044 267412 116045 267476
rect 115979 267411 116045 267412
rect 114323 266388 114389 266389
rect 114323 266324 114324 266388
rect 114388 266324 114389 266388
rect 114323 266323 114389 266324
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 250308 114134 258618
rect 117234 262894 117854 268000
rect 118006 266661 118066 269590
rect 118374 267477 118434 269590
rect 119110 267749 119170 269590
rect 120766 267749 120826 269590
rect 119107 267748 119173 267749
rect 119107 267684 119108 267748
rect 119172 267684 119173 267748
rect 119107 267683 119173 267684
rect 120763 267748 120829 267749
rect 120763 267684 120764 267748
rect 120828 267684 120829 267748
rect 120763 267683 120829 267684
rect 118371 267476 118437 267477
rect 118371 267412 118372 267476
rect 118436 267412 118437 267476
rect 118371 267411 118437 267412
rect 118003 266660 118069 266661
rect 118003 266596 118004 266660
rect 118068 266596 118069 266660
rect 118003 266595 118069 266596
rect 120954 266614 121574 268000
rect 123526 267613 123586 269590
rect 125918 269590 126028 269650
rect 128280 269650 128340 270106
rect 131000 269650 131060 270106
rect 133448 269789 133508 270106
rect 135896 269789 135956 270106
rect 138480 269789 138540 270106
rect 140928 269789 140988 270106
rect 133445 269788 133511 269789
rect 133445 269724 133446 269788
rect 133510 269724 133511 269788
rect 133445 269723 133511 269724
rect 135893 269788 135959 269789
rect 135893 269724 135894 269788
rect 135958 269724 135959 269788
rect 135893 269723 135959 269724
rect 138477 269788 138543 269789
rect 138477 269724 138478 269788
rect 138542 269724 138543 269788
rect 138477 269723 138543 269724
rect 140925 269788 140991 269789
rect 140925 269724 140926 269788
rect 140990 269724 140991 269788
rect 140925 269723 140991 269724
rect 143512 269653 143572 270106
rect 145960 269653 146020 270106
rect 148544 269925 148604 270106
rect 148541 269924 148607 269925
rect 148541 269860 148542 269924
rect 148606 269860 148607 269924
rect 148541 269859 148607 269860
rect 128280 269590 128370 269650
rect 125918 267749 125978 269590
rect 128310 268157 128370 269590
rect 130886 269590 131060 269650
rect 143509 269652 143575 269653
rect 128307 268156 128373 268157
rect 128307 268092 128308 268156
rect 128372 268092 128373 268156
rect 128307 268091 128373 268092
rect 125915 267748 125981 267749
rect 125915 267684 125916 267748
rect 125980 267684 125981 267748
rect 125915 267683 125981 267684
rect 123523 267612 123589 267613
rect 123523 267548 123524 267612
rect 123588 267548 123589 267612
rect 123523 267547 123589 267548
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 250308 117854 262338
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 250308 121574 266058
rect 127794 256394 128414 268000
rect 130886 267613 130946 269590
rect 143509 269588 143510 269652
rect 143574 269588 143575 269652
rect 143509 269587 143575 269588
rect 145957 269652 146023 269653
rect 145957 269588 145958 269652
rect 146022 269588 146023 269652
rect 150992 269650 151052 270106
rect 145957 269587 146023 269588
rect 150942 269590 151052 269650
rect 153440 269650 153500 270106
rect 155888 269650 155948 270106
rect 158472 269650 158532 270106
rect 160920 269650 160980 270106
rect 153440 269590 154130 269650
rect 155888 269590 155970 269650
rect 158472 269590 158546 269650
rect 130883 267612 130949 267613
rect 130883 267548 130884 267612
rect 130948 267548 130949 267612
rect 130883 267547 130949 267548
rect 127794 256158 127826 256394
rect 128062 256158 128146 256394
rect 128382 256158 128414 256394
rect 127794 256074 128414 256158
rect 127794 255838 127826 256074
rect 128062 255838 128146 256074
rect 128382 255838 128414 256074
rect 127794 250308 128414 255838
rect 131514 260114 132134 268000
rect 131514 259878 131546 260114
rect 131782 259878 131866 260114
rect 132102 259878 132134 260114
rect 131514 259794 132134 259878
rect 131514 259558 131546 259794
rect 131782 259558 131866 259794
rect 132102 259558 132134 259794
rect 131514 250308 132134 259558
rect 135234 261954 135854 268000
rect 135234 261718 135266 261954
rect 135502 261718 135586 261954
rect 135822 261718 135854 261954
rect 135234 261634 135854 261718
rect 135234 261398 135266 261634
rect 135502 261398 135586 261634
rect 135822 261398 135854 261634
rect 135234 250308 135854 261398
rect 138954 265674 139574 268000
rect 138954 265438 138986 265674
rect 139222 265438 139306 265674
rect 139542 265438 139574 265674
rect 138954 265354 139574 265438
rect 138954 265118 138986 265354
rect 139222 265118 139306 265354
rect 139542 265118 139574 265354
rect 138954 250308 139574 265118
rect 145794 255454 146414 268000
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 250308 146414 254898
rect 149514 259174 150134 268000
rect 150942 267749 151002 269590
rect 150939 267748 151005 267749
rect 150939 267684 150940 267748
rect 151004 267684 151005 267748
rect 150939 267683 151005 267684
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 250308 150134 258618
rect 153234 262894 153854 268000
rect 154070 267477 154130 269590
rect 155910 267613 155970 269590
rect 155907 267612 155973 267613
rect 155907 267548 155908 267612
rect 155972 267548 155973 267612
rect 155907 267547 155973 267548
rect 154067 267476 154133 267477
rect 154067 267412 154068 267476
rect 154132 267412 154133 267476
rect 154067 267411 154133 267412
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 250308 153854 262338
rect 156954 266614 157574 268000
rect 158486 267749 158546 269590
rect 160878 269590 160980 269650
rect 163368 269650 163428 270106
rect 165952 269650 166012 270106
rect 183224 269650 183284 270106
rect 163368 269590 163514 269650
rect 158483 267748 158549 267749
rect 158483 267684 158484 267748
rect 158548 267684 158549 267748
rect 158483 267683 158549 267684
rect 160878 267613 160938 269590
rect 163454 267749 163514 269590
rect 165846 269590 166012 269650
rect 183142 269590 183284 269650
rect 183360 269650 183420 270106
rect 183360 269590 183570 269650
rect 163451 267748 163517 267749
rect 163451 267684 163452 267748
rect 163516 267684 163517 267748
rect 163451 267683 163517 267684
rect 160875 267612 160941 267613
rect 160875 267548 160876 267612
rect 160940 267548 160941 267612
rect 160875 267547 160941 267548
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 250308 157574 266058
rect 163794 256394 164414 268000
rect 165846 266933 165906 269590
rect 165843 266932 165909 266933
rect 165843 266868 165844 266932
rect 165908 266868 165909 266932
rect 165843 266867 165909 266868
rect 163794 256158 163826 256394
rect 164062 256158 164146 256394
rect 164382 256158 164414 256394
rect 163794 256074 164414 256158
rect 163794 255838 163826 256074
rect 164062 255838 164146 256074
rect 164382 255838 164414 256074
rect 163794 250308 164414 255838
rect 167514 260114 168134 268000
rect 167514 259878 167546 260114
rect 167782 259878 167866 260114
rect 168102 259878 168134 260114
rect 167514 259794 168134 259878
rect 167514 259558 167546 259794
rect 167782 259558 167866 259794
rect 168102 259558 168134 259794
rect 167514 250308 168134 259558
rect 171234 261954 171854 268000
rect 171234 261718 171266 261954
rect 171502 261718 171586 261954
rect 171822 261718 171854 261954
rect 171234 261634 171854 261718
rect 171234 261398 171266 261634
rect 171502 261398 171586 261634
rect 171822 261398 171854 261634
rect 171234 250308 171854 261398
rect 174954 265674 175574 268000
rect 174954 265438 174986 265674
rect 175222 265438 175306 265674
rect 175542 265438 175574 265674
rect 174954 265354 175574 265438
rect 174954 265118 174986 265354
rect 175222 265118 175306 265354
rect 175542 265118 175574 265354
rect 174954 250308 175574 265118
rect 181794 255454 182414 268000
rect 183142 267341 183202 269590
rect 183139 267340 183205 267341
rect 183139 267276 183140 267340
rect 183204 267276 183205 267340
rect 183139 267275 183205 267276
rect 183510 267069 183570 269590
rect 183507 267068 183573 267069
rect 183507 267004 183508 267068
rect 183572 267004 183573 267068
rect 183507 267003 183573 267004
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 250308 182414 254898
rect 185514 259174 186134 268000
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 250308 186134 258618
rect 189234 262894 189854 268000
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 250308 189854 262338
rect 192954 266614 193574 268000
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 250308 193574 266058
rect 178539 249932 178605 249933
rect 178539 249868 178540 249932
rect 178604 249868 178605 249932
rect 178539 249867 178605 249868
rect 179643 249932 179709 249933
rect 179643 249868 179644 249932
rect 179708 249868 179709 249932
rect 179643 249867 179709 249868
rect 190867 249932 190933 249933
rect 190867 249868 190868 249932
rect 190932 249868 190933 249932
rect 190867 249867 190933 249868
rect 178542 248430 178602 249867
rect 59862 248370 60290 248430
rect 178464 248370 178602 248430
rect 179646 248430 179706 249867
rect 190870 248430 190930 249867
rect 179646 248370 179748 248430
rect 59862 164930 59922 248370
rect 178464 248202 178524 248370
rect 179688 248202 179748 248370
rect 190840 248370 190930 248430
rect 190840 248202 190900 248370
rect 60272 237454 60620 237486
rect 60272 237218 60328 237454
rect 60564 237218 60620 237454
rect 60272 237134 60620 237218
rect 60272 236898 60328 237134
rect 60564 236898 60620 237134
rect 60272 236866 60620 236898
rect 196000 237454 196348 237486
rect 196000 237218 196056 237454
rect 196292 237218 196348 237454
rect 196000 237134 196348 237218
rect 196000 236898 196056 237134
rect 196292 236898 196348 237134
rect 196000 236866 196348 236898
rect 60952 219454 61300 219486
rect 60952 219218 61008 219454
rect 61244 219218 61300 219454
rect 60952 219134 61300 219218
rect 60952 218898 61008 219134
rect 61244 218898 61300 219134
rect 60952 218866 61300 218898
rect 195320 219454 195668 219486
rect 195320 219218 195376 219454
rect 195612 219218 195668 219454
rect 195320 219134 195668 219218
rect 195320 218898 195376 219134
rect 195612 218898 195668 219134
rect 195320 218866 195668 218898
rect 60272 201454 60620 201486
rect 60272 201218 60328 201454
rect 60564 201218 60620 201454
rect 60272 201134 60620 201218
rect 60272 200898 60328 201134
rect 60564 200898 60620 201134
rect 60272 200866 60620 200898
rect 196000 201454 196348 201486
rect 196000 201218 196056 201454
rect 196292 201218 196348 201454
rect 196000 201134 196348 201218
rect 196000 200898 196056 201134
rect 196292 200898 196348 201134
rect 196000 200866 196348 200898
rect 60952 183454 61300 183486
rect 60952 183218 61008 183454
rect 61244 183218 61300 183454
rect 60952 183134 61300 183218
rect 60952 182898 61008 183134
rect 61244 182898 61300 183134
rect 60952 182866 61300 182898
rect 195320 183454 195668 183486
rect 195320 183218 195376 183454
rect 195612 183218 195668 183454
rect 195320 183134 195668 183218
rect 195320 182898 195376 183134
rect 195612 182898 195668 183134
rect 195320 182866 195668 182898
rect 76056 164930 76116 165106
rect 59862 164870 60290 164930
rect 59514 152114 60134 163000
rect 59514 151878 59546 152114
rect 59782 151878 59866 152114
rect 60102 151878 60134 152114
rect 59514 151794 60134 151878
rect 59514 151558 59546 151794
rect 59782 151558 59866 151794
rect 60102 151558 60134 151794
rect 59514 145308 60134 151558
rect 60230 145210 60290 164870
rect 76054 164870 76116 164930
rect 77144 164930 77204 165106
rect 78232 164930 78292 165106
rect 79592 164930 79652 165106
rect 80544 164930 80604 165106
rect 77144 164870 77218 164930
rect 78232 164870 78322 164930
rect 63234 153954 63854 163000
rect 63234 153718 63266 153954
rect 63502 153718 63586 153954
rect 63822 153718 63854 153954
rect 63234 153634 63854 153718
rect 63234 153398 63266 153634
rect 63502 153398 63586 153634
rect 63822 153398 63854 153634
rect 63234 145308 63854 153398
rect 66954 157674 67574 163000
rect 66954 157438 66986 157674
rect 67222 157438 67306 157674
rect 67542 157438 67574 157674
rect 66954 157354 67574 157438
rect 66954 157118 66986 157354
rect 67222 157118 67306 157354
rect 67542 157118 67574 157354
rect 66954 145308 67574 157118
rect 73794 147454 74414 163000
rect 76054 162757 76114 164870
rect 76051 162756 76117 162757
rect 76051 162692 76052 162756
rect 76116 162692 76117 162756
rect 76051 162691 76117 162692
rect 77158 162213 77218 164870
rect 77155 162212 77221 162213
rect 77155 162148 77156 162212
rect 77220 162148 77221 162212
rect 77155 162147 77221 162148
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 145308 74414 146898
rect 77514 151174 78134 163000
rect 78262 162757 78322 164870
rect 79550 164870 79652 164930
rect 80470 164870 80604 164930
rect 81768 164930 81828 165106
rect 83128 164930 83188 165106
rect 81768 164870 82002 164930
rect 79550 162757 79610 164870
rect 80470 162757 80530 164870
rect 78259 162756 78325 162757
rect 78259 162692 78260 162756
rect 78324 162692 78325 162756
rect 78259 162691 78325 162692
rect 79547 162756 79613 162757
rect 79547 162692 79548 162756
rect 79612 162692 79613 162756
rect 79547 162691 79613 162692
rect 80467 162756 80533 162757
rect 80467 162692 80468 162756
rect 80532 162692 80533 162756
rect 80467 162691 80533 162692
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 145308 78134 150618
rect 81234 154894 81854 163000
rect 81942 162757 82002 164870
rect 83046 164870 83188 164930
rect 84216 164930 84276 165106
rect 84216 164870 84394 164930
rect 83046 162757 83106 164870
rect 84334 162757 84394 164870
rect 85440 164661 85500 165106
rect 86528 164930 86588 165106
rect 87616 164930 87676 165106
rect 88296 164930 88356 165106
rect 88704 164930 88764 165106
rect 90064 164930 90124 165106
rect 86528 164870 86602 164930
rect 87616 164870 87706 164930
rect 88296 164870 88442 164930
rect 88704 164870 88810 164930
rect 85437 164660 85503 164661
rect 85437 164596 85438 164660
rect 85502 164596 85503 164660
rect 85437 164595 85503 164596
rect 81939 162756 82005 162757
rect 81939 162692 81940 162756
rect 82004 162692 82005 162756
rect 81939 162691 82005 162692
rect 83043 162756 83109 162757
rect 83043 162692 83044 162756
rect 83108 162692 83109 162756
rect 83043 162691 83109 162692
rect 84331 162756 84397 162757
rect 84331 162692 84332 162756
rect 84396 162692 84397 162756
rect 84331 162691 84397 162692
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 145308 81854 154338
rect 84954 158614 85574 163000
rect 86542 162757 86602 164870
rect 87646 162757 87706 164870
rect 86539 162756 86605 162757
rect 86539 162692 86540 162756
rect 86604 162692 86605 162756
rect 86539 162691 86605 162692
rect 87643 162756 87709 162757
rect 87643 162692 87644 162756
rect 87708 162692 87709 162756
rect 87643 162691 87709 162692
rect 88382 162213 88442 164870
rect 88750 162757 88810 164870
rect 90038 164870 90124 164930
rect 90744 164930 90804 165106
rect 91288 164930 91348 165106
rect 92376 164930 92436 165106
rect 93464 164930 93524 165106
rect 90744 164870 90834 164930
rect 91288 164870 91386 164930
rect 90038 162757 90098 164870
rect 90774 162757 90834 164870
rect 91326 162757 91386 164870
rect 91510 164870 92436 164930
rect 93350 164870 93524 164930
rect 93600 164930 93660 165106
rect 94552 164930 94612 165106
rect 93600 164870 93778 164930
rect 88747 162756 88813 162757
rect 88747 162692 88748 162756
rect 88812 162692 88813 162756
rect 88747 162691 88813 162692
rect 90035 162756 90101 162757
rect 90035 162692 90036 162756
rect 90100 162692 90101 162756
rect 90035 162691 90101 162692
rect 90771 162756 90837 162757
rect 90771 162692 90772 162756
rect 90836 162692 90837 162756
rect 90771 162691 90837 162692
rect 91323 162756 91389 162757
rect 91323 162692 91324 162756
rect 91388 162692 91389 162756
rect 91323 162691 91389 162692
rect 91510 162485 91570 164870
rect 91507 162484 91573 162485
rect 91507 162420 91508 162484
rect 91572 162420 91573 162484
rect 91507 162419 91573 162420
rect 88379 162212 88445 162213
rect 88379 162148 88380 162212
rect 88444 162148 88445 162212
rect 88379 162147 88445 162148
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 145308 85574 158058
rect 91794 148394 92414 163000
rect 93350 162757 93410 164870
rect 93347 162756 93413 162757
rect 93347 162692 93348 162756
rect 93412 162692 93413 162756
rect 93347 162691 93413 162692
rect 93718 162213 93778 164870
rect 94454 164870 94612 164930
rect 95912 164930 95972 165106
rect 96048 164933 96108 165106
rect 96048 164932 96173 164933
rect 95912 164870 95986 164930
rect 96048 164870 96108 164932
rect 94454 162757 94514 164870
rect 95926 163165 95986 164870
rect 96107 164868 96108 164870
rect 96172 164868 96173 164932
rect 97000 164930 97060 165106
rect 98088 164930 98148 165106
rect 98496 164930 98556 165106
rect 99448 164930 99508 165106
rect 97000 164870 97090 164930
rect 98088 164870 98194 164930
rect 98496 164870 98562 164930
rect 96107 164867 96173 164868
rect 95923 163164 95989 163165
rect 95923 163100 95924 163164
rect 95988 163100 95989 163164
rect 95923 163099 95989 163100
rect 94451 162756 94517 162757
rect 94451 162692 94452 162756
rect 94516 162692 94517 162756
rect 94451 162691 94517 162692
rect 93715 162212 93781 162213
rect 93715 162148 93716 162212
rect 93780 162148 93781 162212
rect 93715 162147 93781 162148
rect 91794 148158 91826 148394
rect 92062 148158 92146 148394
rect 92382 148158 92414 148394
rect 91794 148074 92414 148158
rect 91794 147838 91826 148074
rect 92062 147838 92146 148074
rect 92382 147838 92414 148074
rect 91794 145308 92414 147838
rect 95514 152114 96134 163000
rect 97030 162757 97090 164870
rect 98134 162757 98194 164870
rect 98502 164253 98562 164870
rect 99422 164870 99508 164930
rect 100672 164930 100732 165106
rect 101080 164930 101140 165106
rect 100672 164870 100770 164930
rect 98499 164252 98565 164253
rect 98499 164188 98500 164252
rect 98564 164188 98565 164252
rect 98499 164187 98565 164188
rect 99422 163165 99482 164870
rect 99419 163164 99485 163165
rect 99419 163100 99420 163164
rect 99484 163100 99485 163164
rect 99419 163099 99485 163100
rect 97027 162756 97093 162757
rect 97027 162692 97028 162756
rect 97092 162692 97093 162756
rect 97027 162691 97093 162692
rect 98131 162756 98197 162757
rect 98131 162692 98132 162756
rect 98196 162692 98197 162756
rect 98131 162691 98197 162692
rect 95514 151878 95546 152114
rect 95782 151878 95866 152114
rect 96102 151878 96134 152114
rect 95514 151794 96134 151878
rect 95514 151558 95546 151794
rect 95782 151558 95866 151794
rect 96102 151558 96134 151794
rect 95514 145308 96134 151558
rect 99234 153954 99854 163000
rect 100710 162757 100770 164870
rect 101078 164870 101140 164930
rect 101760 164930 101820 165106
rect 102848 164930 102908 165106
rect 101760 164870 101874 164930
rect 101078 164253 101138 164870
rect 101075 164252 101141 164253
rect 101075 164188 101076 164252
rect 101140 164188 101141 164252
rect 101075 164187 101141 164188
rect 100707 162756 100773 162757
rect 100707 162692 100708 162756
rect 100772 162692 100773 162756
rect 100707 162691 100773 162692
rect 101814 162077 101874 164870
rect 102734 164870 102908 164930
rect 102734 162757 102794 164870
rect 103528 164661 103588 165106
rect 103936 164930 103996 165106
rect 103838 164870 103996 164930
rect 105296 164930 105356 165106
rect 105296 164870 105370 164930
rect 103525 164660 103591 164661
rect 103525 164596 103526 164660
rect 103590 164596 103591 164660
rect 103525 164595 103591 164596
rect 102731 162756 102797 162757
rect 102731 162692 102732 162756
rect 102796 162692 102797 162756
rect 102731 162691 102797 162692
rect 101811 162076 101877 162077
rect 101811 162012 101812 162076
rect 101876 162012 101877 162076
rect 101811 162011 101877 162012
rect 99234 153718 99266 153954
rect 99502 153718 99586 153954
rect 99822 153718 99854 153954
rect 99234 153634 99854 153718
rect 99234 153398 99266 153634
rect 99502 153398 99586 153634
rect 99822 153398 99854 153634
rect 99234 145308 99854 153398
rect 102954 157674 103574 163000
rect 103838 162757 103898 164870
rect 105310 162757 105370 164870
rect 105976 164661 106036 165106
rect 106384 164930 106444 165106
rect 107608 164930 107668 165106
rect 108288 164930 108348 165106
rect 108696 164930 108756 165106
rect 109784 164930 109844 165106
rect 106384 164870 106474 164930
rect 105973 164660 106039 164661
rect 105973 164596 105974 164660
rect 106038 164596 106039 164660
rect 105973 164595 106039 164596
rect 106414 162757 106474 164870
rect 107518 164870 107668 164930
rect 108254 164870 108348 164930
rect 108622 164870 108756 164930
rect 109542 164870 109844 164930
rect 111008 164930 111068 165106
rect 111144 164930 111204 165106
rect 112232 164930 112292 165106
rect 113320 164930 113380 165106
rect 113592 164930 113652 165106
rect 111008 164870 111074 164930
rect 111144 164870 111258 164930
rect 112232 164870 112362 164930
rect 113320 164870 113466 164930
rect 103835 162756 103901 162757
rect 103835 162692 103836 162756
rect 103900 162692 103901 162756
rect 103835 162691 103901 162692
rect 105307 162756 105373 162757
rect 105307 162692 105308 162756
rect 105372 162692 105373 162756
rect 105307 162691 105373 162692
rect 106411 162756 106477 162757
rect 106411 162692 106412 162756
rect 106476 162692 106477 162756
rect 106411 162691 106477 162692
rect 107518 162485 107578 164870
rect 108254 164253 108314 164870
rect 108251 164252 108317 164253
rect 108251 164188 108252 164252
rect 108316 164188 108317 164252
rect 108251 164187 108317 164188
rect 108622 162757 108682 164870
rect 109542 162757 109602 164870
rect 108619 162756 108685 162757
rect 108619 162692 108620 162756
rect 108684 162692 108685 162756
rect 108619 162691 108685 162692
rect 109539 162756 109605 162757
rect 109539 162692 109540 162756
rect 109604 162692 109605 162756
rect 109539 162691 109605 162692
rect 107515 162484 107581 162485
rect 107515 162420 107516 162484
rect 107580 162420 107581 162484
rect 107515 162419 107581 162420
rect 102954 157438 102986 157674
rect 103222 157438 103306 157674
rect 103542 157438 103574 157674
rect 102954 157354 103574 157438
rect 102954 157118 102986 157354
rect 103222 157118 103306 157354
rect 103542 157118 103574 157354
rect 102954 145308 103574 157118
rect 109794 147454 110414 163000
rect 111014 162757 111074 164870
rect 111198 163981 111258 164870
rect 111195 163980 111261 163981
rect 111195 163916 111196 163980
rect 111260 163916 111261 163980
rect 111195 163915 111261 163916
rect 111011 162756 111077 162757
rect 111011 162692 111012 162756
rect 111076 162692 111077 162756
rect 111011 162691 111077 162692
rect 112302 162213 112362 164870
rect 113406 163709 113466 164870
rect 113590 164870 113652 164930
rect 113403 163708 113469 163709
rect 113403 163644 113404 163708
rect 113468 163644 113469 163708
rect 113403 163643 113469 163644
rect 113590 163570 113650 164870
rect 114408 164661 114468 165106
rect 115768 164933 115828 165106
rect 115765 164932 115831 164933
rect 115765 164868 115766 164932
rect 115830 164868 115831 164932
rect 116040 164930 116100 165106
rect 116992 164930 117052 165106
rect 115765 164867 115831 164868
rect 115982 164870 116100 164930
rect 116902 164870 117052 164930
rect 114405 164660 114471 164661
rect 114405 164596 114406 164660
rect 114470 164596 114471 164660
rect 114405 164595 114471 164596
rect 113222 163510 113650 163570
rect 113222 162757 113282 163510
rect 113219 162756 113285 162757
rect 113219 162692 113220 162756
rect 113284 162692 113285 162756
rect 113219 162691 113285 162692
rect 112299 162212 112365 162213
rect 112299 162148 112300 162212
rect 112364 162148 112365 162212
rect 112299 162147 112365 162148
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 145308 110414 146898
rect 113514 151174 114134 163000
rect 115982 162485 116042 164870
rect 116902 162757 116962 164870
rect 118080 164661 118140 165106
rect 118488 164930 118548 165106
rect 119168 164930 119228 165106
rect 120936 164930 120996 165106
rect 118374 164870 118548 164930
rect 119110 164870 119228 164930
rect 120766 164870 120996 164930
rect 123520 164930 123580 165106
rect 125968 164930 126028 165106
rect 123520 164870 123586 164930
rect 118077 164660 118143 164661
rect 118077 164596 118078 164660
rect 118142 164596 118143 164660
rect 118077 164595 118143 164596
rect 116899 162756 116965 162757
rect 116899 162692 116900 162756
rect 116964 162692 116965 162756
rect 116899 162691 116965 162692
rect 115979 162484 116045 162485
rect 115979 162420 115980 162484
rect 116044 162420 116045 162484
rect 115979 162419 116045 162420
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 145308 114134 150618
rect 117234 154894 117854 163000
rect 118374 162757 118434 164870
rect 119110 162757 119170 164870
rect 120766 162757 120826 164870
rect 123526 164253 123586 164870
rect 125918 164870 126028 164930
rect 128280 164930 128340 165106
rect 131000 164930 131060 165106
rect 128280 164870 128370 164930
rect 123523 164252 123589 164253
rect 123523 164188 123524 164252
rect 123588 164188 123589 164252
rect 123523 164187 123589 164188
rect 118371 162756 118437 162757
rect 118371 162692 118372 162756
rect 118436 162692 118437 162756
rect 118371 162691 118437 162692
rect 119107 162756 119173 162757
rect 119107 162692 119108 162756
rect 119172 162692 119173 162756
rect 119107 162691 119173 162692
rect 120763 162756 120829 162757
rect 120763 162692 120764 162756
rect 120828 162692 120829 162756
rect 120763 162691 120829 162692
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 145308 117854 154338
rect 120954 158614 121574 163000
rect 125918 162757 125978 164870
rect 128310 163165 128370 164870
rect 130886 164870 131060 164930
rect 133448 164930 133508 165106
rect 135896 164930 135956 165106
rect 133448 164870 133522 164930
rect 135896 164870 136098 164930
rect 128307 163164 128373 163165
rect 128307 163100 128308 163164
rect 128372 163100 128373 163164
rect 128307 163099 128373 163100
rect 125915 162756 125981 162757
rect 125915 162692 125916 162756
rect 125980 162692 125981 162756
rect 125915 162691 125981 162692
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 145308 121574 158058
rect 127794 148394 128414 163000
rect 130886 162757 130946 164870
rect 130883 162756 130949 162757
rect 130883 162692 130884 162756
rect 130948 162692 130949 162756
rect 130883 162691 130949 162692
rect 127794 148158 127826 148394
rect 128062 148158 128146 148394
rect 128382 148158 128414 148394
rect 127794 148074 128414 148158
rect 127794 147838 127826 148074
rect 128062 147838 128146 148074
rect 128382 147838 128414 148074
rect 127794 145308 128414 147838
rect 131514 152114 132134 163000
rect 133462 162757 133522 164870
rect 133459 162756 133525 162757
rect 133459 162692 133460 162756
rect 133524 162692 133525 162756
rect 133459 162691 133525 162692
rect 131514 151878 131546 152114
rect 131782 151878 131866 152114
rect 132102 151878 132134 152114
rect 131514 151794 132134 151878
rect 131514 151558 131546 151794
rect 131782 151558 131866 151794
rect 132102 151558 132134 151794
rect 131514 145308 132134 151558
rect 135234 153954 135854 163000
rect 136038 162757 136098 164870
rect 138480 164797 138540 165106
rect 140928 164797 140988 165106
rect 143512 164797 143572 165106
rect 145960 164930 146020 165106
rect 148544 164930 148604 165106
rect 150992 164930 151052 165106
rect 145960 164870 146034 164930
rect 148544 164870 148610 164930
rect 138477 164796 138543 164797
rect 138477 164732 138478 164796
rect 138542 164732 138543 164796
rect 138477 164731 138543 164732
rect 140925 164796 140991 164797
rect 140925 164732 140926 164796
rect 140990 164732 140991 164796
rect 140925 164731 140991 164732
rect 143509 164796 143575 164797
rect 143509 164732 143510 164796
rect 143574 164732 143575 164796
rect 143509 164731 143575 164732
rect 145974 164253 146034 164870
rect 148550 164253 148610 164870
rect 150942 164870 151052 164930
rect 150942 164253 151002 164870
rect 153440 164661 153500 165106
rect 155888 164930 155948 165106
rect 158472 164930 158532 165106
rect 160920 164930 160980 165106
rect 155888 164870 155970 164930
rect 158472 164870 158546 164930
rect 153437 164660 153503 164661
rect 153437 164596 153438 164660
rect 153502 164596 153503 164660
rect 153437 164595 153503 164596
rect 145971 164252 146037 164253
rect 145971 164188 145972 164252
rect 146036 164188 146037 164252
rect 145971 164187 146037 164188
rect 148547 164252 148613 164253
rect 148547 164188 148548 164252
rect 148612 164188 148613 164252
rect 148547 164187 148613 164188
rect 150939 164252 151005 164253
rect 150939 164188 150940 164252
rect 151004 164188 151005 164252
rect 150939 164187 151005 164188
rect 136035 162756 136101 162757
rect 136035 162692 136036 162756
rect 136100 162692 136101 162756
rect 136035 162691 136101 162692
rect 135234 153718 135266 153954
rect 135502 153718 135586 153954
rect 135822 153718 135854 153954
rect 135234 153634 135854 153718
rect 135234 153398 135266 153634
rect 135502 153398 135586 153634
rect 135822 153398 135854 153634
rect 135234 145308 135854 153398
rect 138954 157674 139574 163000
rect 138954 157438 138986 157674
rect 139222 157438 139306 157674
rect 139542 157438 139574 157674
rect 138954 157354 139574 157438
rect 138954 157118 138986 157354
rect 139222 157118 139306 157354
rect 139542 157118 139574 157354
rect 138954 145308 139574 157118
rect 145794 147454 146414 163000
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 145308 146414 146898
rect 149514 151174 150134 163000
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 145308 150134 150618
rect 153234 154894 153854 163000
rect 155910 162757 155970 164870
rect 155907 162756 155973 162757
rect 155907 162692 155908 162756
rect 155972 162692 155973 162756
rect 155907 162691 155973 162692
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 145308 153854 154338
rect 156954 158614 157574 163000
rect 158486 162621 158546 164870
rect 160878 164870 160980 164930
rect 158483 162620 158549 162621
rect 158483 162556 158484 162620
rect 158548 162556 158549 162620
rect 158483 162555 158549 162556
rect 160878 162349 160938 164870
rect 163368 164797 163428 165106
rect 163365 164796 163431 164797
rect 163365 164732 163366 164796
rect 163430 164732 163431 164796
rect 163365 164731 163431 164732
rect 165952 164661 166012 165106
rect 183224 164930 183284 165106
rect 183142 164870 183284 164930
rect 183360 164930 183420 165106
rect 183360 164870 183570 164930
rect 165949 164660 166015 164661
rect 165949 164596 165950 164660
rect 166014 164596 166015 164660
rect 165949 164595 166015 164596
rect 160875 162348 160941 162349
rect 160875 162284 160876 162348
rect 160940 162284 160941 162348
rect 160875 162283 160941 162284
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 145308 157574 158058
rect 163794 148394 164414 163000
rect 163794 148158 163826 148394
rect 164062 148158 164146 148394
rect 164382 148158 164414 148394
rect 163794 148074 164414 148158
rect 163794 147838 163826 148074
rect 164062 147838 164146 148074
rect 164382 147838 164414 148074
rect 163794 145308 164414 147838
rect 167514 152114 168134 163000
rect 167514 151878 167546 152114
rect 167782 151878 167866 152114
rect 168102 151878 168134 152114
rect 167514 151794 168134 151878
rect 167514 151558 167546 151794
rect 167782 151558 167866 151794
rect 168102 151558 168134 151794
rect 167514 145308 168134 151558
rect 171234 153954 171854 163000
rect 171234 153718 171266 153954
rect 171502 153718 171586 153954
rect 171822 153718 171854 153954
rect 171234 153634 171854 153718
rect 171234 153398 171266 153634
rect 171502 153398 171586 153634
rect 171822 153398 171854 153634
rect 171234 145308 171854 153398
rect 174954 157674 175574 163000
rect 174954 157438 174986 157674
rect 175222 157438 175306 157674
rect 175542 157438 175574 157674
rect 174954 157354 175574 157438
rect 174954 157118 174986 157354
rect 175222 157118 175306 157354
rect 175542 157118 175574 157354
rect 174954 145308 175574 157118
rect 181794 147454 182414 163000
rect 183142 162621 183202 164870
rect 183510 162757 183570 164870
rect 196574 163845 196634 478619
rect 198043 478548 198109 478549
rect 198043 478484 198044 478548
rect 198108 478484 198109 478548
rect 198043 478483 198109 478484
rect 197859 478276 197925 478277
rect 197859 478212 197860 478276
rect 197924 478212 197925 478276
rect 197859 478211 197925 478212
rect 196755 478004 196821 478005
rect 196755 477940 196756 478004
rect 196820 477940 196821 478004
rect 196755 477939 196821 477940
rect 196758 269109 196818 477939
rect 196755 269108 196821 269109
rect 196755 269044 196756 269108
rect 196820 269044 196821 269108
rect 196755 269043 196821 269044
rect 196571 163844 196637 163845
rect 196571 163780 196572 163844
rect 196636 163780 196637 163844
rect 196571 163779 196637 163780
rect 183507 162756 183573 162757
rect 183507 162692 183508 162756
rect 183572 162692 183573 162756
rect 183507 162691 183573 162692
rect 183139 162620 183205 162621
rect 183139 162556 183140 162620
rect 183204 162556 183205 162620
rect 183139 162555 183205 162556
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 145308 182414 146898
rect 185514 151174 186134 163000
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 145308 186134 150618
rect 189234 154894 189854 163000
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 145308 189854 154338
rect 192954 158614 193574 163000
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 190867 145484 190933 145485
rect 190867 145420 190868 145484
rect 190932 145420 190933 145484
rect 190867 145419 190933 145420
rect 59862 145150 60290 145210
rect 59862 59530 59922 145150
rect 178539 144940 178605 144941
rect 178539 144876 178540 144940
rect 178604 144876 178605 144940
rect 178539 144875 178605 144876
rect 179643 144940 179709 144941
rect 179643 144876 179644 144940
rect 179708 144876 179709 144940
rect 179643 144875 179709 144876
rect 178542 143850 178602 144875
rect 178464 143790 178602 143850
rect 179646 143850 179706 144875
rect 190870 143850 190930 145419
rect 192954 145308 193574 158058
rect 179646 143790 179748 143850
rect 178464 143202 178524 143790
rect 179688 143202 179748 143790
rect 190840 143790 190930 143850
rect 190840 143202 190900 143790
rect 60272 129454 60620 129486
rect 60272 129218 60328 129454
rect 60564 129218 60620 129454
rect 60272 129134 60620 129218
rect 60272 128898 60328 129134
rect 60564 128898 60620 129134
rect 60272 128866 60620 128898
rect 196000 129454 196348 129486
rect 196000 129218 196056 129454
rect 196292 129218 196348 129454
rect 196000 129134 196348 129218
rect 196000 128898 196056 129134
rect 196292 128898 196348 129134
rect 196000 128866 196348 128898
rect 60952 111454 61300 111486
rect 60952 111218 61008 111454
rect 61244 111218 61300 111454
rect 60952 111134 61300 111218
rect 60952 110898 61008 111134
rect 61244 110898 61300 111134
rect 60952 110866 61300 110898
rect 195320 111454 195668 111486
rect 195320 111218 195376 111454
rect 195612 111218 195668 111454
rect 195320 111134 195668 111218
rect 195320 110898 195376 111134
rect 195612 110898 195668 111134
rect 195320 110866 195668 110898
rect 60272 93454 60620 93486
rect 60272 93218 60328 93454
rect 60564 93218 60620 93454
rect 60272 93134 60620 93218
rect 60272 92898 60328 93134
rect 60564 92898 60620 93134
rect 60272 92866 60620 92898
rect 196000 93454 196348 93486
rect 196000 93218 196056 93454
rect 196292 93218 196348 93454
rect 196000 93134 196348 93218
rect 196000 92898 196056 93134
rect 196292 92898 196348 93134
rect 196000 92866 196348 92898
rect 60952 75454 61300 75486
rect 60952 75218 61008 75454
rect 61244 75218 61300 75454
rect 60952 75134 61300 75218
rect 60952 74898 61008 75134
rect 61244 74898 61300 75134
rect 60952 74866 61300 74898
rect 195320 75454 195668 75486
rect 195320 75218 195376 75454
rect 195612 75218 195668 75454
rect 195320 75134 195668 75218
rect 195320 74898 195376 75134
rect 195612 74898 195668 75134
rect 195320 74866 195668 74898
rect 76056 59530 76116 60106
rect 77144 59805 77204 60106
rect 77141 59804 77207 59805
rect 77141 59740 77142 59804
rect 77206 59740 77207 59804
rect 77141 59739 77207 59740
rect 59862 59470 60290 59530
rect 59307 58716 59373 58717
rect 59307 58652 59308 58716
rect 59372 58652 59373 58716
rect 59307 58651 59373 58652
rect 59123 57220 59189 57221
rect 59123 57156 59124 57220
rect 59188 57156 59189 57220
rect 59123 57155 59189 57156
rect 58571 57084 58637 57085
rect 58571 57020 58572 57084
rect 58636 57020 58637 57084
rect 58571 57019 58637 57020
rect 57835 54636 57901 54637
rect 57835 54572 57836 54636
rect 57900 54572 57901 54636
rect 57835 54571 57901 54572
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 25174 60134 58000
rect 60230 57765 60290 59470
rect 76054 59470 76116 59530
rect 78232 59530 78292 60106
rect 79592 59530 79652 60106
rect 80544 59530 80604 60106
rect 78232 59470 78322 59530
rect 60227 57764 60293 57765
rect 60227 57700 60228 57764
rect 60292 57700 60293 57764
rect 60227 57699 60293 57700
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 28894 63854 58000
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 32614 67574 58000
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 39454 74414 58000
rect 76054 57901 76114 59470
rect 76051 57900 76117 57901
rect 76051 57836 76052 57900
rect 76116 57836 76117 57900
rect 76051 57835 76117 57836
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 43174 78134 58000
rect 78262 57901 78322 59470
rect 79550 59470 79652 59530
rect 80470 59470 80604 59530
rect 81768 59530 81828 60106
rect 83128 59805 83188 60106
rect 83125 59804 83191 59805
rect 83125 59740 83126 59804
rect 83190 59740 83191 59804
rect 83125 59739 83191 59740
rect 84216 59530 84276 60106
rect 85440 59530 85500 60106
rect 81768 59470 82002 59530
rect 79550 57901 79610 59470
rect 80470 57901 80530 59470
rect 78259 57900 78325 57901
rect 78259 57836 78260 57900
rect 78324 57836 78325 57900
rect 78259 57835 78325 57836
rect 79547 57900 79613 57901
rect 79547 57836 79548 57900
rect 79612 57836 79613 57900
rect 79547 57835 79613 57836
rect 80467 57900 80533 57901
rect 80467 57836 80468 57900
rect 80532 57836 80533 57900
rect 80467 57835 80533 57836
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 46894 81854 58000
rect 81942 57901 82002 59470
rect 83966 59470 84276 59530
rect 85438 59470 85500 59530
rect 86528 59530 86588 60106
rect 87616 59530 87676 60106
rect 88296 59530 88356 60106
rect 88704 59530 88764 60106
rect 90064 59530 90124 60106
rect 86528 59470 86602 59530
rect 87616 59470 87706 59530
rect 88296 59470 88442 59530
rect 88704 59470 88810 59530
rect 83966 58037 84026 59470
rect 85438 58173 85498 59470
rect 85435 58172 85501 58173
rect 85435 58108 85436 58172
rect 85500 58108 85501 58172
rect 85435 58107 85501 58108
rect 83963 58036 84029 58037
rect 83963 57972 83964 58036
rect 84028 57972 84029 58036
rect 83963 57971 84029 57972
rect 81939 57900 82005 57901
rect 81939 57836 81940 57900
rect 82004 57836 82005 57900
rect 81939 57835 82005 57836
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 50614 85574 58000
rect 86542 57901 86602 59470
rect 87646 57901 87706 59470
rect 88382 57901 88442 59470
rect 88750 57901 88810 59470
rect 90038 59470 90124 59530
rect 90744 59530 90804 60106
rect 91288 59530 91348 60106
rect 92376 59530 92436 60106
rect 93464 59530 93524 60106
rect 90744 59470 90834 59530
rect 91288 59470 91386 59530
rect 90038 57901 90098 59470
rect 90774 57901 90834 59470
rect 91326 57901 91386 59470
rect 92246 59470 92436 59530
rect 93350 59470 93524 59530
rect 93600 59530 93660 60106
rect 94552 59669 94612 60106
rect 94549 59668 94615 59669
rect 94549 59604 94550 59668
rect 94614 59604 94615 59668
rect 95912 59666 95972 60106
rect 95912 59606 95986 59666
rect 94549 59603 94615 59604
rect 93600 59470 93778 59530
rect 92246 58173 92306 59470
rect 92243 58172 92309 58173
rect 92243 58108 92244 58172
rect 92308 58108 92309 58172
rect 92243 58107 92309 58108
rect 86539 57900 86605 57901
rect 86539 57836 86540 57900
rect 86604 57836 86605 57900
rect 86539 57835 86605 57836
rect 87643 57900 87709 57901
rect 87643 57836 87644 57900
rect 87708 57836 87709 57900
rect 87643 57835 87709 57836
rect 88379 57900 88445 57901
rect 88379 57836 88380 57900
rect 88444 57836 88445 57900
rect 88379 57835 88445 57836
rect 88747 57900 88813 57901
rect 88747 57836 88748 57900
rect 88812 57836 88813 57900
rect 88747 57835 88813 57836
rect 90035 57900 90101 57901
rect 90035 57836 90036 57900
rect 90100 57836 90101 57900
rect 90035 57835 90101 57836
rect 90771 57900 90837 57901
rect 90771 57836 90772 57900
rect 90836 57836 90837 57900
rect 90771 57835 90837 57836
rect 91323 57900 91389 57901
rect 91323 57836 91324 57900
rect 91388 57836 91389 57900
rect 91323 57835 91389 57836
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 58000
rect 93350 57901 93410 59470
rect 93718 57901 93778 59470
rect 95926 59397 95986 59606
rect 96048 59530 96108 60106
rect 97000 59666 97060 60106
rect 97000 59606 97090 59666
rect 96048 59470 96354 59530
rect 95923 59396 95989 59397
rect 95923 59332 95924 59396
rect 95988 59332 95989 59396
rect 95923 59331 95989 59332
rect 93347 57900 93413 57901
rect 93347 57836 93348 57900
rect 93412 57836 93413 57900
rect 93347 57835 93413 57836
rect 93715 57900 93781 57901
rect 93715 57836 93716 57900
rect 93780 57836 93781 57900
rect 93715 57835 93781 57836
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 25174 96134 58000
rect 96294 57085 96354 59470
rect 97030 59397 97090 59606
rect 98088 59530 98148 60106
rect 98496 59530 98556 60106
rect 99448 59805 99508 60106
rect 99445 59804 99511 59805
rect 99445 59740 99446 59804
rect 99510 59740 99511 59804
rect 99445 59739 99511 59740
rect 100672 59666 100732 60106
rect 101080 59669 101140 60106
rect 101077 59668 101143 59669
rect 100672 59606 100770 59666
rect 100710 59533 100770 59606
rect 101077 59604 101078 59668
rect 101142 59604 101143 59668
rect 101077 59603 101143 59604
rect 100707 59532 100773 59533
rect 98088 59470 98194 59530
rect 98496 59470 98562 59530
rect 97027 59396 97093 59397
rect 97027 59332 97028 59396
rect 97092 59332 97093 59396
rect 97027 59331 97093 59332
rect 98134 57901 98194 59470
rect 98131 57900 98197 57901
rect 98131 57836 98132 57900
rect 98196 57836 98197 57900
rect 98131 57835 98197 57836
rect 98502 57221 98562 59470
rect 100707 59468 100708 59532
rect 100772 59468 100773 59532
rect 101760 59530 101820 60106
rect 102848 59669 102908 60106
rect 102845 59668 102911 59669
rect 102845 59604 102846 59668
rect 102910 59604 102911 59668
rect 102845 59603 102911 59604
rect 103528 59530 103588 60106
rect 103936 59669 103996 60106
rect 103933 59668 103999 59669
rect 103933 59604 103934 59668
rect 103998 59604 103999 59668
rect 103933 59603 103999 59604
rect 105296 59530 105356 60106
rect 105976 59530 106036 60106
rect 101760 59470 101874 59530
rect 103528 59470 103898 59530
rect 105296 59470 105370 59530
rect 100707 59467 100773 59468
rect 101814 59397 101874 59470
rect 101811 59396 101877 59397
rect 101811 59332 101812 59396
rect 101876 59332 101877 59396
rect 101811 59331 101877 59332
rect 98499 57220 98565 57221
rect 98499 57156 98500 57220
rect 98564 57156 98565 57220
rect 98499 57155 98565 57156
rect 96291 57084 96357 57085
rect 96291 57020 96292 57084
rect 96356 57020 96357 57084
rect 96291 57019 96357 57020
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 28894 99854 58000
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 32614 103574 58000
rect 103838 57357 103898 59470
rect 103835 57356 103901 57357
rect 103835 57292 103836 57356
rect 103900 57292 103901 57356
rect 103835 57291 103901 57292
rect 105310 56269 105370 59470
rect 105862 59470 106036 59530
rect 106384 59530 106444 60106
rect 107608 59530 107668 60106
rect 108288 59530 108348 60106
rect 108696 59530 108756 60106
rect 109784 59530 109844 60106
rect 106384 59470 106474 59530
rect 105862 57085 105922 59470
rect 106414 57901 106474 59470
rect 107518 59470 107668 59530
rect 108254 59470 108348 59530
rect 108622 59470 108756 59530
rect 109542 59470 109844 59530
rect 111008 59530 111068 60106
rect 111144 59530 111204 60106
rect 112232 59530 112292 60106
rect 113320 59530 113380 60106
rect 113592 59805 113652 60106
rect 113589 59804 113655 59805
rect 113589 59740 113590 59804
rect 113654 59740 113655 59804
rect 113589 59739 113655 59740
rect 114408 59530 114468 60106
rect 111008 59470 111074 59530
rect 111144 59470 111258 59530
rect 107518 57901 107578 59470
rect 108254 58581 108314 59470
rect 108251 58580 108317 58581
rect 108251 58516 108252 58580
rect 108316 58516 108317 58580
rect 108251 58515 108317 58516
rect 108622 57901 108682 59470
rect 106411 57900 106477 57901
rect 106411 57836 106412 57900
rect 106476 57836 106477 57900
rect 106411 57835 106477 57836
rect 107515 57900 107581 57901
rect 107515 57836 107516 57900
rect 107580 57836 107581 57900
rect 107515 57835 107581 57836
rect 108619 57900 108685 57901
rect 108619 57836 108620 57900
rect 108684 57836 108685 57900
rect 108619 57835 108685 57836
rect 109542 57629 109602 59470
rect 111014 58445 111074 59470
rect 111198 59397 111258 59470
rect 112118 59470 112292 59530
rect 113222 59470 113380 59530
rect 114326 59470 114468 59530
rect 115768 59530 115828 60106
rect 116040 59530 116100 60106
rect 116992 59530 117052 60106
rect 118080 59530 118140 60106
rect 118488 59530 118548 60106
rect 119168 59530 119228 60106
rect 115768 59470 115858 59530
rect 111195 59396 111261 59397
rect 111195 59332 111196 59396
rect 111260 59332 111261 59396
rect 111195 59331 111261 59332
rect 111011 58444 111077 58445
rect 111011 58380 111012 58444
rect 111076 58380 111077 58444
rect 111011 58379 111077 58380
rect 109539 57628 109605 57629
rect 109539 57564 109540 57628
rect 109604 57564 109605 57628
rect 109539 57563 109605 57564
rect 105859 57084 105925 57085
rect 105859 57020 105860 57084
rect 105924 57020 105925 57084
rect 105859 57019 105925 57020
rect 105307 56268 105373 56269
rect 105307 56204 105308 56268
rect 105372 56204 105373 56268
rect 105307 56203 105373 56204
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 39454 110414 58000
rect 112118 57901 112178 59470
rect 113222 57901 113282 59470
rect 112115 57900 112181 57901
rect 112115 57836 112116 57900
rect 112180 57836 112181 57900
rect 112115 57835 112181 57836
rect 113219 57900 113285 57901
rect 113219 57836 113220 57900
rect 113284 57836 113285 57900
rect 113219 57835 113285 57836
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 43174 114134 58000
rect 114326 57629 114386 59470
rect 115798 57629 115858 59470
rect 115982 59470 116100 59530
rect 116902 59470 117052 59530
rect 118006 59470 118140 59530
rect 118374 59470 118548 59530
rect 119110 59470 119228 59530
rect 120936 59530 120996 60106
rect 123520 59530 123580 60106
rect 125968 59530 126028 60106
rect 120936 59470 121010 59530
rect 123520 59470 123586 59530
rect 115982 59397 116042 59470
rect 115979 59396 116045 59397
rect 115979 59332 115980 59396
rect 116044 59332 116045 59396
rect 115979 59331 116045 59332
rect 116902 57629 116962 59470
rect 114323 57628 114389 57629
rect 114323 57564 114324 57628
rect 114388 57564 114389 57628
rect 114323 57563 114389 57564
rect 115795 57628 115861 57629
rect 115795 57564 115796 57628
rect 115860 57564 115861 57628
rect 115795 57563 115861 57564
rect 116899 57628 116965 57629
rect 116899 57564 116900 57628
rect 116964 57564 116965 57628
rect 116899 57563 116965 57564
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 46894 117854 58000
rect 118006 57629 118066 59470
rect 118003 57628 118069 57629
rect 118003 57564 118004 57628
rect 118068 57564 118069 57628
rect 118003 57563 118069 57564
rect 118374 57493 118434 59470
rect 119110 57629 119170 59470
rect 120950 58717 121010 59470
rect 120947 58716 121013 58717
rect 120947 58652 120948 58716
rect 121012 58652 121013 58716
rect 120947 58651 121013 58652
rect 119107 57628 119173 57629
rect 119107 57564 119108 57628
rect 119172 57564 119173 57628
rect 119107 57563 119173 57564
rect 118371 57492 118437 57493
rect 118371 57428 118372 57492
rect 118436 57428 118437 57492
rect 118371 57427 118437 57428
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 50614 121574 58000
rect 123526 57901 123586 59470
rect 125918 59470 126028 59530
rect 128280 59530 128340 60106
rect 131000 59530 131060 60106
rect 128280 59470 128738 59530
rect 123523 57900 123589 57901
rect 123523 57836 123524 57900
rect 123588 57836 123589 57900
rect 123523 57835 123589 57836
rect 125918 57765 125978 59470
rect 125915 57764 125981 57765
rect 125915 57700 125916 57764
rect 125980 57700 125981 57764
rect 125915 57699 125981 57700
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 58000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 128678 56677 128738 59470
rect 130886 59470 131060 59530
rect 133448 59530 133508 60106
rect 135896 59530 135956 60106
rect 138480 59530 138540 60106
rect 140928 59530 140988 60106
rect 133448 59470 133522 59530
rect 130886 57901 130946 59470
rect 130883 57900 130949 57901
rect 130883 57836 130884 57900
rect 130948 57836 130949 57900
rect 130883 57835 130949 57836
rect 128675 56676 128741 56677
rect 128675 56612 128676 56676
rect 128740 56612 128741 56676
rect 128675 56611 128741 56612
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 25174 132134 58000
rect 133462 57901 133522 59470
rect 135854 59470 135956 59530
rect 138430 59470 138540 59530
rect 140822 59470 140988 59530
rect 143512 59530 143572 60106
rect 145960 59530 146020 60106
rect 143512 59470 143642 59530
rect 135854 58853 135914 59470
rect 138430 58989 138490 59470
rect 140822 59125 140882 59470
rect 143582 59261 143642 59470
rect 145606 59470 146020 59530
rect 148544 59530 148604 60106
rect 150992 59530 151052 60106
rect 153440 59530 153500 60106
rect 148544 59470 148610 59530
rect 143579 59260 143645 59261
rect 143579 59196 143580 59260
rect 143644 59196 143645 59260
rect 143579 59195 143645 59196
rect 140819 59124 140885 59125
rect 140819 59060 140820 59124
rect 140884 59060 140885 59124
rect 140819 59059 140885 59060
rect 138427 58988 138493 58989
rect 138427 58924 138428 58988
rect 138492 58924 138493 58988
rect 138427 58923 138493 58924
rect 135851 58852 135917 58853
rect 135851 58788 135852 58852
rect 135916 58788 135917 58852
rect 135851 58787 135917 58788
rect 133459 57900 133525 57901
rect 133459 57836 133460 57900
rect 133524 57836 133525 57900
rect 133459 57835 133525 57836
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 28894 135854 58000
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 32614 139574 58000
rect 145606 57901 145666 59470
rect 148550 59261 148610 59470
rect 150942 59470 151052 59530
rect 153334 59470 153500 59530
rect 155888 59530 155948 60106
rect 158472 59530 158532 60106
rect 160920 59530 160980 60106
rect 163368 59530 163428 60106
rect 165952 59530 166012 60106
rect 183224 59530 183284 60106
rect 155888 59470 155970 59530
rect 158472 59470 158546 59530
rect 150942 59261 151002 59470
rect 148547 59260 148613 59261
rect 148547 59196 148548 59260
rect 148612 59196 148613 59260
rect 148547 59195 148613 59196
rect 150939 59260 151005 59261
rect 150939 59196 150940 59260
rect 151004 59196 151005 59260
rect 150939 59195 151005 59196
rect 153334 58173 153394 59470
rect 153331 58172 153397 58173
rect 153331 58108 153332 58172
rect 153396 58108 153397 58172
rect 153331 58107 153397 58108
rect 145603 57900 145669 57901
rect 145603 57836 145604 57900
rect 145668 57836 145669 57900
rect 145603 57835 145669 57836
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 39454 146414 58000
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 43174 150134 58000
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 46894 153854 58000
rect 155910 57629 155970 59470
rect 155907 57628 155973 57629
rect 155907 57564 155908 57628
rect 155972 57564 155973 57628
rect 155907 57563 155973 57564
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 50614 157574 58000
rect 158486 57901 158546 59470
rect 160878 59470 160980 59530
rect 163270 59470 163428 59530
rect 165846 59470 166012 59530
rect 183142 59470 183284 59530
rect 183360 59530 183420 60106
rect 183360 59470 183570 59530
rect 158483 57900 158549 57901
rect 158483 57836 158484 57900
rect 158548 57836 158549 57900
rect 158483 57835 158549 57836
rect 160878 57629 160938 59470
rect 160875 57628 160941 57629
rect 160875 57564 160876 57628
rect 160940 57564 160941 57628
rect 160875 57563 160941 57564
rect 163270 56677 163330 59470
rect 163794 57454 164414 58000
rect 165846 57629 165906 59470
rect 165843 57628 165909 57629
rect 165843 57564 165844 57628
rect 165908 57564 165909 57628
rect 165843 57563 165909 57564
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163267 56676 163333 56677
rect 163267 56612 163268 56676
rect 163332 56612 163333 56676
rect 163267 56611 163333 56612
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 25174 168134 58000
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 28894 171854 58000
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 32614 175574 58000
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 39454 182414 58000
rect 183142 57901 183202 59470
rect 183139 57900 183205 57901
rect 183139 57836 183140 57900
rect 183204 57836 183205 57900
rect 183139 57835 183205 57836
rect 183510 57765 183570 59470
rect 197862 58717 197922 478211
rect 198046 59397 198106 478483
rect 198230 164117 198290 478755
rect 198595 477732 198661 477733
rect 198595 477668 198596 477732
rect 198660 477668 198661 477732
rect 198595 477667 198661 477668
rect 198227 164116 198293 164117
rect 198227 164052 198228 164116
rect 198292 164052 198293 164116
rect 198227 164051 198293 164052
rect 198043 59396 198109 59397
rect 198043 59332 198044 59396
rect 198108 59332 198109 59396
rect 198043 59331 198109 59332
rect 198598 59125 198658 477667
rect 198782 394637 198842 478891
rect 205403 478548 205469 478549
rect 205403 478484 205404 478548
rect 205468 478484 205469 478548
rect 205403 478483 205469 478484
rect 200619 478412 200685 478413
rect 200619 478348 200620 478412
rect 200684 478348 200685 478412
rect 200619 478347 200685 478348
rect 198963 474060 199029 474061
rect 198963 473996 198964 474060
rect 199028 473996 199029 474060
rect 198963 473995 199029 473996
rect 198779 394636 198845 394637
rect 198779 394572 198780 394636
rect 198844 394572 198845 394636
rect 198779 394571 198845 394572
rect 198779 392052 198845 392053
rect 198779 391988 198780 392052
rect 198844 391988 198845 392052
rect 198779 391987 198845 391988
rect 198782 267613 198842 391987
rect 198966 388517 199026 473995
rect 199794 470514 200414 478000
rect 199794 470278 199826 470514
rect 200062 470278 200146 470514
rect 200382 470278 200414 470514
rect 199794 470194 200414 470278
rect 199794 469958 199826 470194
rect 200062 469958 200146 470194
rect 200382 469958 200414 470194
rect 199147 458828 199213 458829
rect 199147 458764 199148 458828
rect 199212 458764 199213 458828
rect 199147 458763 199213 458764
rect 199150 390693 199210 458763
rect 199794 453454 200414 469958
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199331 392188 199397 392189
rect 199331 392124 199332 392188
rect 199396 392124 199397 392188
rect 199331 392123 199397 392124
rect 199147 390692 199213 390693
rect 199147 390628 199148 390692
rect 199212 390628 199213 390692
rect 199147 390627 199213 390628
rect 199147 389060 199213 389061
rect 199147 388996 199148 389060
rect 199212 388996 199213 389060
rect 199147 388995 199213 388996
rect 198963 388516 199029 388517
rect 198963 388452 198964 388516
rect 199028 388452 199029 388516
rect 198963 388451 199029 388452
rect 199150 373965 199210 388995
rect 199147 373964 199213 373965
rect 199147 373900 199148 373964
rect 199212 373900 199213 373964
rect 199147 373899 199213 373900
rect 199150 372741 199210 373899
rect 199334 373829 199394 392123
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199331 373828 199397 373829
rect 199331 373764 199332 373828
rect 199396 373764 199397 373828
rect 199331 373763 199397 373764
rect 199147 372740 199213 372741
rect 199147 372676 199148 372740
rect 199212 372676 199213 372740
rect 199147 372675 199213 372676
rect 199794 364394 200414 380898
rect 199794 364158 199826 364394
rect 200062 364158 200146 364394
rect 200382 364158 200414 364394
rect 199794 364074 200414 364158
rect 199794 363838 199826 364074
rect 200062 363838 200146 364074
rect 200382 363838 200414 364074
rect 199794 345454 200414 363838
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 198779 267612 198845 267613
rect 198779 267548 198780 267612
rect 198844 267548 198845 267612
rect 198779 267547 198845 267548
rect 199794 256394 200414 272898
rect 199794 256158 199826 256394
rect 200062 256158 200146 256394
rect 200382 256158 200414 256394
rect 199794 256074 200414 256158
rect 199794 255838 199826 256074
rect 200062 255838 200146 256074
rect 200382 255838 200414 256074
rect 199794 237454 200414 255838
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 148394 200414 164898
rect 199794 148158 199826 148394
rect 200062 148158 200146 148394
rect 200382 148158 200414 148394
rect 199794 148074 200414 148158
rect 199794 147838 199826 148074
rect 200062 147838 200146 148074
rect 200382 147838 200414 148074
rect 199794 129454 200414 147838
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 198595 59124 198661 59125
rect 198595 59060 198596 59124
rect 198660 59060 198661 59124
rect 198595 59059 198661 59060
rect 197859 58716 197925 58717
rect 197859 58652 197860 58716
rect 197924 58652 197925 58716
rect 197859 58651 197925 58652
rect 183507 57764 183573 57765
rect 183507 57700 183508 57764
rect 183572 57700 183573 57764
rect 183507 57699 183573 57700
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 43174 186134 58000
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 46894 189854 58000
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 50614 193574 58000
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 200622 56405 200682 478347
rect 200987 478276 201053 478277
rect 200987 478212 200988 478276
rect 201052 478212 201053 478276
rect 200987 478211 201053 478212
rect 200803 459508 200869 459509
rect 200803 459444 200804 459508
rect 200868 459444 200869 459508
rect 200803 459443 200869 459444
rect 200806 174997 200866 459443
rect 200990 375325 201050 478211
rect 202091 478140 202157 478141
rect 202091 478076 202092 478140
rect 202156 478076 202157 478140
rect 202091 478075 202157 478076
rect 201355 477732 201421 477733
rect 201355 477668 201356 477732
rect 201420 477668 201421 477732
rect 201355 477667 201421 477668
rect 200987 375324 201053 375325
rect 200987 375260 200988 375324
rect 201052 375260 201053 375324
rect 200987 375259 201053 375260
rect 200803 174996 200869 174997
rect 200803 174932 200804 174996
rect 200868 174932 200869 174996
rect 200803 174931 200869 174932
rect 201358 59261 201418 477667
rect 201355 59260 201421 59261
rect 201355 59196 201356 59260
rect 201420 59196 201421 59260
rect 201355 59195 201421 59196
rect 202094 58581 202154 478075
rect 202643 478004 202709 478005
rect 202643 477940 202644 478004
rect 202708 477940 202709 478004
rect 202643 477939 202709 477940
rect 202275 463044 202341 463045
rect 202275 462980 202276 463044
rect 202340 462980 202341 463044
rect 202275 462979 202341 462980
rect 202091 58580 202157 58581
rect 202091 58516 202092 58580
rect 202156 58516 202157 58580
rect 202091 58515 202157 58516
rect 202278 57493 202338 462979
rect 202459 460868 202525 460869
rect 202459 460804 202460 460868
rect 202524 460804 202525 460868
rect 202459 460803 202525 460804
rect 202462 163981 202522 460803
rect 202646 375325 202706 477939
rect 203514 474234 204134 478000
rect 203514 473998 203546 474234
rect 203782 473998 203866 474234
rect 204102 473998 204134 474234
rect 203514 473914 204134 473998
rect 203514 473678 203546 473914
rect 203782 473678 203866 473914
rect 204102 473678 204134 473914
rect 203195 466172 203261 466173
rect 203195 466108 203196 466172
rect 203260 466108 203261 466172
rect 203195 466107 203261 466108
rect 203011 463180 203077 463181
rect 203011 463116 203012 463180
rect 203076 463116 203077 463180
rect 203011 463115 203077 463116
rect 202643 375324 202709 375325
rect 202643 375260 202644 375324
rect 202708 375260 202709 375324
rect 202643 375259 202709 375260
rect 203014 164253 203074 463115
rect 203011 164252 203077 164253
rect 203011 164188 203012 164252
rect 203076 164188 203077 164252
rect 203011 164187 203077 164188
rect 202459 163980 202525 163981
rect 202459 163916 202460 163980
rect 202524 163916 202525 163980
rect 202459 163915 202525 163916
rect 203198 162485 203258 466107
rect 203514 457174 204134 473678
rect 204851 471340 204917 471341
rect 204851 471276 204852 471340
rect 204916 471276 204917 471340
rect 204851 471275 204917 471276
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 366234 204134 384618
rect 203514 365998 203546 366234
rect 203782 365998 203866 366234
rect 204102 365998 204134 366234
rect 203514 365914 204134 365998
rect 203514 365678 203546 365914
rect 203782 365678 203866 365914
rect 204102 365678 204134 365914
rect 203514 349174 204134 365678
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 277174 204134 312618
rect 203514 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 204134 277174
rect 203514 276854 204134 276938
rect 203514 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 204134 276854
rect 203514 260114 204134 276618
rect 203514 259878 203546 260114
rect 203782 259878 203866 260114
rect 204102 259878 204134 260114
rect 203514 259794 204134 259878
rect 203514 259558 203546 259794
rect 203782 259558 203866 259794
rect 204102 259558 204134 259794
rect 203514 241174 204134 259558
rect 203514 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 204134 241174
rect 203514 240854 204134 240938
rect 203514 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 204134 240854
rect 203514 205174 204134 240618
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203195 162484 203261 162485
rect 203195 162420 203196 162484
rect 203260 162420 203261 162484
rect 203195 162419 203261 162420
rect 203514 152114 204134 168618
rect 203514 151878 203546 152114
rect 203782 151878 203866 152114
rect 204102 151878 204134 152114
rect 203514 151794 204134 151878
rect 203514 151558 203546 151794
rect 203782 151558 203866 151794
rect 204102 151558 204134 151794
rect 203514 133174 204134 151558
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 202275 57492 202341 57493
rect 202275 57428 202276 57492
rect 202340 57428 202341 57492
rect 202275 57427 202341 57428
rect 200619 56404 200685 56405
rect 200619 56340 200620 56404
rect 200684 56340 200685 56404
rect 200619 56339 200685 56340
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 25174 204134 60618
rect 204854 57357 204914 471275
rect 205219 460732 205285 460733
rect 205219 460668 205220 460732
rect 205284 460668 205285 460732
rect 205219 460667 205285 460668
rect 205035 460324 205101 460325
rect 205035 460260 205036 460324
rect 205100 460260 205101 460324
rect 205035 460259 205101 460260
rect 205038 68101 205098 460259
rect 205222 164389 205282 460667
rect 205406 456925 205466 478483
rect 205403 456924 205469 456925
rect 205403 456860 205404 456924
rect 205468 456860 205469 456924
rect 205403 456859 205469 456860
rect 205219 164388 205285 164389
rect 205219 164324 205220 164388
rect 205284 164324 205285 164388
rect 205219 164323 205285 164324
rect 205035 68100 205101 68101
rect 205035 68036 205036 68100
rect 205100 68036 205101 68100
rect 205035 68035 205101 68036
rect 204851 57356 204917 57357
rect 204851 57292 204852 57356
rect 204916 57292 204917 57356
rect 204851 57291 204917 57292
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 206142 3909 206202 479435
rect 206875 478684 206941 478685
rect 206875 478620 206876 478684
rect 206940 478620 206941 478684
rect 206875 478619 206941 478620
rect 206507 478412 206573 478413
rect 206507 478348 206508 478412
rect 206572 478348 206573 478412
rect 206507 478347 206573 478348
rect 206323 470116 206389 470117
rect 206323 470052 206324 470116
rect 206388 470052 206389 470116
rect 206323 470051 206389 470052
rect 206326 161805 206386 470051
rect 206510 375325 206570 478347
rect 206507 375324 206573 375325
rect 206507 375260 206508 375324
rect 206572 375260 206573 375324
rect 206507 375259 206573 375260
rect 206323 161804 206389 161805
rect 206323 161740 206324 161804
rect 206388 161740 206389 161804
rect 206323 161739 206389 161740
rect 206878 58989 206938 478619
rect 207234 470078 207854 478000
rect 207234 469842 207266 470078
rect 207502 469842 207586 470078
rect 207822 469842 207854 470078
rect 207234 469758 207854 469842
rect 207234 469522 207266 469758
rect 207502 469522 207586 469758
rect 207822 469522 207854 469758
rect 207059 467260 207125 467261
rect 207059 467196 207060 467260
rect 207124 467196 207125 467260
rect 207059 467195 207125 467196
rect 207062 407829 207122 467195
rect 207234 460894 207854 469522
rect 207979 464404 208045 464405
rect 207979 464340 207980 464404
rect 208044 464340 208045 464404
rect 207979 464339 208045 464340
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207059 407828 207125 407829
rect 207059 407764 207060 407828
rect 207124 407764 207125 407828
rect 207059 407763 207125 407764
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 369954 207854 388338
rect 207234 369718 207266 369954
rect 207502 369718 207586 369954
rect 207822 369718 207854 369954
rect 207234 369634 207854 369718
rect 207234 369398 207266 369634
rect 207502 369398 207586 369634
rect 207822 369398 207854 369634
rect 207234 352894 207854 369398
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 280894 207854 316338
rect 207234 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 207854 280894
rect 207234 280574 207854 280658
rect 207234 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 207854 280574
rect 207234 261954 207854 280338
rect 207234 261718 207266 261954
rect 207502 261718 207586 261954
rect 207822 261718 207854 261954
rect 207234 261634 207854 261718
rect 207234 261398 207266 261634
rect 207502 261398 207586 261634
rect 207822 261398 207854 261634
rect 207234 244894 207854 261398
rect 207234 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 207854 244894
rect 207234 244574 207854 244658
rect 207234 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 207854 244574
rect 207234 208894 207854 244338
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 153954 207854 172338
rect 207982 162621 208042 464339
rect 207979 162620 208045 162621
rect 207979 162556 207980 162620
rect 208044 162556 208045 162620
rect 207979 162555 208045 162556
rect 207234 153718 207266 153954
rect 207502 153718 207586 153954
rect 207822 153718 207854 153954
rect 207234 153634 207854 153718
rect 207234 153398 207266 153634
rect 207502 153398 207586 153634
rect 207822 153398 207854 153634
rect 207234 136894 207854 153398
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 206875 58988 206941 58989
rect 206875 58924 206876 58988
rect 206940 58924 206941 58988
rect 206875 58923 206941 58924
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 206139 3908 206205 3909
rect 206139 3844 206140 3908
rect 206204 3844 206205 3908
rect 206139 3843 206205 3844
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 -5146 207854 28338
rect 208902 4045 208962 479571
rect 214787 478684 214853 478685
rect 214787 478620 214788 478684
rect 214852 478620 214853 478684
rect 214787 478619 214853 478620
rect 209267 478548 209333 478549
rect 209267 478484 209268 478548
rect 209332 478484 209333 478548
rect 209267 478483 209333 478484
rect 209083 467124 209149 467125
rect 209083 467060 209084 467124
rect 209148 467060 209149 467124
rect 209083 467059 209149 467060
rect 209086 57629 209146 467059
rect 209270 369205 209330 478483
rect 213683 478140 213749 478141
rect 213683 478076 213684 478140
rect 213748 478076 213749 478140
rect 213683 478075 213749 478076
rect 209819 476780 209885 476781
rect 209819 476716 209820 476780
rect 209884 476716 209885 476780
rect 209819 476715 209885 476716
rect 209822 375325 209882 476715
rect 210371 474060 210437 474061
rect 210371 473996 210372 474060
rect 210436 473996 210437 474060
rect 210371 473995 210437 473996
rect 210003 468756 210069 468757
rect 210003 468692 210004 468756
rect 210068 468692 210069 468756
rect 210003 468691 210069 468692
rect 209819 375324 209885 375325
rect 209819 375260 209820 375324
rect 209884 375260 209885 375324
rect 209819 375259 209885 375260
rect 210006 372741 210066 468691
rect 210003 372740 210069 372741
rect 210003 372676 210004 372740
rect 210068 372676 210069 372740
rect 210003 372675 210069 372676
rect 209267 369204 209333 369205
rect 209267 369140 209268 369204
rect 209332 369140 209333 369204
rect 209267 369139 209333 369140
rect 209083 57628 209149 57629
rect 209083 57564 209084 57628
rect 209148 57564 209149 57628
rect 209083 57563 209149 57564
rect 208899 4044 208965 4045
rect 208899 3980 208900 4044
rect 208964 3980 208965 4044
rect 208899 3979 208965 3980
rect 210374 3229 210434 473995
rect 210954 464614 211574 478000
rect 213315 474332 213381 474333
rect 213315 474268 213316 474332
rect 213380 474268 213381 474332
rect 213315 474267 213381 474268
rect 212027 472564 212093 472565
rect 212027 472500 212028 472564
rect 212092 472500 212093 472564
rect 212027 472499 212093 472500
rect 211843 469980 211909 469981
rect 211843 469916 211844 469980
rect 211908 469916 211909 469980
rect 211843 469915 211909 469916
rect 211659 468484 211725 468485
rect 211659 468420 211660 468484
rect 211724 468420 211725 468484
rect 211659 468419 211725 468420
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 356614 211574 392058
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 284614 211574 320058
rect 210954 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 211574 284614
rect 210954 284294 211574 284378
rect 210954 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 211574 284294
rect 210954 265674 211574 284058
rect 210954 265438 210986 265674
rect 211222 265438 211306 265674
rect 211542 265438 211574 265674
rect 210954 265354 211574 265438
rect 210954 265118 210986 265354
rect 211222 265118 211306 265354
rect 211542 265118 211574 265354
rect 210954 248614 211574 265118
rect 210954 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 211574 248614
rect 210954 248294 211574 248378
rect 210954 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 211574 248294
rect 210954 212614 211574 248058
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 157674 211574 176058
rect 210954 157438 210986 157674
rect 211222 157438 211306 157674
rect 211542 157438 211574 157674
rect 210954 157354 211574 157438
rect 210954 157118 210986 157354
rect 211222 157118 211306 157354
rect 211542 157118 211574 157354
rect 210954 140614 211574 157118
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 211662 57085 211722 468419
rect 211846 375325 211906 469915
rect 212030 382397 212090 472499
rect 212579 469844 212645 469845
rect 212579 469780 212580 469844
rect 212644 469780 212645 469844
rect 212579 469779 212645 469780
rect 212027 382396 212093 382397
rect 212027 382332 212028 382396
rect 212092 382332 212093 382396
rect 212027 382331 212093 382332
rect 211843 375324 211909 375325
rect 211843 375260 211844 375324
rect 211908 375260 211909 375324
rect 211843 375259 211909 375260
rect 212582 369205 212642 469779
rect 213131 462908 213197 462909
rect 213131 462844 213132 462908
rect 213196 462844 213197 462908
rect 213131 462843 213197 462844
rect 212579 369204 212645 369205
rect 212579 369140 212580 369204
rect 212644 369140 212645 369204
rect 212579 369139 212645 369140
rect 213134 57221 213194 462843
rect 213318 162349 213378 474267
rect 213315 162348 213381 162349
rect 213315 162284 213316 162348
rect 213380 162284 213381 162348
rect 213315 162283 213381 162284
rect 213686 58853 213746 478075
rect 214419 474196 214485 474197
rect 214419 474132 214420 474196
rect 214484 474132 214485 474196
rect 214419 474131 214485 474132
rect 213683 58852 213749 58853
rect 213683 58788 213684 58852
rect 213748 58788 213749 58852
rect 213683 58787 213749 58788
rect 214422 57765 214482 474131
rect 214603 468620 214669 468621
rect 214603 468556 214604 468620
rect 214668 468556 214669 468620
rect 214603 468555 214669 468556
rect 214419 57764 214485 57765
rect 214419 57700 214420 57764
rect 214484 57700 214485 57764
rect 214419 57699 214485 57700
rect 213131 57220 213197 57221
rect 213131 57156 213132 57220
rect 213196 57156 213197 57220
rect 213131 57155 213197 57156
rect 211659 57084 211725 57085
rect 211659 57020 211660 57084
rect 211724 57020 211725 57084
rect 211659 57019 211725 57020
rect 214606 56677 214666 468555
rect 214790 369885 214850 478619
rect 219203 478276 219269 478277
rect 219203 478212 219204 478276
rect 219268 478212 219269 478276
rect 219203 478211 219269 478212
rect 216995 477732 217061 477733
rect 216995 477668 216996 477732
rect 217060 477668 217061 477732
rect 216995 477667 217061 477668
rect 215339 475556 215405 475557
rect 215339 475492 215340 475556
rect 215404 475492 215405 475556
rect 215339 475491 215405 475492
rect 214787 369884 214853 369885
rect 214787 369820 214788 369884
rect 214852 369820 214853 369884
rect 214787 369819 214853 369820
rect 215342 266525 215402 475491
rect 215523 471204 215589 471205
rect 215523 471140 215524 471204
rect 215588 471140 215589 471204
rect 215523 471139 215589 471140
rect 215339 266524 215405 266525
rect 215339 266460 215340 266524
rect 215404 266460 215405 266524
rect 215339 266459 215405 266460
rect 215526 266389 215586 471139
rect 215891 460596 215957 460597
rect 215891 460532 215892 460596
rect 215956 460532 215957 460596
rect 215891 460531 215957 460532
rect 215523 266388 215589 266389
rect 215523 266324 215524 266388
rect 215588 266324 215589 266388
rect 215523 266323 215589 266324
rect 215894 162213 215954 460531
rect 216998 372741 217058 477667
rect 217547 477596 217613 477597
rect 217547 477532 217548 477596
rect 217612 477532 217613 477596
rect 217547 477531 217613 477532
rect 217179 472700 217245 472701
rect 217179 472636 217180 472700
rect 217244 472636 217245 472700
rect 217179 472635 217245 472636
rect 216995 372740 217061 372741
rect 216995 372676 216996 372740
rect 217060 372676 217061 372740
rect 216995 372675 217061 372676
rect 216995 370972 217061 370973
rect 216995 370908 216996 370972
rect 217060 370908 217061 370972
rect 216995 370907 217061 370908
rect 216998 267885 217058 370907
rect 216995 267884 217061 267885
rect 216995 267820 216996 267884
rect 217060 267820 217061 267884
rect 216995 267819 217061 267820
rect 217182 267205 217242 472635
rect 217363 463316 217429 463317
rect 217363 463252 217364 463316
rect 217428 463252 217429 463316
rect 217363 463251 217429 463252
rect 217366 268973 217426 463251
rect 217550 373693 217610 477531
rect 217794 471454 218414 478000
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 460308 218414 470898
rect 218651 460460 218717 460461
rect 218651 460396 218652 460460
rect 218716 460396 218717 460460
rect 218651 460395 218717 460396
rect 217547 373692 217613 373693
rect 217547 373628 217548 373692
rect 217612 373628 217613 373692
rect 217547 373627 217613 373628
rect 217550 370973 217610 373627
rect 217547 370972 217613 370973
rect 217547 370908 217548 370972
rect 217612 370908 217613 370972
rect 217547 370907 217613 370908
rect 217794 363454 218414 373000
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 355308 218414 362898
rect 217363 268972 217429 268973
rect 217363 268908 217364 268972
rect 217428 268908 217429 268972
rect 217363 268907 217429 268908
rect 217547 268836 217613 268837
rect 217547 268772 217548 268836
rect 217612 268772 217613 268836
rect 217547 268771 217613 268772
rect 217550 268021 217610 268771
rect 217547 268020 217613 268021
rect 217547 267956 217548 268020
rect 217612 267956 217613 268020
rect 217547 267955 217613 267956
rect 217179 267204 217245 267205
rect 217179 267140 217180 267204
rect 217244 267140 217245 267204
rect 217179 267139 217245 267140
rect 215891 162212 215957 162213
rect 215891 162148 215892 162212
rect 215956 162148 215957 162212
rect 215891 162147 215957 162148
rect 217550 161125 217610 267955
rect 217794 255454 218414 268000
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 250308 218414 254898
rect 217547 161124 217613 161125
rect 217547 161060 217548 161124
rect 217612 161060 217613 161124
rect 217547 161059 217613 161060
rect 217363 148340 217429 148341
rect 217363 148276 217364 148340
rect 217428 148276 217429 148340
rect 217363 148275 217429 148276
rect 217179 146436 217245 146437
rect 217179 146372 217180 146436
rect 217244 146372 217245 146436
rect 217179 146371 217245 146372
rect 214603 56676 214669 56677
rect 214603 56612 214604 56676
rect 214668 56612 214669 56676
rect 214603 56611 214669 56612
rect 217182 55181 217242 146371
rect 217366 56269 217426 148275
rect 217550 58445 217610 161059
rect 217794 147454 218414 163000
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 145308 218414 146898
rect 218654 60621 218714 460395
rect 218835 460188 218901 460189
rect 218835 460124 218836 460188
rect 218900 460124 218901 460188
rect 218835 460123 218901 460124
rect 218838 163709 218898 460123
rect 218835 163708 218901 163709
rect 218835 163644 218836 163708
rect 218900 163644 218901 163708
rect 218835 163643 218901 163644
rect 219206 60621 219266 478211
rect 219939 477596 220005 477597
rect 219939 477532 219940 477596
rect 220004 477532 220005 477596
rect 219939 477531 220005 477532
rect 218651 60620 218717 60621
rect 218651 60556 218652 60620
rect 218716 60556 218717 60620
rect 218651 60555 218717 60556
rect 219203 60620 219269 60621
rect 219203 60556 219204 60620
rect 219268 60556 219269 60620
rect 219203 60555 219269 60556
rect 217547 58444 217613 58445
rect 217547 58380 217548 58444
rect 217612 58380 217613 58444
rect 217547 58379 217613 58380
rect 217363 56268 217429 56269
rect 217363 56204 217364 56268
rect 217428 56204 217429 56268
rect 217363 56203 217429 56204
rect 217179 55180 217245 55181
rect 217179 55116 217180 55180
rect 217244 55116 217245 55180
rect 217179 55115 217245 55116
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 210371 3228 210437 3229
rect 210371 3164 210372 3228
rect 210436 3164 210437 3228
rect 210371 3163 210437 3164
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 39454 218414 58000
rect 219942 56541 220002 477531
rect 221514 475174 222134 478000
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 460308 222134 474618
rect 225234 469138 225854 478000
rect 225234 468902 225266 469138
rect 225502 468902 225586 469138
rect 225822 468902 225854 469138
rect 225234 468818 225854 468902
rect 225234 468582 225266 468818
rect 225502 468582 225586 468818
rect 225822 468582 225854 468818
rect 225234 460308 225854 468582
rect 228954 465554 229574 478000
rect 228954 465318 228986 465554
rect 229222 465318 229306 465554
rect 229542 465318 229574 465554
rect 228954 465234 229574 465318
rect 228954 464998 228986 465234
rect 229222 464998 229306 465234
rect 229542 464998 229574 465234
rect 228954 460308 229574 464998
rect 235794 470514 236414 478000
rect 235794 470278 235826 470514
rect 236062 470278 236146 470514
rect 236382 470278 236414 470514
rect 235794 470194 236414 470278
rect 235794 469958 235826 470194
rect 236062 469958 236146 470194
rect 236382 469958 236414 470194
rect 235794 460308 236414 469958
rect 239514 474234 240134 478000
rect 239514 473998 239546 474234
rect 239782 473998 239866 474234
rect 240102 473998 240134 474234
rect 239514 473914 240134 473998
rect 239514 473678 239546 473914
rect 239782 473678 239866 473914
rect 240102 473678 240134 473914
rect 239514 460308 240134 473678
rect 243234 470078 243854 478000
rect 243234 469842 243266 470078
rect 243502 469842 243586 470078
rect 243822 469842 243854 470078
rect 243234 469758 243854 469842
rect 243234 469522 243266 469758
rect 243502 469522 243586 469758
rect 243822 469522 243854 469758
rect 243234 460308 243854 469522
rect 246954 464614 247574 478000
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 460308 247574 464058
rect 253794 471454 254414 478000
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 460308 254414 470898
rect 257514 475174 258134 478000
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 460308 258134 474618
rect 261234 469138 261854 478000
rect 261234 468902 261266 469138
rect 261502 468902 261586 469138
rect 261822 468902 261854 469138
rect 261234 468818 261854 468902
rect 261234 468582 261266 468818
rect 261502 468582 261586 468818
rect 261822 468582 261854 468818
rect 261234 460308 261854 468582
rect 264954 465554 265574 478000
rect 264954 465318 264986 465554
rect 265222 465318 265306 465554
rect 265542 465318 265574 465554
rect 264954 465234 265574 465318
rect 264954 464998 264986 465234
rect 265222 464998 265306 465234
rect 265542 464998 265574 465234
rect 264954 460308 265574 464998
rect 271794 470514 272414 478000
rect 271794 470278 271826 470514
rect 272062 470278 272146 470514
rect 272382 470278 272414 470514
rect 271794 470194 272414 470278
rect 271794 469958 271826 470194
rect 272062 469958 272146 470194
rect 272382 469958 272414 470194
rect 271794 460308 272414 469958
rect 275514 474234 276134 478000
rect 275514 473998 275546 474234
rect 275782 473998 275866 474234
rect 276102 473998 276134 474234
rect 275514 473914 276134 473998
rect 275514 473678 275546 473914
rect 275782 473678 275866 473914
rect 276102 473678 276134 473914
rect 275514 460308 276134 473678
rect 279234 470078 279854 478000
rect 279234 469842 279266 470078
rect 279502 469842 279586 470078
rect 279822 469842 279854 470078
rect 279234 469758 279854 469842
rect 279234 469522 279266 469758
rect 279502 469522 279586 469758
rect 279822 469522 279854 469758
rect 279234 460308 279854 469522
rect 282954 464614 283574 478000
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 460308 283574 464058
rect 289794 471454 290414 478000
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 460308 290414 470898
rect 293514 475174 294134 478000
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 460308 294134 474618
rect 297234 469138 297854 478000
rect 297234 468902 297266 469138
rect 297502 468902 297586 469138
rect 297822 468902 297854 469138
rect 297234 468818 297854 468902
rect 297234 468582 297266 468818
rect 297502 468582 297586 468818
rect 297822 468582 297854 468818
rect 297234 460308 297854 468582
rect 300954 465554 301574 478000
rect 300954 465318 300986 465554
rect 301222 465318 301306 465554
rect 301542 465318 301574 465554
rect 300954 465234 301574 465318
rect 300954 464998 300986 465234
rect 301222 464998 301306 465234
rect 301542 464998 301574 465234
rect 300954 460308 301574 464998
rect 307794 460308 308414 488898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 460308 312134 492618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 633033 319574 644058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 633033 326414 650898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 633033 330134 654618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 633033 333854 658338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 633033 337574 662058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633033 344414 668898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 633033 348134 636618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 633033 351854 640338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 633033 355574 644058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 633033 362414 650898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 633033 366134 654618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 633033 369854 658338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 633033 373574 662058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633033 380414 668898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 633033 384134 636618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 633033 387854 640338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 633033 391574 644058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 633033 398414 650898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 633033 402134 654618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 633033 405854 658338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 633033 409574 662058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633033 416414 668898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 633033 420134 636618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 633033 423854 640338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 633033 427574 644058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 324208 615454 324528 615486
rect 324208 615218 324250 615454
rect 324486 615218 324528 615454
rect 324208 615134 324528 615218
rect 324208 614898 324250 615134
rect 324486 614898 324528 615134
rect 324208 614866 324528 614898
rect 354928 615454 355248 615486
rect 354928 615218 354970 615454
rect 355206 615218 355248 615454
rect 354928 615134 355248 615218
rect 354928 614898 354970 615134
rect 355206 614898 355248 615134
rect 354928 614866 355248 614898
rect 385648 615454 385968 615486
rect 385648 615218 385690 615454
rect 385926 615218 385968 615454
rect 385648 615134 385968 615218
rect 385648 614898 385690 615134
rect 385926 614898 385968 615134
rect 385648 614866 385968 614898
rect 416368 615454 416688 615486
rect 416368 615218 416410 615454
rect 416646 615218 416688 615454
rect 416368 615134 416688 615218
rect 416368 614898 416410 615134
rect 416646 614898 416688 615134
rect 416368 614866 416688 614898
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 430619 601764 430685 601765
rect 430619 601700 430620 601764
rect 430684 601700 430685 601764
rect 430619 601699 430685 601700
rect 339568 597454 339888 597486
rect 339568 597218 339610 597454
rect 339846 597218 339888 597454
rect 339568 597134 339888 597218
rect 339568 596898 339610 597134
rect 339846 596898 339888 597134
rect 339568 596866 339888 596898
rect 370288 597454 370608 597486
rect 370288 597218 370330 597454
rect 370566 597218 370608 597454
rect 370288 597134 370608 597218
rect 370288 596898 370330 597134
rect 370566 596898 370608 597134
rect 370288 596866 370608 596898
rect 401008 597454 401328 597486
rect 401008 597218 401050 597454
rect 401286 597218 401328 597454
rect 401008 597134 401328 597218
rect 401008 596898 401050 597134
rect 401286 596898 401328 597134
rect 401008 596866 401328 596898
rect 324208 579454 324528 579486
rect 324208 579218 324250 579454
rect 324486 579218 324528 579454
rect 324208 579134 324528 579218
rect 324208 578898 324250 579134
rect 324486 578898 324528 579134
rect 324208 578866 324528 578898
rect 354928 579454 355248 579486
rect 354928 579218 354970 579454
rect 355206 579218 355248 579454
rect 354928 579134 355248 579218
rect 354928 578898 354970 579134
rect 355206 578898 355248 579134
rect 354928 578866 355248 578898
rect 385648 579454 385968 579486
rect 385648 579218 385690 579454
rect 385926 579218 385968 579454
rect 385648 579134 385968 579218
rect 385648 578898 385690 579134
rect 385926 578898 385968 579134
rect 385648 578866 385968 578898
rect 416368 579454 416688 579486
rect 416368 579218 416410 579454
rect 416646 579218 416688 579454
rect 416368 579134 416688 579218
rect 416368 578898 416410 579134
rect 416646 578898 416688 579134
rect 416368 578866 416688 578898
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 339568 561454 339888 561486
rect 339568 561218 339610 561454
rect 339846 561218 339888 561454
rect 339568 561134 339888 561218
rect 339568 560898 339610 561134
rect 339846 560898 339888 561134
rect 339568 560866 339888 560898
rect 370288 561454 370608 561486
rect 370288 561218 370330 561454
rect 370566 561218 370608 561454
rect 370288 561134 370608 561218
rect 370288 560898 370330 561134
rect 370566 560898 370608 561134
rect 370288 560866 370608 560898
rect 401008 561454 401328 561486
rect 401008 561218 401050 561454
rect 401286 561218 401328 561454
rect 401008 561134 401328 561218
rect 401008 560898 401050 561134
rect 401286 560898 401328 561134
rect 401008 560866 401328 560898
rect 324208 543454 324528 543486
rect 324208 543218 324250 543454
rect 324486 543218 324528 543454
rect 324208 543134 324528 543218
rect 324208 542898 324250 543134
rect 324486 542898 324528 543134
rect 324208 542866 324528 542898
rect 354928 543454 355248 543486
rect 354928 543218 354970 543454
rect 355206 543218 355248 543454
rect 354928 543134 355248 543218
rect 354928 542898 354970 543134
rect 355206 542898 355248 543134
rect 354928 542866 355248 542898
rect 385648 543454 385968 543486
rect 385648 543218 385690 543454
rect 385926 543218 385968 543454
rect 385648 543134 385968 543218
rect 385648 542898 385690 543134
rect 385926 542898 385968 543134
rect 385648 542866 385968 542898
rect 416368 543454 416688 543486
rect 416368 543218 416410 543454
rect 416646 543218 416688 543454
rect 416368 543134 416688 543218
rect 416368 542898 416410 543134
rect 416646 542898 416688 543134
rect 416368 542866 416688 542898
rect 320587 541108 320653 541109
rect 320587 541044 320588 541108
rect 320652 541044 320653 541108
rect 320587 541043 320653 541044
rect 320590 538230 320650 541043
rect 320590 538170 320834 538230
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 320774 518669 320834 538170
rect 339568 525454 339888 525486
rect 339568 525218 339610 525454
rect 339846 525218 339888 525454
rect 339568 525134 339888 525218
rect 339568 524898 339610 525134
rect 339846 524898 339888 525134
rect 339568 524866 339888 524898
rect 370288 525454 370608 525486
rect 370288 525218 370330 525454
rect 370566 525218 370608 525454
rect 370288 525134 370608 525218
rect 370288 524898 370330 525134
rect 370566 524898 370608 525134
rect 370288 524866 370608 524898
rect 401008 525454 401328 525486
rect 401008 525218 401050 525454
rect 401286 525218 401328 525454
rect 401008 525134 401328 525218
rect 401008 524898 401050 525134
rect 401286 524898 401328 525134
rect 401008 524866 401328 524898
rect 430622 520165 430682 601699
rect 430803 597684 430869 597685
rect 430803 597620 430804 597684
rect 430868 597620 430869 597684
rect 430803 597619 430869 597620
rect 430619 520164 430685 520165
rect 430619 520100 430620 520164
rect 430684 520100 430685 520164
rect 430619 520099 430685 520100
rect 430806 518805 430866 597619
rect 430987 592244 431053 592245
rect 430987 592180 430988 592244
rect 431052 592180 431053 592244
rect 430987 592179 431053 592180
rect 430803 518804 430869 518805
rect 430803 518740 430804 518804
rect 430868 518740 430869 518804
rect 430803 518739 430869 518740
rect 320771 518668 320837 518669
rect 320771 518604 320772 518668
rect 320836 518604 320837 518668
rect 320771 518603 320837 518604
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460308 315854 496338
rect 318954 500614 319574 518000
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 460308 319574 464058
rect 325794 507454 326414 518000
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 460308 326414 470898
rect 329514 511174 330134 518000
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 460308 330134 474618
rect 333234 514894 333854 518000
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 460308 333854 478338
rect 336954 482614 337574 518000
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 460308 337574 482058
rect 343794 489454 344414 518000
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 338251 461004 338317 461005
rect 338251 460940 338252 461004
rect 338316 460950 338317 461004
rect 339723 461004 339789 461005
rect 338316 460940 338498 460950
rect 338251 460939 338498 460940
rect 339723 460940 339724 461004
rect 339788 460940 339789 461004
rect 339723 460939 339789 460940
rect 338254 460890 338498 460939
rect 338438 458690 338498 460890
rect 339726 458690 339786 460939
rect 343794 460308 344414 488898
rect 347514 493174 348134 518000
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 460308 348134 492618
rect 351234 496894 351854 518000
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 350947 461004 351013 461005
rect 350947 460940 350948 461004
rect 351012 460940 351013 461004
rect 350947 460939 351013 460940
rect 350950 458690 351010 460939
rect 351234 460308 351854 496338
rect 354954 500614 355574 518000
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 361794 507454 362414 518000
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 360883 485076 360949 485077
rect 360883 485012 360884 485076
rect 360948 485012 360949 485076
rect 360883 485011 360949 485012
rect 360699 478820 360765 478821
rect 360699 478756 360700 478820
rect 360764 478756 360765 478820
rect 360699 478755 360765 478756
rect 357939 478004 358005 478005
rect 357939 477940 357940 478004
rect 358004 477940 358005 478004
rect 357939 477939 358005 477940
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 460308 355574 464058
rect 338438 458630 338524 458690
rect 338464 458202 338524 458630
rect 339688 458630 339786 458690
rect 350840 458630 351010 458690
rect 339688 458202 339748 458630
rect 350840 458202 350900 458630
rect 220272 453454 220620 453486
rect 220272 453218 220328 453454
rect 220564 453218 220620 453454
rect 220272 453134 220620 453218
rect 220272 452898 220328 453134
rect 220564 452898 220620 453134
rect 220272 452866 220620 452898
rect 356000 453454 356348 453486
rect 356000 453218 356056 453454
rect 356292 453218 356348 453454
rect 356000 453134 356348 453218
rect 356000 452898 356056 453134
rect 356292 452898 356348 453134
rect 356000 452866 356348 452898
rect 220952 435454 221300 435486
rect 220952 435218 221008 435454
rect 221244 435218 221300 435454
rect 220952 435134 221300 435218
rect 220952 434898 221008 435134
rect 221244 434898 221300 435134
rect 220952 434866 221300 434898
rect 355320 435454 355668 435486
rect 355320 435218 355376 435454
rect 355612 435218 355668 435454
rect 355320 435134 355668 435218
rect 355320 434898 355376 435134
rect 355612 434898 355668 435134
rect 355320 434866 355668 434898
rect 220272 417454 220620 417486
rect 220272 417218 220328 417454
rect 220564 417218 220620 417454
rect 220272 417134 220620 417218
rect 220272 416898 220328 417134
rect 220564 416898 220620 417134
rect 220272 416866 220620 416898
rect 356000 417454 356348 417486
rect 356000 417218 356056 417454
rect 356292 417218 356348 417454
rect 356000 417134 356348 417218
rect 356000 416898 356056 417134
rect 356292 416898 356348 417134
rect 356000 416866 356348 416898
rect 220952 399454 221300 399486
rect 220952 399218 221008 399454
rect 221244 399218 221300 399454
rect 220952 399134 221300 399218
rect 220952 398898 221008 399134
rect 221244 398898 221300 399134
rect 220952 398866 221300 398898
rect 355320 399454 355668 399486
rect 355320 399218 355376 399454
rect 355612 399218 355668 399454
rect 355320 399134 355668 399218
rect 355320 398898 355376 399134
rect 355612 398898 355668 399134
rect 355320 398866 355668 398898
rect 220272 381454 220620 381486
rect 220272 381218 220328 381454
rect 220564 381218 220620 381454
rect 220272 381134 220620 381218
rect 220272 380898 220328 381134
rect 220564 380898 220620 381134
rect 220272 380866 220620 380898
rect 356000 381454 356348 381486
rect 356000 381218 356056 381454
rect 356292 381218 356348 381454
rect 356000 381134 356348 381218
rect 356000 380898 356056 381134
rect 356292 380898 356348 381134
rect 356000 380866 356348 380898
rect 244779 375052 244845 375053
rect 235950 374990 236086 375050
rect 236502 374990 237174 375050
rect 238158 374990 238262 375050
rect 239262 374990 239622 375050
rect 240366 374990 240574 375050
rect 241470 374990 241798 375050
rect 242942 374990 243158 375050
rect 235950 373149 236010 374990
rect 235947 373148 236013 373149
rect 235947 373084 235948 373148
rect 236012 373084 236013 373148
rect 235947 373083 236013 373084
rect 221514 367174 222134 373000
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 355308 222134 366618
rect 225234 370894 225854 373000
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 355308 225854 370338
rect 228954 357554 229574 373000
rect 228954 357318 228986 357554
rect 229222 357318 229306 357554
rect 229542 357318 229574 357554
rect 228954 357234 229574 357318
rect 228954 356998 228986 357234
rect 229222 356998 229306 357234
rect 229542 356998 229574 357234
rect 228954 355308 229574 356998
rect 235794 364394 236414 373000
rect 236502 372605 236562 374990
rect 238158 372605 238218 374990
rect 239262 372605 239322 374990
rect 236499 372604 236565 372605
rect 236499 372540 236500 372604
rect 236564 372540 236565 372604
rect 236499 372539 236565 372540
rect 238155 372604 238221 372605
rect 238155 372540 238156 372604
rect 238220 372540 238221 372604
rect 238155 372539 238221 372540
rect 239259 372604 239325 372605
rect 239259 372540 239260 372604
rect 239324 372540 239325 372604
rect 239259 372539 239325 372540
rect 235794 364158 235826 364394
rect 236062 364158 236146 364394
rect 236382 364158 236414 364394
rect 235794 364074 236414 364158
rect 235794 363838 235826 364074
rect 236062 363838 236146 364074
rect 236382 363838 236414 364074
rect 235794 355308 236414 363838
rect 239514 366234 240134 373000
rect 240366 372605 240426 374990
rect 241470 372605 241530 374990
rect 242942 373285 243002 374990
rect 244230 374509 244290 375050
rect 244779 374988 244780 375052
rect 244844 375050 244845 375052
rect 270539 375052 270605 375053
rect 244844 374990 245470 375050
rect 245886 374990 246558 375050
rect 244844 374988 244845 374990
rect 244779 374987 244845 374988
rect 244227 374508 244293 374509
rect 244227 374444 244228 374508
rect 244292 374444 244293 374508
rect 244227 374443 244293 374444
rect 242939 373284 243005 373285
rect 242939 373220 242940 373284
rect 243004 373220 243005 373284
rect 242939 373219 243005 373220
rect 240363 372604 240429 372605
rect 240363 372540 240364 372604
rect 240428 372540 240429 372604
rect 240363 372539 240429 372540
rect 241467 372604 241533 372605
rect 241467 372540 241468 372604
rect 241532 372540 241533 372604
rect 241467 372539 241533 372540
rect 239514 365998 239546 366234
rect 239782 365998 239866 366234
rect 240102 365998 240134 366234
rect 239514 365914 240134 365998
rect 239514 365678 239546 365914
rect 239782 365678 239866 365914
rect 240102 365678 240134 365914
rect 239514 355308 240134 365678
rect 243234 369954 243854 373000
rect 245886 372605 245946 374990
rect 247616 374509 247676 375020
rect 247910 374990 248326 375050
rect 248462 374990 248734 375050
rect 249934 374990 250094 375050
rect 250302 374990 250774 375050
rect 251222 374990 251318 375050
rect 251958 374990 252406 375050
rect 247613 374508 247679 374509
rect 247613 374444 247614 374508
rect 247678 374444 247679 374508
rect 247613 374443 247679 374444
rect 245883 372604 245949 372605
rect 245883 372540 245884 372604
rect 245948 372540 245949 372604
rect 245883 372539 245949 372540
rect 243234 369718 243266 369954
rect 243502 369718 243586 369954
rect 243822 369718 243854 369954
rect 243234 369634 243854 369718
rect 243234 369398 243266 369634
rect 243502 369398 243586 369634
rect 243822 369398 243854 369634
rect 243234 355308 243854 369398
rect 246954 356614 247574 373000
rect 247910 371653 247970 374990
rect 248462 372605 248522 374990
rect 248459 372604 248525 372605
rect 248459 372540 248460 372604
rect 248524 372540 248525 372604
rect 248459 372539 248525 372540
rect 247907 371652 247973 371653
rect 247907 371588 247908 371652
rect 247972 371588 247973 371652
rect 247907 371587 247973 371588
rect 249934 371381 249994 374990
rect 250302 371653 250362 374990
rect 251222 372605 251282 374990
rect 251219 372604 251285 372605
rect 251219 372540 251220 372604
rect 251284 372540 251285 372604
rect 251219 372539 251285 372540
rect 251958 371653 252018 374990
rect 253464 374509 253524 375020
rect 253461 374508 253527 374509
rect 253461 374444 253462 374508
rect 253526 374444 253527 374508
rect 253461 374443 253527 374444
rect 250299 371652 250365 371653
rect 250299 371588 250300 371652
rect 250364 371588 250365 371652
rect 250299 371587 250365 371588
rect 251955 371652 252021 371653
rect 251955 371588 251956 371652
rect 252020 371588 252021 371652
rect 251955 371587 252021 371588
rect 253614 371381 253674 375050
rect 253982 374990 254582 375050
rect 255454 374990 255942 375050
rect 256078 374990 256250 375050
rect 253982 373149 254042 374990
rect 255454 373149 255514 374990
rect 253979 373148 254045 373149
rect 253979 373084 253980 373148
rect 254044 373084 254045 373148
rect 253979 373083 254045 373084
rect 255451 373148 255517 373149
rect 255451 373084 255452 373148
rect 255516 373084 255517 373148
rect 255451 373083 255517 373084
rect 249931 371380 249997 371381
rect 249931 371316 249932 371380
rect 249996 371316 249997 371380
rect 249931 371315 249997 371316
rect 253611 371380 253677 371381
rect 253611 371316 253612 371380
rect 253676 371316 253677 371380
rect 253611 371315 253677 371316
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 246954 355308 247574 356058
rect 253794 363454 254414 373000
rect 256190 371381 256250 374990
rect 256742 374990 257030 375050
rect 258118 374990 258274 375050
rect 256742 372605 256802 374990
rect 258214 374010 258274 374990
rect 258030 373950 258274 374010
rect 258398 374990 258526 375050
rect 259478 374990 259562 375050
rect 258030 373829 258090 373950
rect 258027 373828 258093 373829
rect 258027 373764 258028 373828
rect 258092 373764 258093 373828
rect 258027 373763 258093 373764
rect 256739 372604 256805 372605
rect 256739 372540 256740 372604
rect 256804 372540 256805 372604
rect 256739 372539 256805 372540
rect 256187 371380 256253 371381
rect 256187 371316 256188 371380
rect 256252 371316 256253 371380
rect 256187 371315 256253 371316
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 355308 254414 362898
rect 257514 367174 258134 373000
rect 258398 371381 258458 374990
rect 259502 372605 259562 374990
rect 260054 374990 260702 375050
rect 260974 374990 261110 375050
rect 261342 374990 261790 375050
rect 262262 374990 262878 375050
rect 260054 372605 260114 374990
rect 259499 372604 259565 372605
rect 259499 372540 259500 372604
rect 259564 372540 259565 372604
rect 259499 372539 259565 372540
rect 260051 372604 260117 372605
rect 260051 372540 260052 372604
rect 260116 372540 260117 372604
rect 260051 372539 260117 372540
rect 260974 371381 261034 374990
rect 261342 373285 261402 374990
rect 262262 374373 262322 374990
rect 262259 374372 262325 374373
rect 262259 374308 262260 374372
rect 262324 374308 262325 374372
rect 262259 374307 262325 374308
rect 261339 373284 261405 373285
rect 261339 373220 261340 373284
rect 261404 373220 261405 373284
rect 261339 373219 261405 373220
rect 258395 371380 258461 371381
rect 258395 371316 258396 371380
rect 258460 371316 258461 371380
rect 258395 371315 258461 371316
rect 260971 371380 261037 371381
rect 260971 371316 260972 371380
rect 261036 371316 261037 371380
rect 260971 371315 261037 371316
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 355308 258134 366618
rect 261234 370894 261854 373000
rect 263550 371381 263610 375050
rect 263734 374990 263966 375050
rect 263734 373557 263794 374990
rect 265296 374509 265356 375020
rect 265758 374990 266006 375050
rect 266310 374990 266414 375050
rect 267046 374990 267638 375050
rect 267782 374990 268318 375050
rect 268518 374990 268726 375050
rect 269254 374990 269814 375050
rect 265293 374508 265359 374509
rect 265293 374444 265294 374508
rect 265358 374444 265359 374508
rect 265293 374443 265359 374444
rect 263731 373556 263797 373557
rect 263731 373492 263732 373556
rect 263796 373492 263797 373556
rect 263731 373491 263797 373492
rect 263547 371380 263613 371381
rect 263547 371316 263548 371380
rect 263612 371316 263613 371380
rect 263547 371315 263613 371316
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 355308 261854 370338
rect 264954 357554 265574 373000
rect 265758 371517 265818 374990
rect 266310 373693 266370 374990
rect 266307 373692 266373 373693
rect 266307 373628 266308 373692
rect 266372 373628 266373 373692
rect 266307 373627 266373 373628
rect 265755 371516 265821 371517
rect 265755 371452 265756 371516
rect 265820 371452 265821 371516
rect 265755 371451 265821 371452
rect 267046 371381 267106 374990
rect 267782 371381 267842 374990
rect 268518 373829 268578 374990
rect 268515 373828 268581 373829
rect 268515 373764 268516 373828
rect 268580 373764 268581 373828
rect 268515 373763 268581 373764
rect 269254 373421 269314 374990
rect 270539 374988 270540 375052
rect 270604 375050 270605 375052
rect 283051 375052 283117 375053
rect 270604 374990 271038 375050
rect 271174 374990 271338 375050
rect 270604 374988 270605 374990
rect 270539 374987 270605 374988
rect 271278 374101 271338 374990
rect 272014 374990 272262 375050
rect 271275 374100 271341 374101
rect 271275 374036 271276 374100
rect 271340 374036 271341 374100
rect 271275 374035 271341 374036
rect 269251 373420 269317 373421
rect 269251 373356 269252 373420
rect 269316 373356 269317 373420
rect 269251 373355 269317 373356
rect 272014 373149 272074 374990
rect 272011 373148 272077 373149
rect 272011 373084 272012 373148
rect 272076 373084 272077 373148
rect 272011 373083 272077 373084
rect 267043 371380 267109 371381
rect 267043 371316 267044 371380
rect 267108 371316 267109 371380
rect 267043 371315 267109 371316
rect 267779 371380 267845 371381
rect 267779 371316 267780 371380
rect 267844 371316 267845 371380
rect 267779 371315 267845 371316
rect 264954 357318 264986 357554
rect 265222 357318 265306 357554
rect 265542 357318 265574 357554
rect 264954 357234 265574 357318
rect 264954 356998 264986 357234
rect 265222 356998 265306 357234
rect 265542 356998 265574 357234
rect 264954 355308 265574 356998
rect 271794 364394 272414 373000
rect 273302 372605 273362 375050
rect 273622 374990 273730 375050
rect 273299 372604 273365 372605
rect 273299 372540 273300 372604
rect 273364 372540 273365 372604
rect 273299 372539 273365 372540
rect 273670 371517 273730 374990
rect 273854 374990 274438 375050
rect 275326 374990 275798 375050
rect 276070 374990 276306 375050
rect 277022 374990 277226 375050
rect 273854 374237 273914 374990
rect 273851 374236 273917 374237
rect 273851 374172 273852 374236
rect 273916 374172 273917 374236
rect 273851 374171 273917 374172
rect 275326 371789 275386 374990
rect 275323 371788 275389 371789
rect 275323 371724 275324 371788
rect 275388 371724 275389 371788
rect 275323 371723 275389 371724
rect 273667 371516 273733 371517
rect 273667 371452 273668 371516
rect 273732 371452 273733 371516
rect 273667 371451 273733 371452
rect 271794 364158 271826 364394
rect 272062 364158 272146 364394
rect 272382 364158 272414 364394
rect 271794 364074 272414 364158
rect 271794 363838 271826 364074
rect 272062 363838 272146 364074
rect 272382 363838 272414 364074
rect 271794 355308 272414 363838
rect 275514 366234 276134 373000
rect 276246 371381 276306 374990
rect 277166 372469 277226 374990
rect 277534 374990 278110 375050
rect 278270 374990 278518 375050
rect 277163 372468 277229 372469
rect 277163 372404 277164 372468
rect 277228 372404 277229 372468
rect 277163 372403 277229 372404
rect 277534 372333 277594 374990
rect 277531 372332 277597 372333
rect 277531 372268 277532 372332
rect 277596 372268 277597 372332
rect 277531 372267 277597 372268
rect 278270 371381 278330 374990
rect 279190 373965 279250 375050
rect 280294 374990 280966 375050
rect 279187 373964 279253 373965
rect 279187 373900 279188 373964
rect 279252 373900 279253 373964
rect 279187 373899 279253 373900
rect 279190 373285 279250 373899
rect 279187 373284 279253 373285
rect 279187 373220 279188 373284
rect 279252 373220 279253 373284
rect 279187 373219 279253 373220
rect 276243 371380 276309 371381
rect 276243 371316 276244 371380
rect 276308 371316 276309 371380
rect 276243 371315 276309 371316
rect 278267 371380 278333 371381
rect 278267 371316 278268 371380
rect 278332 371316 278333 371380
rect 278267 371315 278333 371316
rect 275514 365998 275546 366234
rect 275782 365998 275866 366234
rect 276102 365998 276134 366234
rect 275514 365914 276134 365998
rect 275514 365678 275546 365914
rect 275782 365678 275866 365914
rect 276102 365678 276134 365914
rect 275514 355308 276134 365678
rect 279234 369954 279854 373000
rect 280294 371381 280354 374990
rect 283051 374988 283052 375052
rect 283116 375050 283117 375052
rect 315251 375052 315317 375053
rect 283116 374990 283550 375050
rect 285814 374990 285998 375050
rect 287654 374990 288310 375050
rect 290598 374990 291030 375050
rect 292806 374990 293478 375050
rect 295382 374990 295926 375050
rect 298142 374990 298510 375050
rect 283116 374988 283117 374990
rect 283051 374987 283117 374988
rect 280291 371380 280357 371381
rect 280291 371316 280292 371380
rect 280356 371316 280357 371380
rect 280291 371315 280357 371316
rect 279234 369718 279266 369954
rect 279502 369718 279586 369954
rect 279822 369718 279854 369954
rect 279234 369634 279854 369718
rect 279234 369398 279266 369634
rect 279502 369398 279586 369634
rect 279822 369398 279854 369634
rect 279234 355308 279854 369398
rect 282954 356614 283574 373000
rect 285814 371381 285874 374990
rect 287654 371381 287714 374990
rect 285811 371380 285877 371381
rect 285811 371316 285812 371380
rect 285876 371316 285877 371380
rect 285811 371315 285877 371316
rect 287651 371380 287717 371381
rect 287651 371316 287652 371380
rect 287716 371316 287717 371380
rect 287651 371315 287717 371316
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 355308 283574 356058
rect 289794 363454 290414 373000
rect 290598 371381 290658 374990
rect 292806 371381 292866 374990
rect 290595 371380 290661 371381
rect 290595 371316 290596 371380
rect 290660 371316 290661 371380
rect 290595 371315 290661 371316
rect 292803 371380 292869 371381
rect 292803 371316 292804 371380
rect 292868 371316 292869 371380
rect 292803 371315 292869 371316
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 355308 290414 362898
rect 293514 367174 294134 373000
rect 295382 371381 295442 374990
rect 295379 371380 295445 371381
rect 295379 371316 295380 371380
rect 295444 371316 295445 371380
rect 295379 371315 295445 371316
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 355308 294134 366618
rect 297234 370894 297854 373000
rect 298142 371381 298202 374990
rect 300902 373149 300962 375050
rect 302926 374990 303542 375050
rect 305318 374990 305990 375050
rect 308574 374990 308690 375050
rect 300899 373148 300965 373149
rect 300899 373084 300900 373148
rect 300964 373084 300965 373148
rect 300899 373083 300965 373084
rect 298139 371380 298205 371381
rect 298139 371316 298140 371380
rect 298204 371316 298205 371380
rect 298139 371315 298205 371316
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 355308 297854 370338
rect 300954 357554 301574 373000
rect 302926 371381 302986 374990
rect 305318 372469 305378 374990
rect 305315 372468 305381 372469
rect 305315 372404 305316 372468
rect 305380 372404 305381 372468
rect 305315 372403 305381 372404
rect 302923 371380 302989 371381
rect 302923 371316 302924 371380
rect 302988 371316 302989 371380
rect 302923 371315 302989 371316
rect 300954 357318 300986 357554
rect 301222 357318 301306 357554
rect 301542 357318 301574 357554
rect 300954 357234 301574 357318
rect 300954 356998 300986 357234
rect 301222 356998 301306 357234
rect 301542 356998 301574 357234
rect 300954 355308 301574 356998
rect 307794 364394 308414 373000
rect 308630 371381 308690 374990
rect 310654 374990 311022 375050
rect 310654 372605 310714 374990
rect 310651 372604 310717 372605
rect 310651 372540 310652 372604
rect 310716 372540 310717 372604
rect 310651 372539 310717 372540
rect 308627 371380 308693 371381
rect 308627 371316 308628 371380
rect 308692 371316 308693 371380
rect 308627 371315 308693 371316
rect 307794 364158 307826 364394
rect 308062 364158 308146 364394
rect 308382 364158 308414 364394
rect 307794 364074 308414 364158
rect 307794 363838 307826 364074
rect 308062 363838 308146 364074
rect 308382 363838 308414 364074
rect 307794 355308 308414 363838
rect 311514 366234 312134 373000
rect 313414 372605 313474 375050
rect 315251 374988 315252 375052
rect 315316 375050 315317 375052
rect 315316 374990 315918 375050
rect 317830 374990 318502 375050
rect 315316 374988 315317 374990
rect 315251 374987 315317 374988
rect 313411 372604 313477 372605
rect 313411 372540 313412 372604
rect 313476 372540 313477 372604
rect 313411 372539 313477 372540
rect 311514 365998 311546 366234
rect 311782 365998 311866 366234
rect 312102 365998 312134 366234
rect 311514 365914 312134 365998
rect 311514 365678 311546 365914
rect 311782 365678 311866 365914
rect 312102 365678 312134 365914
rect 311514 355308 312134 365678
rect 315234 369954 315854 373000
rect 317830 371789 317890 374990
rect 320920 374645 320980 375020
rect 322982 374990 323398 375050
rect 325982 374990 326722 375050
rect 320917 374644 320983 374645
rect 320917 374580 320918 374644
rect 320982 374580 320983 374644
rect 320917 374579 320983 374580
rect 317827 371788 317893 371789
rect 317827 371724 317828 371788
rect 317892 371724 317893 371788
rect 317827 371723 317893 371724
rect 315234 369718 315266 369954
rect 315502 369718 315586 369954
rect 315822 369718 315854 369954
rect 315234 369634 315854 369718
rect 315234 369398 315266 369634
rect 315502 369398 315586 369634
rect 315822 369398 315854 369634
rect 315234 355308 315854 369398
rect 318954 356614 319574 373000
rect 322982 371381 323042 374990
rect 322979 371380 323045 371381
rect 322979 371316 322980 371380
rect 323044 371316 323045 371380
rect 322979 371315 323045 371316
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 355308 319574 356058
rect 325794 363454 326414 373000
rect 326662 371653 326722 374990
rect 326659 371652 326725 371653
rect 326659 371588 326660 371652
rect 326724 371588 326725 371652
rect 326659 371587 326725 371588
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 355308 326414 362898
rect 329514 367174 330134 373000
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 355308 330134 366618
rect 333234 370894 333854 373000
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 355308 333854 370338
rect 336954 357554 337574 373000
rect 343222 371381 343282 375050
rect 343390 374990 343466 375050
rect 343406 371381 343466 374990
rect 343219 371380 343285 371381
rect 343219 371316 343220 371380
rect 343284 371316 343285 371380
rect 343219 371315 343285 371316
rect 343403 371380 343469 371381
rect 343403 371316 343404 371380
rect 343468 371316 343469 371380
rect 343403 371315 343469 371316
rect 336954 357318 336986 357554
rect 337222 357318 337306 357554
rect 337542 357318 337574 357554
rect 336954 357234 337574 357318
rect 336954 356998 336986 357234
rect 337222 356998 337306 357234
rect 337542 356998 337574 357234
rect 336954 355308 337574 356998
rect 343794 364394 344414 373000
rect 343794 364158 343826 364394
rect 344062 364158 344146 364394
rect 344382 364158 344414 364394
rect 343794 364074 344414 364158
rect 343794 363838 343826 364074
rect 344062 363838 344146 364074
rect 344382 363838 344414 364074
rect 343794 355308 344414 363838
rect 347514 366234 348134 373000
rect 347514 365998 347546 366234
rect 347782 365998 347866 366234
rect 348102 365998 348134 366234
rect 347514 365914 348134 365998
rect 347514 365678 347546 365914
rect 347782 365678 347866 365914
rect 348102 365678 348134 365914
rect 347514 355308 348134 365678
rect 351234 369954 351854 373000
rect 351234 369718 351266 369954
rect 351502 369718 351586 369954
rect 351822 369718 351854 369954
rect 351234 369634 351854 369718
rect 351234 369398 351266 369634
rect 351502 369398 351586 369634
rect 351822 369398 351854 369634
rect 351234 355308 351854 369398
rect 354954 356614 355574 373000
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 355308 355574 356058
rect 339723 355060 339789 355061
rect 339723 354996 339724 355060
rect 339788 354996 339789 355060
rect 339723 354995 339789 354996
rect 350947 355060 351013 355061
rect 350947 354996 350948 355060
rect 351012 354996 351013 355060
rect 350947 354995 351013 354996
rect 338067 354788 338133 354789
rect 338067 354724 338068 354788
rect 338132 354724 338133 354788
rect 338067 354723 338133 354724
rect 338070 353970 338130 354723
rect 339726 353970 339786 354995
rect 350950 353970 351010 354995
rect 338070 353910 338524 353970
rect 338464 353260 338524 353910
rect 339688 353910 339786 353970
rect 350840 353910 351010 353970
rect 339688 353260 339748 353910
rect 350840 353260 350900 353910
rect 220272 345454 220620 345486
rect 220272 345218 220328 345454
rect 220564 345218 220620 345454
rect 220272 345134 220620 345218
rect 220272 344898 220328 345134
rect 220564 344898 220620 345134
rect 220272 344866 220620 344898
rect 356000 345454 356348 345486
rect 356000 345218 356056 345454
rect 356292 345218 356348 345454
rect 356000 345134 356348 345218
rect 356000 344898 356056 345134
rect 356292 344898 356348 345134
rect 356000 344866 356348 344898
rect 220952 327454 221300 327486
rect 220952 327218 221008 327454
rect 221244 327218 221300 327454
rect 220952 327134 221300 327218
rect 220952 326898 221008 327134
rect 221244 326898 221300 327134
rect 220952 326866 221300 326898
rect 355320 327454 355668 327486
rect 355320 327218 355376 327454
rect 355612 327218 355668 327454
rect 355320 327134 355668 327218
rect 355320 326898 355376 327134
rect 355612 326898 355668 327134
rect 355320 326866 355668 326898
rect 220272 309454 220620 309486
rect 220272 309218 220328 309454
rect 220564 309218 220620 309454
rect 220272 309134 220620 309218
rect 220272 308898 220328 309134
rect 220564 308898 220620 309134
rect 220272 308866 220620 308898
rect 356000 309454 356348 309486
rect 356000 309218 356056 309454
rect 356292 309218 356348 309454
rect 356000 309134 356348 309218
rect 356000 308898 356056 309134
rect 356292 308898 356348 309134
rect 356000 308866 356348 308898
rect 220952 291454 221300 291486
rect 220952 291218 221008 291454
rect 221244 291218 221300 291454
rect 220952 291134 221300 291218
rect 220952 290898 221008 291134
rect 221244 290898 221300 291134
rect 220952 290866 221300 290898
rect 355320 291454 355668 291486
rect 355320 291218 355376 291454
rect 355612 291218 355668 291454
rect 355320 291134 355668 291218
rect 355320 290898 355376 291134
rect 355612 290898 355668 291134
rect 355320 290866 355668 290898
rect 220272 273454 220620 273486
rect 220272 273218 220328 273454
rect 220564 273218 220620 273454
rect 220272 273134 220620 273218
rect 220272 272898 220328 273134
rect 220564 272898 220620 273134
rect 220272 272866 220620 272898
rect 356000 273454 356348 273486
rect 356000 273218 356056 273454
rect 356292 273218 356348 273454
rect 356000 273134 356348 273218
rect 356000 272898 356056 273134
rect 356292 272898 356348 273134
rect 356000 272866 356348 272898
rect 236056 269650 236116 270106
rect 237144 269650 237204 270106
rect 238232 269650 238292 270106
rect 239592 269650 239652 270106
rect 236056 269590 236562 269650
rect 221514 259174 222134 268000
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221514 250308 222134 258618
rect 225234 262894 225854 268000
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 225234 250308 225854 262338
rect 228954 266614 229574 268000
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 228954 250308 229574 266058
rect 235794 256394 236414 268000
rect 236502 267069 236562 269590
rect 237054 269590 237204 269650
rect 238158 269590 238292 269650
rect 239262 269590 239652 269650
rect 240544 269650 240604 270106
rect 241768 269650 241828 270106
rect 243128 269650 243188 270106
rect 240544 269590 240610 269650
rect 236499 267068 236565 267069
rect 236499 267004 236500 267068
rect 236564 267004 236565 267068
rect 236499 267003 236565 267004
rect 237054 266933 237114 269590
rect 237051 266932 237117 266933
rect 237051 266868 237052 266932
rect 237116 266868 237117 266932
rect 237051 266867 237117 266868
rect 238158 265573 238218 269590
rect 239262 265709 239322 269590
rect 239259 265708 239325 265709
rect 239259 265644 239260 265708
rect 239324 265644 239325 265708
rect 239259 265643 239325 265644
rect 238155 265572 238221 265573
rect 238155 265508 238156 265572
rect 238220 265508 238221 265572
rect 238155 265507 238221 265508
rect 235794 256158 235826 256394
rect 236062 256158 236146 256394
rect 236382 256158 236414 256394
rect 235794 256074 236414 256158
rect 235794 255838 235826 256074
rect 236062 255838 236146 256074
rect 236382 255838 236414 256074
rect 235794 250308 236414 255838
rect 239514 260114 240134 268000
rect 240550 266117 240610 269590
rect 241654 269590 241828 269650
rect 243126 269590 243188 269650
rect 244216 269650 244276 270106
rect 245440 269650 245500 270106
rect 246528 269650 246588 270106
rect 244216 269590 244290 269650
rect 240547 266116 240613 266117
rect 240547 266052 240548 266116
rect 240612 266052 240613 266116
rect 240547 266051 240613 266052
rect 241654 265981 241714 269590
rect 243126 268837 243186 269590
rect 243123 268836 243189 268837
rect 243123 268772 243124 268836
rect 243188 268772 243189 268836
rect 243123 268771 243189 268772
rect 241651 265980 241717 265981
rect 241651 265916 241652 265980
rect 241716 265916 241717 265980
rect 241651 265915 241717 265916
rect 239514 259878 239546 260114
rect 239782 259878 239866 260114
rect 240102 259878 240134 260114
rect 239514 259794 240134 259878
rect 239514 259558 239546 259794
rect 239782 259558 239866 259794
rect 240102 259558 240134 259794
rect 239514 250308 240134 259558
rect 243234 261954 243854 268000
rect 244230 266525 244290 269590
rect 245334 269590 245500 269650
rect 246438 269590 246588 269650
rect 247616 269650 247676 270106
rect 248296 269650 248356 270106
rect 248704 269650 248764 270106
rect 247616 269590 247786 269650
rect 244227 266524 244293 266525
rect 244227 266460 244228 266524
rect 244292 266460 244293 266524
rect 244227 266459 244293 266460
rect 245334 266389 245394 269590
rect 246438 266389 246498 269590
rect 245331 266388 245397 266389
rect 245331 266324 245332 266388
rect 245396 266324 245397 266388
rect 245331 266323 245397 266324
rect 246435 266388 246501 266389
rect 246435 266324 246436 266388
rect 246500 266324 246501 266388
rect 246435 266323 246501 266324
rect 243234 261718 243266 261954
rect 243502 261718 243586 261954
rect 243822 261718 243854 261954
rect 243234 261634 243854 261718
rect 243234 261398 243266 261634
rect 243502 261398 243586 261634
rect 243822 261398 243854 261634
rect 243234 250308 243854 261398
rect 246954 265674 247574 268000
rect 247726 266389 247786 269590
rect 248278 269590 248356 269650
rect 248646 269590 248764 269650
rect 250064 269650 250124 270106
rect 250744 269789 250804 270106
rect 250741 269788 250807 269789
rect 250741 269724 250742 269788
rect 250806 269724 250807 269788
rect 250741 269723 250807 269724
rect 251288 269650 251348 270106
rect 252376 269650 252436 270106
rect 253464 269650 253524 270106
rect 250064 269590 250178 269650
rect 248278 266933 248338 269590
rect 248275 266932 248341 266933
rect 248275 266868 248276 266932
rect 248340 266868 248341 266932
rect 248275 266867 248341 266868
rect 248646 266389 248706 269590
rect 250118 266661 250178 269590
rect 251222 269590 251348 269650
rect 252326 269590 252436 269650
rect 253430 269590 253524 269650
rect 253600 269650 253660 270106
rect 254552 269650 254612 270106
rect 255912 269650 255972 270106
rect 253600 269590 253674 269650
rect 250115 266660 250181 266661
rect 250115 266596 250116 266660
rect 250180 266596 250181 266660
rect 250115 266595 250181 266596
rect 251222 266389 251282 269590
rect 252326 266525 252386 269590
rect 252323 266524 252389 266525
rect 252323 266460 252324 266524
rect 252388 266460 252389 266524
rect 252323 266459 252389 266460
rect 253430 266389 253490 269590
rect 253614 266933 253674 269590
rect 254534 269590 254612 269650
rect 255822 269590 255972 269650
rect 256048 269650 256108 270106
rect 257000 269650 257060 270106
rect 258088 269650 258148 270106
rect 258496 269650 258556 270106
rect 256048 269590 256250 269650
rect 253611 266932 253677 266933
rect 253611 266868 253612 266932
rect 253676 266868 253677 266932
rect 253611 266867 253677 266868
rect 247723 266388 247789 266389
rect 247723 266324 247724 266388
rect 247788 266324 247789 266388
rect 247723 266323 247789 266324
rect 248643 266388 248709 266389
rect 248643 266324 248644 266388
rect 248708 266324 248709 266388
rect 248643 266323 248709 266324
rect 251219 266388 251285 266389
rect 251219 266324 251220 266388
rect 251284 266324 251285 266388
rect 251219 266323 251285 266324
rect 253427 266388 253493 266389
rect 253427 266324 253428 266388
rect 253492 266324 253493 266388
rect 253427 266323 253493 266324
rect 246954 265438 246986 265674
rect 247222 265438 247306 265674
rect 247542 265438 247574 265674
rect 246954 265354 247574 265438
rect 246954 265118 246986 265354
rect 247222 265118 247306 265354
rect 247542 265118 247574 265354
rect 246954 250308 247574 265118
rect 253794 255454 254414 268000
rect 254534 266389 254594 269590
rect 255822 267749 255882 269590
rect 255819 267748 255885 267749
rect 255819 267684 255820 267748
rect 255884 267684 255885 267748
rect 255819 267683 255885 267684
rect 256190 267069 256250 269590
rect 256926 269590 257060 269650
rect 257846 269590 258148 269650
rect 258398 269590 258556 269650
rect 259448 269650 259508 270106
rect 260672 269650 260732 270106
rect 261080 269650 261140 270106
rect 261760 269650 261820 270106
rect 262848 269650 262908 270106
rect 259448 269590 259562 269650
rect 256187 267068 256253 267069
rect 256187 267004 256188 267068
rect 256252 267004 256253 267068
rect 256187 267003 256253 267004
rect 256926 266389 256986 269590
rect 257846 268837 257906 269590
rect 257843 268836 257909 268837
rect 257843 268772 257844 268836
rect 257908 268772 257909 268836
rect 257843 268771 257909 268772
rect 254531 266388 254597 266389
rect 254531 266324 254532 266388
rect 254596 266324 254597 266388
rect 254531 266323 254597 266324
rect 256923 266388 256989 266389
rect 256923 266324 256924 266388
rect 256988 266324 256989 266388
rect 256923 266323 256989 266324
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 250308 254414 254898
rect 257514 259174 258134 268000
rect 258398 267749 258458 269590
rect 258395 267748 258461 267749
rect 258395 267684 258396 267748
rect 258460 267684 258461 267748
rect 258395 267683 258461 267684
rect 259502 266389 259562 269590
rect 260606 269590 260732 269650
rect 260974 269590 261140 269650
rect 261710 269590 261820 269650
rect 262814 269590 262908 269650
rect 263528 269650 263588 270106
rect 263936 269650 263996 270106
rect 265296 269650 265356 270106
rect 265976 269650 266036 270106
rect 266384 269650 266444 270106
rect 267608 269650 267668 270106
rect 263528 269590 263610 269650
rect 260606 266525 260666 269590
rect 260974 267749 261034 269590
rect 261710 268837 261770 269590
rect 261707 268836 261773 268837
rect 261707 268772 261708 268836
rect 261772 268772 261773 268836
rect 261707 268771 261773 268772
rect 260971 267748 261037 267749
rect 260971 267684 260972 267748
rect 261036 267684 261037 267748
rect 260971 267683 261037 267684
rect 260603 266524 260669 266525
rect 260603 266460 260604 266524
rect 260668 266460 260669 266524
rect 260603 266459 260669 266460
rect 259499 266388 259565 266389
rect 259499 266324 259500 266388
rect 259564 266324 259565 266388
rect 259499 266323 259565 266324
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 250308 258134 258618
rect 261234 262894 261854 268000
rect 262814 266389 262874 269590
rect 263550 267749 263610 269590
rect 263918 269590 263996 269650
rect 265206 269590 265356 269650
rect 265942 269590 266036 269650
rect 266310 269590 266444 269650
rect 267598 269590 267668 269650
rect 268288 269650 268348 270106
rect 268696 269650 268756 270106
rect 269784 269650 269844 270106
rect 271008 269650 271068 270106
rect 268288 269590 268394 269650
rect 268696 269590 268762 269650
rect 269784 269590 269866 269650
rect 263547 267748 263613 267749
rect 263547 267684 263548 267748
rect 263612 267684 263613 267748
rect 263547 267683 263613 267684
rect 263918 266389 263978 269590
rect 265206 268157 265266 269590
rect 265203 268156 265269 268157
rect 265203 268092 265204 268156
rect 265268 268092 265269 268156
rect 265203 268091 265269 268092
rect 264954 266614 265574 268000
rect 265942 267749 266002 269590
rect 265939 267748 266005 267749
rect 265939 267684 265940 267748
rect 266004 267684 266005 267748
rect 265939 267683 266005 267684
rect 262811 266388 262877 266389
rect 262811 266324 262812 266388
rect 262876 266324 262877 266388
rect 262811 266323 262877 266324
rect 263915 266388 263981 266389
rect 263915 266324 263916 266388
rect 263980 266324 263981 266388
rect 263915 266323 263981 266324
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 266310 266389 266370 269590
rect 267598 266525 267658 269590
rect 268334 267749 268394 269590
rect 268331 267748 268397 267749
rect 268331 267684 268332 267748
rect 268396 267684 268397 267748
rect 268331 267683 268397 267684
rect 267595 266524 267661 266525
rect 267595 266460 267596 266524
rect 267660 266460 267661 266524
rect 267595 266459 267661 266460
rect 268702 266389 268762 269590
rect 269806 266389 269866 269590
rect 270910 269590 271068 269650
rect 271144 269650 271204 270106
rect 272232 269650 272292 270106
rect 273320 269650 273380 270106
rect 273592 269650 273652 270106
rect 274408 269650 274468 270106
rect 271144 269590 271338 269650
rect 272232 269590 272626 269650
rect 270910 267749 270970 269590
rect 270907 267748 270973 267749
rect 270907 267684 270908 267748
rect 270972 267684 270973 267748
rect 270907 267683 270973 267684
rect 271278 266389 271338 269590
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 250308 261854 262338
rect 264954 266294 265574 266378
rect 266307 266388 266373 266389
rect 266307 266324 266308 266388
rect 266372 266324 266373 266388
rect 266307 266323 266373 266324
rect 268699 266388 268765 266389
rect 268699 266324 268700 266388
rect 268764 266324 268765 266388
rect 268699 266323 268765 266324
rect 269803 266388 269869 266389
rect 269803 266324 269804 266388
rect 269868 266324 269869 266388
rect 269803 266323 269869 266324
rect 271275 266388 271341 266389
rect 271275 266324 271276 266388
rect 271340 266324 271341 266388
rect 271275 266323 271341 266324
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 250308 265574 266058
rect 271794 256394 272414 268000
rect 272566 266253 272626 269590
rect 273302 269590 273380 269650
rect 273486 269590 273652 269650
rect 274406 269590 274468 269650
rect 275768 269650 275828 270106
rect 276040 269650 276100 270106
rect 276992 269650 277052 270106
rect 275768 269590 275938 269650
rect 276040 269590 276306 269650
rect 273302 267069 273362 269590
rect 273486 267749 273546 269590
rect 273483 267748 273549 267749
rect 273483 267684 273484 267748
rect 273548 267684 273549 267748
rect 273483 267683 273549 267684
rect 273299 267068 273365 267069
rect 273299 267004 273300 267068
rect 273364 267004 273365 267068
rect 273299 267003 273365 267004
rect 274406 266389 274466 269590
rect 275878 268157 275938 269590
rect 275875 268156 275941 268157
rect 275875 268092 275876 268156
rect 275940 268092 275941 268156
rect 275875 268091 275941 268092
rect 274403 266388 274469 266389
rect 274403 266324 274404 266388
rect 274468 266324 274469 266388
rect 274403 266323 274469 266324
rect 272563 266252 272629 266253
rect 272563 266188 272564 266252
rect 272628 266188 272629 266252
rect 272563 266187 272629 266188
rect 271794 256158 271826 256394
rect 272062 256158 272146 256394
rect 272382 256158 272414 256394
rect 271794 256074 272414 256158
rect 271794 255838 271826 256074
rect 272062 255838 272146 256074
rect 272382 255838 272414 256074
rect 271794 250308 272414 255838
rect 275514 260114 276134 268000
rect 276246 267749 276306 269590
rect 276982 269590 277052 269650
rect 278080 269650 278140 270106
rect 278488 269650 278548 270106
rect 279168 269650 279228 270106
rect 280936 269650 280996 270106
rect 283520 269653 283580 270106
rect 278080 269590 278146 269650
rect 276982 267749 277042 269590
rect 278086 267749 278146 269590
rect 278454 269590 278548 269650
rect 279006 269590 279228 269650
rect 280846 269590 280996 269650
rect 283517 269652 283583 269653
rect 276243 267748 276309 267749
rect 276243 267684 276244 267748
rect 276308 267684 276309 267748
rect 276243 267683 276309 267684
rect 276979 267748 277045 267749
rect 276979 267684 276980 267748
rect 277044 267684 277045 267748
rect 276979 267683 277045 267684
rect 278083 267748 278149 267749
rect 278083 267684 278084 267748
rect 278148 267684 278149 267748
rect 278083 267683 278149 267684
rect 278454 267205 278514 269590
rect 279006 267205 279066 269590
rect 278451 267204 278517 267205
rect 278451 267140 278452 267204
rect 278516 267140 278517 267204
rect 278451 267139 278517 267140
rect 279003 267204 279069 267205
rect 279003 267140 279004 267204
rect 279068 267140 279069 267204
rect 279003 267139 279069 267140
rect 275514 259878 275546 260114
rect 275782 259878 275866 260114
rect 276102 259878 276134 260114
rect 275514 259794 276134 259878
rect 275514 259558 275546 259794
rect 275782 259558 275866 259794
rect 276102 259558 276134 259794
rect 275514 250308 276134 259558
rect 279234 261954 279854 268000
rect 280846 267749 280906 269590
rect 283517 269588 283518 269652
rect 283582 269588 283583 269652
rect 285968 269650 286028 270106
rect 288280 269653 288340 270106
rect 291000 269653 291060 270106
rect 293448 269653 293508 270106
rect 288277 269652 288343 269653
rect 285968 269590 286058 269650
rect 283517 269587 283583 269588
rect 280843 267748 280909 267749
rect 280843 267684 280844 267748
rect 280908 267684 280909 267748
rect 280843 267683 280909 267684
rect 279234 261718 279266 261954
rect 279502 261718 279586 261954
rect 279822 261718 279854 261954
rect 279234 261634 279854 261718
rect 279234 261398 279266 261634
rect 279502 261398 279586 261634
rect 279822 261398 279854 261634
rect 279234 250308 279854 261398
rect 282954 265674 283574 268000
rect 285998 266933 286058 269590
rect 288277 269588 288278 269652
rect 288342 269588 288343 269652
rect 288277 269587 288343 269588
rect 290997 269652 291063 269653
rect 290997 269588 290998 269652
rect 291062 269588 291063 269652
rect 290997 269587 291063 269588
rect 293445 269652 293511 269653
rect 293445 269588 293446 269652
rect 293510 269588 293511 269652
rect 295896 269650 295956 270106
rect 298480 269650 298540 270106
rect 300928 269650 300988 270106
rect 303512 269650 303572 270106
rect 305960 269653 306020 270106
rect 295896 269590 295994 269650
rect 298480 269590 298570 269650
rect 293445 269587 293511 269588
rect 295934 268837 295994 269590
rect 298510 268837 298570 269590
rect 300902 269590 300988 269650
rect 303478 269590 303572 269650
rect 305957 269652 306023 269653
rect 300902 268837 300962 269590
rect 303478 268837 303538 269590
rect 305957 269588 305958 269652
rect 306022 269588 306023 269652
rect 308544 269650 308604 270106
rect 310992 269650 311052 270106
rect 313440 269650 313500 270106
rect 315888 269650 315948 270106
rect 318472 269653 318532 270106
rect 308544 269590 308690 269650
rect 310992 269590 311082 269650
rect 305957 269587 306023 269588
rect 295931 268836 295997 268837
rect 295931 268772 295932 268836
rect 295996 268772 295997 268836
rect 295931 268771 295997 268772
rect 298507 268836 298573 268837
rect 298507 268772 298508 268836
rect 298572 268772 298573 268836
rect 298507 268771 298573 268772
rect 300899 268836 300965 268837
rect 300899 268772 300900 268836
rect 300964 268772 300965 268836
rect 300899 268771 300965 268772
rect 303475 268836 303541 268837
rect 303475 268772 303476 268836
rect 303540 268772 303541 268836
rect 303475 268771 303541 268772
rect 285995 266932 286061 266933
rect 285995 266868 285996 266932
rect 286060 266868 286061 266932
rect 285995 266867 286061 266868
rect 282954 265438 282986 265674
rect 283222 265438 283306 265674
rect 283542 265438 283574 265674
rect 282954 265354 283574 265438
rect 282954 265118 282986 265354
rect 283222 265118 283306 265354
rect 283542 265118 283574 265354
rect 282954 250308 283574 265118
rect 289794 255454 290414 268000
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 250308 290414 254898
rect 293514 259174 294134 268000
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 250308 294134 258618
rect 297234 262894 297854 268000
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 250308 297854 262338
rect 300954 266614 301574 268000
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 250308 301574 266058
rect 307794 256394 308414 268000
rect 308630 267341 308690 269590
rect 311022 269109 311082 269590
rect 313414 269590 313500 269650
rect 315806 269590 315948 269650
rect 318469 269652 318535 269653
rect 311019 269108 311085 269109
rect 311019 269044 311020 269108
rect 311084 269044 311085 269108
rect 311019 269043 311085 269044
rect 308627 267340 308693 267341
rect 308627 267276 308628 267340
rect 308692 267276 308693 267340
rect 308627 267275 308693 267276
rect 307794 256158 307826 256394
rect 308062 256158 308146 256394
rect 308382 256158 308414 256394
rect 307794 256074 308414 256158
rect 307794 255838 307826 256074
rect 308062 255838 308146 256074
rect 308382 255838 308414 256074
rect 307794 250308 308414 255838
rect 311514 260114 312134 268000
rect 313414 267477 313474 269590
rect 315806 268290 315866 269590
rect 318469 269588 318470 269652
rect 318534 269588 318535 269652
rect 320920 269650 320980 270106
rect 323368 269650 323428 270106
rect 320920 269590 321018 269650
rect 318469 269587 318535 269588
rect 320958 268973 321018 269590
rect 323350 269590 323428 269650
rect 325952 269650 326012 270106
rect 343224 269650 343284 270106
rect 325952 269590 326722 269650
rect 323350 269109 323410 269590
rect 323347 269108 323413 269109
rect 323347 269044 323348 269108
rect 323412 269044 323413 269108
rect 323347 269043 323413 269044
rect 320955 268972 321021 268973
rect 320955 268908 320956 268972
rect 321020 268908 321021 268972
rect 320955 268907 321021 268908
rect 315806 268230 316050 268290
rect 313411 267476 313477 267477
rect 313411 267412 313412 267476
rect 313476 267412 313477 267476
rect 313411 267411 313477 267412
rect 311514 259878 311546 260114
rect 311782 259878 311866 260114
rect 312102 259878 312134 260114
rect 311514 259794 312134 259878
rect 311514 259558 311546 259794
rect 311782 259558 311866 259794
rect 312102 259558 312134 259794
rect 311514 250308 312134 259558
rect 315234 261954 315854 268000
rect 315990 267613 316050 268230
rect 315987 267612 316053 267613
rect 315987 267548 315988 267612
rect 316052 267548 316053 267612
rect 315987 267547 316053 267548
rect 315234 261718 315266 261954
rect 315502 261718 315586 261954
rect 315822 261718 315854 261954
rect 315234 261634 315854 261718
rect 315234 261398 315266 261634
rect 315502 261398 315586 261634
rect 315822 261398 315854 261634
rect 315234 250308 315854 261398
rect 318954 265674 319574 268000
rect 318954 265438 318986 265674
rect 319222 265438 319306 265674
rect 319542 265438 319574 265674
rect 318954 265354 319574 265438
rect 318954 265118 318986 265354
rect 319222 265118 319306 265354
rect 319542 265118 319574 265354
rect 318954 250308 319574 265118
rect 325794 255454 326414 268000
rect 326662 266797 326722 269590
rect 343222 269590 343284 269650
rect 343360 269650 343420 270106
rect 343360 269590 343466 269650
rect 326659 266796 326725 266797
rect 326659 266732 326660 266796
rect 326724 266732 326725 266796
rect 326659 266731 326725 266732
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 250308 326414 254898
rect 329514 259174 330134 268000
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 250308 330134 258618
rect 333234 262894 333854 268000
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 250308 333854 262338
rect 336954 266614 337574 268000
rect 343222 267477 343282 269590
rect 343219 267476 343285 267477
rect 343219 267412 343220 267476
rect 343284 267412 343285 267476
rect 343219 267411 343285 267412
rect 343406 267069 343466 269590
rect 343403 267068 343469 267069
rect 343403 267004 343404 267068
rect 343468 267004 343469 267068
rect 343403 267003 343469 267004
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 250308 337574 266058
rect 343794 256394 344414 268000
rect 343794 256158 343826 256394
rect 344062 256158 344146 256394
rect 344382 256158 344414 256394
rect 343794 256074 344414 256158
rect 343794 255838 343826 256074
rect 344062 255838 344146 256074
rect 344382 255838 344414 256074
rect 343794 250308 344414 255838
rect 347514 260114 348134 268000
rect 347514 259878 347546 260114
rect 347782 259878 347866 260114
rect 348102 259878 348134 260114
rect 347514 259794 348134 259878
rect 347514 259558 347546 259794
rect 347782 259558 347866 259794
rect 348102 259558 348134 259794
rect 347514 250308 348134 259558
rect 351234 261954 351854 268000
rect 351234 261718 351266 261954
rect 351502 261718 351586 261954
rect 351822 261718 351854 261954
rect 351234 261634 351854 261718
rect 351234 261398 351266 261634
rect 351502 261398 351586 261634
rect 351822 261398 351854 261634
rect 351234 250308 351854 261398
rect 354954 265674 355574 268000
rect 354954 265438 354986 265674
rect 355222 265438 355306 265674
rect 355542 265438 355574 265674
rect 354954 265354 355574 265438
rect 354954 265118 354986 265354
rect 355222 265118 355306 265354
rect 355542 265118 355574 265354
rect 354954 250308 355574 265118
rect 338435 249932 338501 249933
rect 338435 249868 338436 249932
rect 338500 249868 338501 249932
rect 338435 249867 338501 249868
rect 339723 249932 339789 249933
rect 339723 249868 339724 249932
rect 339788 249868 339789 249932
rect 339723 249867 339789 249868
rect 350947 249932 351013 249933
rect 350947 249868 350948 249932
rect 351012 249868 351013 249932
rect 350947 249867 351013 249868
rect 338438 248430 338498 249867
rect 339726 248430 339786 249867
rect 350950 248430 351010 249867
rect 338438 248370 338524 248430
rect 338464 248202 338524 248370
rect 339688 248370 339786 248430
rect 350840 248370 351010 248430
rect 339688 248202 339748 248370
rect 350840 248202 350900 248370
rect 220272 237454 220620 237486
rect 220272 237218 220328 237454
rect 220564 237218 220620 237454
rect 220272 237134 220620 237218
rect 220272 236898 220328 237134
rect 220564 236898 220620 237134
rect 220272 236866 220620 236898
rect 356000 237454 356348 237486
rect 356000 237218 356056 237454
rect 356292 237218 356348 237454
rect 356000 237134 356348 237218
rect 356000 236898 356056 237134
rect 356292 236898 356348 237134
rect 356000 236866 356348 236898
rect 220952 219454 221300 219486
rect 220952 219218 221008 219454
rect 221244 219218 221300 219454
rect 220952 219134 221300 219218
rect 220952 218898 221008 219134
rect 221244 218898 221300 219134
rect 220952 218866 221300 218898
rect 355320 219454 355668 219486
rect 355320 219218 355376 219454
rect 355612 219218 355668 219454
rect 355320 219134 355668 219218
rect 355320 218898 355376 219134
rect 355612 218898 355668 219134
rect 355320 218866 355668 218898
rect 220272 201454 220620 201486
rect 220272 201218 220328 201454
rect 220564 201218 220620 201454
rect 220272 201134 220620 201218
rect 220272 200898 220328 201134
rect 220564 200898 220620 201134
rect 220272 200866 220620 200898
rect 356000 201454 356348 201486
rect 356000 201218 356056 201454
rect 356292 201218 356348 201454
rect 356000 201134 356348 201218
rect 356000 200898 356056 201134
rect 356292 200898 356348 201134
rect 356000 200866 356348 200898
rect 220952 183454 221300 183486
rect 220952 183218 221008 183454
rect 221244 183218 221300 183454
rect 220952 183134 221300 183218
rect 220952 182898 221008 183134
rect 221244 182898 221300 183134
rect 220952 182866 221300 182898
rect 355320 183454 355668 183486
rect 355320 183218 355376 183454
rect 355612 183218 355668 183454
rect 355320 183134 355668 183218
rect 355320 182898 355376 183134
rect 355612 182898 355668 183134
rect 355320 182866 355668 182898
rect 236056 164930 236116 165106
rect 237144 164930 237204 165106
rect 238232 164930 238292 165106
rect 239592 164930 239652 165106
rect 235950 164870 236116 164930
rect 237054 164870 237204 164930
rect 238158 164870 238292 164930
rect 239446 164870 239652 164930
rect 240544 164930 240604 165106
rect 241768 164930 241828 165106
rect 243128 164930 243188 165106
rect 240544 164870 240610 164930
rect 235950 163165 236010 164870
rect 235947 163164 236013 163165
rect 235947 163100 235948 163164
rect 236012 163100 236013 163164
rect 235947 163099 236013 163100
rect 221514 151174 222134 163000
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 145308 222134 150618
rect 225234 154894 225854 163000
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 225234 145308 225854 154338
rect 228954 158614 229574 163000
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228954 145308 229574 158058
rect 235794 148394 236414 163000
rect 237054 162757 237114 164870
rect 238158 162757 238218 164870
rect 239446 164250 239506 164870
rect 238526 164190 239506 164250
rect 237051 162756 237117 162757
rect 237051 162692 237052 162756
rect 237116 162692 237117 162756
rect 237051 162691 237117 162692
rect 238155 162756 238221 162757
rect 238155 162692 238156 162756
rect 238220 162692 238221 162756
rect 238155 162691 238221 162692
rect 238526 161530 238586 164190
rect 238707 161532 238773 161533
rect 238707 161530 238708 161532
rect 238526 161470 238708 161530
rect 238707 161468 238708 161470
rect 238772 161468 238773 161532
rect 238707 161467 238773 161468
rect 235794 148158 235826 148394
rect 236062 148158 236146 148394
rect 236382 148158 236414 148394
rect 235794 148074 236414 148158
rect 235794 147838 235826 148074
rect 236062 147838 236146 148074
rect 236382 147838 236414 148074
rect 235794 145308 236414 147838
rect 239514 152114 240134 163000
rect 240550 162757 240610 164870
rect 241654 164870 241828 164930
rect 242942 164870 243188 164930
rect 244216 164930 244276 165106
rect 245440 164930 245500 165106
rect 246528 164930 246588 165106
rect 244216 164870 244290 164930
rect 241654 162757 241714 164870
rect 242942 162757 243002 164870
rect 240547 162756 240613 162757
rect 240547 162692 240548 162756
rect 240612 162692 240613 162756
rect 240547 162691 240613 162692
rect 241651 162756 241717 162757
rect 241651 162692 241652 162756
rect 241716 162692 241717 162756
rect 241651 162691 241717 162692
rect 242939 162756 243005 162757
rect 242939 162692 242940 162756
rect 243004 162692 243005 162756
rect 242939 162691 243005 162692
rect 239514 151878 239546 152114
rect 239782 151878 239866 152114
rect 240102 151878 240134 152114
rect 239514 151794 240134 151878
rect 239514 151558 239546 151794
rect 239782 151558 239866 151794
rect 240102 151558 240134 151794
rect 239514 145308 240134 151558
rect 243234 153954 243854 163000
rect 244230 162757 244290 164870
rect 245334 164870 245500 164930
rect 246438 164870 246588 164930
rect 247616 164930 247676 165106
rect 248296 164930 248356 165106
rect 248704 164930 248764 165106
rect 247616 164870 247786 164930
rect 244227 162756 244293 162757
rect 244227 162692 244228 162756
rect 244292 162692 244293 162756
rect 244227 162691 244293 162692
rect 245334 162077 245394 164870
rect 246438 162757 246498 164870
rect 246435 162756 246501 162757
rect 246435 162692 246436 162756
rect 246500 162692 246501 162756
rect 246435 162691 246501 162692
rect 245331 162076 245397 162077
rect 245331 162012 245332 162076
rect 245396 162012 245397 162076
rect 245331 162011 245397 162012
rect 243234 153718 243266 153954
rect 243502 153718 243586 153954
rect 243822 153718 243854 153954
rect 243234 153634 243854 153718
rect 243234 153398 243266 153634
rect 243502 153398 243586 153634
rect 243822 153398 243854 153634
rect 243234 145308 243854 153398
rect 246954 157674 247574 163000
rect 247726 162757 247786 164870
rect 248278 164870 248356 164930
rect 248646 164870 248764 164930
rect 250064 164930 250124 165106
rect 250744 164930 250804 165106
rect 251288 164930 251348 165106
rect 252376 164930 252436 165106
rect 253464 164930 253524 165106
rect 250064 164870 250178 164930
rect 248278 162757 248338 164870
rect 248646 162757 248706 164870
rect 250118 162757 250178 164870
rect 250670 164870 250804 164930
rect 251222 164870 251348 164930
rect 252326 164870 252436 164930
rect 253430 164870 253524 164930
rect 253600 164930 253660 165106
rect 254552 164930 254612 165106
rect 255912 164930 255972 165106
rect 253600 164870 253674 164930
rect 250670 162757 250730 164870
rect 251222 162757 251282 164870
rect 247723 162756 247789 162757
rect 247723 162692 247724 162756
rect 247788 162692 247789 162756
rect 247723 162691 247789 162692
rect 248275 162756 248341 162757
rect 248275 162692 248276 162756
rect 248340 162692 248341 162756
rect 248275 162691 248341 162692
rect 248643 162756 248709 162757
rect 248643 162692 248644 162756
rect 248708 162692 248709 162756
rect 248643 162691 248709 162692
rect 250115 162756 250181 162757
rect 250115 162692 250116 162756
rect 250180 162692 250181 162756
rect 250115 162691 250181 162692
rect 250667 162756 250733 162757
rect 250667 162692 250668 162756
rect 250732 162692 250733 162756
rect 250667 162691 250733 162692
rect 251219 162756 251285 162757
rect 251219 162692 251220 162756
rect 251284 162692 251285 162756
rect 251219 162691 251285 162692
rect 252326 162077 252386 164870
rect 253430 162757 253490 164870
rect 253614 162757 253674 164870
rect 254534 164870 254612 164930
rect 255822 164870 255972 164930
rect 256048 164930 256108 165106
rect 257000 164930 257060 165106
rect 256048 164870 256250 164930
rect 253427 162756 253493 162757
rect 253427 162692 253428 162756
rect 253492 162692 253493 162756
rect 253427 162691 253493 162692
rect 253611 162756 253677 162757
rect 253611 162692 253612 162756
rect 253676 162692 253677 162756
rect 253611 162691 253677 162692
rect 252323 162076 252389 162077
rect 252323 162012 252324 162076
rect 252388 162012 252389 162076
rect 252323 162011 252389 162012
rect 246954 157438 246986 157674
rect 247222 157438 247306 157674
rect 247542 157438 247574 157674
rect 246954 157354 247574 157438
rect 246954 157118 246986 157354
rect 247222 157118 247306 157354
rect 247542 157118 247574 157354
rect 246954 145308 247574 157118
rect 253794 147454 254414 163000
rect 254534 162757 254594 164870
rect 255822 162757 255882 164870
rect 256190 162757 256250 164870
rect 256926 164870 257060 164930
rect 258088 164930 258148 165106
rect 258496 164930 258556 165106
rect 258088 164870 258274 164930
rect 256926 162757 256986 164870
rect 254531 162756 254597 162757
rect 254531 162692 254532 162756
rect 254596 162692 254597 162756
rect 254531 162691 254597 162692
rect 255819 162756 255885 162757
rect 255819 162692 255820 162756
rect 255884 162692 255885 162756
rect 255819 162691 255885 162692
rect 256187 162756 256253 162757
rect 256187 162692 256188 162756
rect 256252 162692 256253 162756
rect 256187 162691 256253 162692
rect 256923 162756 256989 162757
rect 256923 162692 256924 162756
rect 256988 162692 256989 162756
rect 256923 162691 256989 162692
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 145308 254414 146898
rect 257514 151174 258134 163000
rect 258214 161530 258274 164870
rect 258398 164870 258556 164930
rect 259448 164930 259508 165106
rect 260672 164930 260732 165106
rect 259448 164870 259562 164930
rect 258398 162757 258458 164870
rect 259502 162757 259562 164870
rect 260606 164870 260732 164930
rect 258395 162756 258461 162757
rect 258395 162692 258396 162756
rect 258460 162692 258461 162756
rect 258395 162691 258461 162692
rect 259499 162756 259565 162757
rect 259499 162692 259500 162756
rect 259564 162692 259565 162756
rect 259499 162691 259565 162692
rect 260606 162077 260666 164870
rect 261080 164797 261140 165106
rect 261760 164930 261820 165106
rect 262848 164930 262908 165106
rect 261710 164870 261820 164930
rect 262814 164870 262908 164930
rect 263528 164930 263588 165106
rect 263936 164930 263996 165106
rect 265296 164930 265356 165106
rect 265976 164930 266036 165106
rect 266384 164930 266444 165106
rect 267608 164930 267668 165106
rect 263528 164870 263610 164930
rect 261077 164796 261143 164797
rect 261077 164732 261078 164796
rect 261142 164732 261143 164796
rect 261077 164731 261143 164732
rect 261710 163165 261770 164870
rect 261707 163164 261773 163165
rect 261707 163100 261708 163164
rect 261772 163100 261773 163164
rect 261707 163099 261773 163100
rect 260603 162076 260669 162077
rect 260603 162012 260604 162076
rect 260668 162012 260669 162076
rect 260603 162011 260669 162012
rect 258395 161532 258461 161533
rect 258395 161530 258396 161532
rect 258214 161470 258396 161530
rect 258395 161468 258396 161470
rect 258460 161468 258461 161532
rect 258395 161467 258461 161468
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 145308 258134 150618
rect 261234 154894 261854 163000
rect 262814 162757 262874 164870
rect 263550 162893 263610 164870
rect 263918 164870 263996 164930
rect 265206 164870 265356 164930
rect 265942 164870 266036 164930
rect 266310 164870 266444 164930
rect 267598 164870 267668 164930
rect 263547 162892 263613 162893
rect 263547 162828 263548 162892
rect 263612 162828 263613 162892
rect 263547 162827 263613 162828
rect 263918 162757 263978 164870
rect 265206 163165 265266 164870
rect 265942 164525 266002 164870
rect 265939 164524 266005 164525
rect 265939 164460 265940 164524
rect 266004 164460 266005 164524
rect 265939 164459 266005 164460
rect 265203 163164 265269 163165
rect 265203 163100 265204 163164
rect 265268 163100 265269 163164
rect 265203 163099 265269 163100
rect 262811 162756 262877 162757
rect 262811 162692 262812 162756
rect 262876 162692 262877 162756
rect 262811 162691 262877 162692
rect 263915 162756 263981 162757
rect 263915 162692 263916 162756
rect 263980 162692 263981 162756
rect 263915 162691 263981 162692
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 145308 261854 154338
rect 264954 158614 265574 163000
rect 266310 162757 266370 164870
rect 267598 162757 267658 164870
rect 268288 164658 268348 165106
rect 268696 164658 268756 165106
rect 269784 164658 269844 165106
rect 271008 164930 271068 165106
rect 270910 164870 271068 164930
rect 268288 164598 268394 164658
rect 268696 164598 268762 164658
rect 269784 164598 269866 164658
rect 268334 162893 268394 164598
rect 268331 162892 268397 162893
rect 268331 162828 268332 162892
rect 268396 162828 268397 162892
rect 268331 162827 268397 162828
rect 268702 162757 268762 164598
rect 269806 162757 269866 164598
rect 270910 163845 270970 164870
rect 271144 164658 271204 165106
rect 272232 164658 272292 165106
rect 273320 164658 273380 165106
rect 273592 164930 273652 165106
rect 271094 164598 271204 164658
rect 272198 164598 272292 164658
rect 273302 164598 273380 164658
rect 273486 164870 273652 164930
rect 270907 163844 270973 163845
rect 270907 163780 270908 163844
rect 270972 163780 270973 163844
rect 270907 163779 270973 163780
rect 271094 162757 271154 164598
rect 272198 163165 272258 164598
rect 272195 163164 272261 163165
rect 272195 163100 272196 163164
rect 272260 163100 272261 163164
rect 272195 163099 272261 163100
rect 266307 162756 266373 162757
rect 266307 162692 266308 162756
rect 266372 162692 266373 162756
rect 266307 162691 266373 162692
rect 267595 162756 267661 162757
rect 267595 162692 267596 162756
rect 267660 162692 267661 162756
rect 267595 162691 267661 162692
rect 268699 162756 268765 162757
rect 268699 162692 268700 162756
rect 268764 162692 268765 162756
rect 268699 162691 268765 162692
rect 269803 162756 269869 162757
rect 269803 162692 269804 162756
rect 269868 162692 269869 162756
rect 269803 162691 269869 162692
rect 271091 162756 271157 162757
rect 271091 162692 271092 162756
rect 271156 162692 271157 162756
rect 271091 162691 271157 162692
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 145308 265574 158058
rect 271794 148394 272414 163000
rect 273302 162077 273362 164598
rect 273486 162893 273546 164870
rect 274408 164658 274468 165106
rect 275768 164658 275828 165106
rect 274406 164598 274468 164658
rect 275326 164598 275828 164658
rect 276040 164658 276100 165106
rect 276992 164658 277052 165106
rect 278080 164930 278140 165106
rect 276040 164598 276122 164658
rect 273483 162892 273549 162893
rect 273483 162828 273484 162892
rect 273548 162828 273549 162892
rect 273483 162827 273549 162828
rect 274406 162757 274466 164598
rect 275326 162757 275386 164598
rect 276062 163165 276122 164598
rect 276982 164598 277052 164658
rect 277166 164870 278140 164930
rect 276059 163164 276125 163165
rect 276059 163100 276060 163164
rect 276124 163100 276125 163164
rect 276059 163099 276125 163100
rect 274403 162756 274469 162757
rect 274403 162692 274404 162756
rect 274468 162692 274469 162756
rect 274403 162691 274469 162692
rect 275323 162756 275389 162757
rect 275323 162692 275324 162756
rect 275388 162692 275389 162756
rect 275323 162691 275389 162692
rect 273299 162076 273365 162077
rect 273299 162012 273300 162076
rect 273364 162012 273365 162076
rect 273299 162011 273365 162012
rect 271794 148158 271826 148394
rect 272062 148158 272146 148394
rect 272382 148158 272414 148394
rect 271794 148074 272414 148158
rect 271794 147838 271826 148074
rect 272062 147838 272146 148074
rect 272382 147838 272414 148074
rect 271794 145308 272414 147838
rect 275514 152114 276134 163000
rect 276982 162757 277042 164598
rect 276979 162756 277045 162757
rect 276979 162692 276980 162756
rect 277044 162692 277045 162756
rect 276979 162691 277045 162692
rect 277166 161530 277226 164870
rect 278488 164658 278548 165106
rect 279168 164658 279228 165106
rect 280936 164930 280996 165106
rect 278454 164598 278548 164658
rect 279006 164598 279228 164658
rect 280846 164870 280996 164930
rect 278454 162213 278514 164598
rect 279006 162757 279066 164598
rect 279003 162756 279069 162757
rect 279003 162692 279004 162756
rect 279068 162692 279069 162756
rect 279003 162691 279069 162692
rect 278451 162212 278517 162213
rect 278451 162148 278452 162212
rect 278516 162148 278517 162212
rect 278451 162147 278517 162148
rect 277347 161532 277413 161533
rect 277347 161530 277348 161532
rect 277166 161470 277348 161530
rect 277347 161468 277348 161470
rect 277412 161468 277413 161532
rect 277347 161467 277413 161468
rect 275514 151878 275546 152114
rect 275782 151878 275866 152114
rect 276102 151878 276134 152114
rect 275514 151794 276134 151878
rect 275514 151558 275546 151794
rect 275782 151558 275866 151794
rect 276102 151558 276134 151794
rect 275514 145308 276134 151558
rect 279234 153954 279854 163000
rect 280846 162757 280906 164870
rect 283520 164658 283580 165106
rect 285968 164658 286028 165106
rect 288280 164661 288340 165106
rect 291000 164930 291060 165106
rect 293448 164930 293508 165106
rect 290966 164870 291060 164930
rect 293358 164870 293508 164930
rect 295896 164930 295956 165106
rect 298480 164930 298540 165106
rect 300928 164930 300988 165106
rect 303512 164930 303572 165106
rect 295896 164870 295994 164930
rect 298480 164870 298570 164930
rect 288277 164660 288343 164661
rect 283520 164598 283850 164658
rect 285968 164598 286058 164658
rect 280843 162756 280909 162757
rect 280843 162692 280844 162756
rect 280908 162692 280909 162756
rect 280843 162691 280909 162692
rect 279234 153718 279266 153954
rect 279502 153718 279586 153954
rect 279822 153718 279854 153954
rect 279234 153634 279854 153718
rect 279234 153398 279266 153634
rect 279502 153398 279586 153634
rect 279822 153398 279854 153634
rect 279234 145308 279854 153398
rect 282954 157674 283574 163000
rect 283790 162757 283850 164598
rect 285998 163845 286058 164598
rect 288277 164596 288278 164660
rect 288342 164596 288343 164660
rect 288277 164595 288343 164596
rect 290966 164389 291026 164870
rect 290963 164388 291029 164389
rect 290963 164324 290964 164388
rect 291028 164324 291029 164388
rect 290963 164323 291029 164324
rect 285995 163844 286061 163845
rect 285995 163780 285996 163844
rect 286060 163780 286061 163844
rect 285995 163779 286061 163780
rect 283787 162756 283853 162757
rect 283787 162692 283788 162756
rect 283852 162692 283853 162756
rect 283787 162691 283853 162692
rect 282954 157438 282986 157674
rect 283222 157438 283306 157674
rect 283542 157438 283574 157674
rect 282954 157354 283574 157438
rect 282954 157118 282986 157354
rect 283222 157118 283306 157354
rect 283542 157118 283574 157354
rect 282954 145308 283574 157118
rect 289794 147454 290414 163000
rect 293358 162757 293418 164870
rect 295934 163981 295994 164870
rect 298510 164253 298570 164870
rect 300902 164870 300988 164930
rect 303478 164870 303572 164930
rect 300902 164253 300962 164870
rect 303478 164253 303538 164870
rect 305960 164661 306020 165106
rect 308544 164930 308604 165106
rect 308446 164870 308604 164930
rect 310992 164930 311052 165106
rect 313440 164930 313500 165106
rect 315888 164930 315948 165106
rect 310992 164870 311082 164930
rect 305957 164660 306023 164661
rect 305957 164596 305958 164660
rect 306022 164596 306023 164660
rect 305957 164595 306023 164596
rect 298507 164252 298573 164253
rect 298507 164188 298508 164252
rect 298572 164188 298573 164252
rect 298507 164187 298573 164188
rect 300899 164252 300965 164253
rect 300899 164188 300900 164252
rect 300964 164188 300965 164252
rect 300899 164187 300965 164188
rect 303475 164252 303541 164253
rect 303475 164188 303476 164252
rect 303540 164188 303541 164252
rect 303475 164187 303541 164188
rect 308446 164117 308506 164870
rect 308443 164116 308509 164117
rect 308443 164052 308444 164116
rect 308508 164052 308509 164116
rect 308443 164051 308509 164052
rect 295931 163980 295997 163981
rect 295931 163916 295932 163980
rect 295996 163916 295997 163980
rect 295931 163915 295997 163916
rect 293355 162756 293421 162757
rect 293355 162692 293356 162756
rect 293420 162692 293421 162756
rect 293355 162691 293421 162692
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 145308 290414 146898
rect 293514 151174 294134 163000
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 145308 294134 150618
rect 297234 154894 297854 163000
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 145308 297854 154338
rect 300954 158614 301574 163000
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 145308 301574 158058
rect 307794 148394 308414 163000
rect 311022 162485 311082 164870
rect 313414 164870 313500 164930
rect 315070 164870 315948 164930
rect 313414 164253 313474 164870
rect 313411 164252 313477 164253
rect 313411 164188 313412 164252
rect 313476 164188 313477 164252
rect 313411 164187 313477 164188
rect 311019 162484 311085 162485
rect 311019 162420 311020 162484
rect 311084 162420 311085 162484
rect 311019 162419 311085 162420
rect 307794 148158 307826 148394
rect 308062 148158 308146 148394
rect 308382 148158 308414 148394
rect 307794 148074 308414 148158
rect 307794 147838 307826 148074
rect 308062 147838 308146 148074
rect 308382 147838 308414 148074
rect 307794 145308 308414 147838
rect 311514 152114 312134 163000
rect 315070 162349 315130 164870
rect 318472 164661 318532 165106
rect 320920 164930 320980 165106
rect 323368 164930 323428 165106
rect 320920 164870 321018 164930
rect 318469 164660 318535 164661
rect 318469 164596 318470 164660
rect 318534 164596 318535 164660
rect 318469 164595 318535 164596
rect 315067 162348 315133 162349
rect 315067 162284 315068 162348
rect 315132 162284 315133 162348
rect 315067 162283 315133 162284
rect 311514 151878 311546 152114
rect 311782 151878 311866 152114
rect 312102 151878 312134 152114
rect 311514 151794 312134 151878
rect 311514 151558 311546 151794
rect 311782 151558 311866 151794
rect 312102 151558 312134 151794
rect 311514 145308 312134 151558
rect 315234 153954 315854 163000
rect 315234 153718 315266 153954
rect 315502 153718 315586 153954
rect 315822 153718 315854 153954
rect 315234 153634 315854 153718
rect 315234 153398 315266 153634
rect 315502 153398 315586 153634
rect 315822 153398 315854 153634
rect 315234 145308 315854 153398
rect 318954 157674 319574 163000
rect 320958 162757 321018 164870
rect 323350 164870 323428 164930
rect 325952 164930 326012 165106
rect 343224 164930 343284 165106
rect 325952 164870 326722 164930
rect 320955 162756 321021 162757
rect 320955 162692 320956 162756
rect 321020 162692 321021 162756
rect 320955 162691 321021 162692
rect 323350 162621 323410 164870
rect 323347 162620 323413 162621
rect 323347 162556 323348 162620
rect 323412 162556 323413 162620
rect 323347 162555 323413 162556
rect 318954 157438 318986 157674
rect 319222 157438 319306 157674
rect 319542 157438 319574 157674
rect 318954 157354 319574 157438
rect 318954 157118 318986 157354
rect 319222 157118 319306 157354
rect 319542 157118 319574 157354
rect 318954 145308 319574 157118
rect 325794 147454 326414 163000
rect 326662 161805 326722 164870
rect 343222 164870 343284 164930
rect 343360 164930 343420 165106
rect 343360 164870 343466 164930
rect 326659 161804 326725 161805
rect 326659 161740 326660 161804
rect 326724 161740 326725 161804
rect 326659 161739 326725 161740
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 145308 326414 146898
rect 329514 151174 330134 163000
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 145308 330134 150618
rect 333234 154894 333854 163000
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 145308 333854 154338
rect 336954 158614 337574 163000
rect 343222 162621 343282 164870
rect 343406 162757 343466 164870
rect 343403 162756 343469 162757
rect 343403 162692 343404 162756
rect 343468 162692 343469 162756
rect 343403 162691 343469 162692
rect 343219 162620 343285 162621
rect 343219 162556 343220 162620
rect 343284 162556 343285 162620
rect 343219 162555 343285 162556
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 145308 337574 158058
rect 343794 148394 344414 163000
rect 343794 148158 343826 148394
rect 344062 148158 344146 148394
rect 344382 148158 344414 148394
rect 343794 148074 344414 148158
rect 343794 147838 343826 148074
rect 344062 147838 344146 148074
rect 344382 147838 344414 148074
rect 343794 145308 344414 147838
rect 347514 152114 348134 163000
rect 347514 151878 347546 152114
rect 347782 151878 347866 152114
rect 348102 151878 348134 152114
rect 347514 151794 348134 151878
rect 347514 151558 347546 151794
rect 347782 151558 347866 151794
rect 348102 151558 348134 151794
rect 347514 145308 348134 151558
rect 351234 153954 351854 163000
rect 351234 153718 351266 153954
rect 351502 153718 351586 153954
rect 351822 153718 351854 153954
rect 351234 153634 351854 153718
rect 351234 153398 351266 153634
rect 351502 153398 351586 153634
rect 351822 153398 351854 153634
rect 351234 145308 351854 153398
rect 354954 157674 355574 163000
rect 354954 157438 354986 157674
rect 355222 157438 355306 157674
rect 355542 157438 355574 157674
rect 354954 157354 355574 157438
rect 354954 157118 354986 157354
rect 355222 157118 355306 157354
rect 355542 157118 355574 157354
rect 354954 145308 355574 157118
rect 338435 144940 338501 144941
rect 338435 144876 338436 144940
rect 338500 144876 338501 144940
rect 338435 144875 338501 144876
rect 339723 144940 339789 144941
rect 339723 144876 339724 144940
rect 339788 144876 339789 144940
rect 339723 144875 339789 144876
rect 350947 144940 351013 144941
rect 350947 144876 350948 144940
rect 351012 144876 351013 144940
rect 350947 144875 351013 144876
rect 338438 143850 338498 144875
rect 339726 143850 339786 144875
rect 350950 143850 351010 144875
rect 338438 143790 338524 143850
rect 338464 143202 338524 143790
rect 339688 143790 339786 143850
rect 350840 143790 351010 143850
rect 339688 143202 339748 143790
rect 350840 143202 350900 143790
rect 220272 129454 220620 129486
rect 220272 129218 220328 129454
rect 220564 129218 220620 129454
rect 220272 129134 220620 129218
rect 220272 128898 220328 129134
rect 220564 128898 220620 129134
rect 220272 128866 220620 128898
rect 356000 129454 356348 129486
rect 356000 129218 356056 129454
rect 356292 129218 356348 129454
rect 356000 129134 356348 129218
rect 356000 128898 356056 129134
rect 356292 128898 356348 129134
rect 356000 128866 356348 128898
rect 220952 111454 221300 111486
rect 220952 111218 221008 111454
rect 221244 111218 221300 111454
rect 220952 111134 221300 111218
rect 220952 110898 221008 111134
rect 221244 110898 221300 111134
rect 220952 110866 221300 110898
rect 355320 111454 355668 111486
rect 355320 111218 355376 111454
rect 355612 111218 355668 111454
rect 355320 111134 355668 111218
rect 355320 110898 355376 111134
rect 355612 110898 355668 111134
rect 355320 110866 355668 110898
rect 220272 93454 220620 93486
rect 220272 93218 220328 93454
rect 220564 93218 220620 93454
rect 220272 93134 220620 93218
rect 220272 92898 220328 93134
rect 220564 92898 220620 93134
rect 220272 92866 220620 92898
rect 356000 93454 356348 93486
rect 356000 93218 356056 93454
rect 356292 93218 356348 93454
rect 356000 93134 356348 93218
rect 356000 92898 356056 93134
rect 356292 92898 356348 93134
rect 356000 92866 356348 92898
rect 220952 75454 221300 75486
rect 220952 75218 221008 75454
rect 221244 75218 221300 75454
rect 220952 75134 221300 75218
rect 220952 74898 221008 75134
rect 221244 74898 221300 75134
rect 220952 74866 221300 74898
rect 355320 75454 355668 75486
rect 355320 75218 355376 75454
rect 355612 75218 355668 75454
rect 355320 75134 355668 75218
rect 355320 74898 355376 75134
rect 355612 74898 355668 75134
rect 355320 74866 355668 74898
rect 236056 59530 236116 60106
rect 237144 59805 237204 60106
rect 237141 59804 237207 59805
rect 237141 59740 237142 59804
rect 237206 59740 237207 59804
rect 237141 59739 237207 59740
rect 238232 59530 238292 60106
rect 239592 59530 239652 60106
rect 235950 59470 236116 59530
rect 238158 59470 238292 59530
rect 239262 59470 239652 59530
rect 240544 59530 240604 60106
rect 241768 59530 241828 60106
rect 243128 59530 243188 60106
rect 240544 59470 240610 59530
rect 235950 58173 236010 59470
rect 235947 58172 236013 58173
rect 235947 58108 235948 58172
rect 236012 58108 236013 58172
rect 235947 58107 236013 58108
rect 219939 56540 220005 56541
rect 219939 56476 219940 56540
rect 220004 56476 220005 56540
rect 219939 56475 220005 56476
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 43174 222134 58000
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 46894 225854 58000
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 50614 229574 58000
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 57454 236414 58000
rect 238158 57901 238218 59470
rect 239262 57901 239322 59470
rect 238155 57900 238221 57901
rect 238155 57836 238156 57900
rect 238220 57836 238221 57900
rect 238155 57835 238221 57836
rect 239259 57900 239325 57901
rect 239259 57836 239260 57900
rect 239324 57836 239325 57900
rect 239259 57835 239325 57836
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 25174 240134 58000
rect 240550 57901 240610 59470
rect 241654 59470 241828 59530
rect 242942 59470 243188 59530
rect 244216 59530 244276 60106
rect 245440 59530 245500 60106
rect 246528 59530 246588 60106
rect 244216 59470 244290 59530
rect 241654 57901 241714 59470
rect 242942 57901 243002 59470
rect 240547 57900 240613 57901
rect 240547 57836 240548 57900
rect 240612 57836 240613 57900
rect 240547 57835 240613 57836
rect 241651 57900 241717 57901
rect 241651 57836 241652 57900
rect 241716 57836 241717 57900
rect 241651 57835 241717 57836
rect 242939 57900 243005 57901
rect 242939 57836 242940 57900
rect 243004 57836 243005 57900
rect 242939 57835 243005 57836
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 28894 243854 58000
rect 244230 57901 244290 59470
rect 245334 59470 245500 59530
rect 246438 59470 246588 59530
rect 247616 59530 247676 60106
rect 248296 59530 248356 60106
rect 248704 59530 248764 60106
rect 247616 59470 247786 59530
rect 245334 57901 245394 59470
rect 246438 57901 246498 59470
rect 244227 57900 244293 57901
rect 244227 57836 244228 57900
rect 244292 57836 244293 57900
rect 244227 57835 244293 57836
rect 245331 57900 245397 57901
rect 245331 57836 245332 57900
rect 245396 57836 245397 57900
rect 245331 57835 245397 57836
rect 246435 57900 246501 57901
rect 246435 57836 246436 57900
rect 246500 57836 246501 57900
rect 246435 57835 246501 57836
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 32614 247574 58000
rect 247726 57901 247786 59470
rect 248278 59470 248356 59530
rect 248646 59470 248764 59530
rect 250064 59530 250124 60106
rect 250744 59530 250804 60106
rect 251288 59530 251348 60106
rect 252376 59530 252436 60106
rect 253464 59530 253524 60106
rect 250064 59470 250178 59530
rect 247723 57900 247789 57901
rect 247723 57836 247724 57900
rect 247788 57836 247789 57900
rect 247723 57835 247789 57836
rect 248278 57085 248338 59470
rect 248646 57901 248706 59470
rect 250118 57901 250178 59470
rect 250670 59470 250804 59530
rect 251222 59470 251348 59530
rect 252326 59470 252436 59530
rect 253430 59470 253524 59530
rect 253600 59530 253660 60106
rect 254552 59530 254612 60106
rect 255912 59805 255972 60106
rect 255909 59804 255975 59805
rect 255909 59740 255910 59804
rect 255974 59740 255975 59804
rect 255909 59739 255975 59740
rect 256048 59530 256108 60106
rect 257000 59805 257060 60106
rect 256997 59804 257063 59805
rect 256997 59740 256998 59804
rect 257062 59740 257063 59804
rect 256997 59739 257063 59740
rect 258088 59530 258148 60106
rect 258496 59530 258556 60106
rect 253600 59470 253674 59530
rect 250670 58581 250730 59470
rect 250667 58580 250733 58581
rect 250667 58516 250668 58580
rect 250732 58516 250733 58580
rect 250667 58515 250733 58516
rect 251222 57901 251282 59470
rect 252326 57901 252386 59470
rect 253430 57901 253490 59470
rect 253614 58717 253674 59470
rect 254534 59470 254612 59530
rect 256006 59470 256108 59530
rect 257846 59470 258148 59530
rect 258398 59470 258556 59530
rect 259448 59530 259508 60106
rect 260672 59669 260732 60106
rect 260669 59668 260735 59669
rect 260669 59604 260670 59668
rect 260734 59604 260735 59668
rect 260669 59603 260735 59604
rect 261080 59530 261140 60106
rect 261760 59805 261820 60106
rect 261757 59804 261823 59805
rect 261757 59740 261758 59804
rect 261822 59740 261823 59804
rect 261757 59739 261823 59740
rect 262848 59533 262908 60106
rect 259448 59470 259562 59530
rect 253611 58716 253677 58717
rect 253611 58652 253612 58716
rect 253676 58652 253677 58716
rect 253611 58651 253677 58652
rect 248643 57900 248709 57901
rect 248643 57836 248644 57900
rect 248708 57836 248709 57900
rect 248643 57835 248709 57836
rect 250115 57900 250181 57901
rect 250115 57836 250116 57900
rect 250180 57836 250181 57900
rect 250115 57835 250181 57836
rect 251219 57900 251285 57901
rect 251219 57836 251220 57900
rect 251284 57836 251285 57900
rect 251219 57835 251285 57836
rect 252323 57900 252389 57901
rect 252323 57836 252324 57900
rect 252388 57836 252389 57900
rect 252323 57835 252389 57836
rect 253427 57900 253493 57901
rect 253427 57836 253428 57900
rect 253492 57836 253493 57900
rect 253427 57835 253493 57836
rect 248275 57084 248341 57085
rect 248275 57020 248276 57084
rect 248340 57020 248341 57084
rect 248275 57019 248341 57020
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 39454 254414 58000
rect 254534 57901 254594 59470
rect 254531 57900 254597 57901
rect 254531 57836 254532 57900
rect 254596 57836 254597 57900
rect 254531 57835 254597 57836
rect 256006 57357 256066 59470
rect 257846 58445 257906 59470
rect 257843 58444 257909 58445
rect 257843 58380 257844 58444
rect 257908 58380 257909 58444
rect 257843 58379 257909 58380
rect 256003 57356 256069 57357
rect 256003 57292 256004 57356
rect 256068 57292 256069 57356
rect 256003 57291 256069 57292
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 43174 258134 58000
rect 258398 57493 258458 59470
rect 259502 58717 259562 59470
rect 260974 59470 261140 59530
rect 262811 59532 262908 59533
rect 259499 58716 259565 58717
rect 259499 58652 259500 58716
rect 259564 58652 259565 58716
rect 259499 58651 259565 58652
rect 258395 57492 258461 57493
rect 258395 57428 258396 57492
rect 258460 57428 258461 57492
rect 258395 57427 258461 57428
rect 260974 57221 261034 59470
rect 262811 59468 262812 59532
rect 262876 59470 262908 59532
rect 263528 59530 263588 60106
rect 263936 59805 263996 60106
rect 263933 59804 263999 59805
rect 263933 59740 263934 59804
rect 263998 59740 263999 59804
rect 263933 59739 263999 59740
rect 265296 59530 265356 60106
rect 265976 59530 266036 60106
rect 266384 59530 266444 60106
rect 267608 59530 267668 60106
rect 263528 59470 263610 59530
rect 262876 59468 262877 59470
rect 262811 59467 262877 59468
rect 263550 59397 263610 59470
rect 265206 59470 265356 59530
rect 265942 59470 266036 59530
rect 266310 59470 266444 59530
rect 267598 59470 267668 59530
rect 268288 59530 268348 60106
rect 268696 59530 268756 60106
rect 269784 59530 269844 60106
rect 271008 59530 271068 60106
rect 268288 59470 268394 59530
rect 268696 59470 268762 59530
rect 269784 59470 269866 59530
rect 263547 59396 263613 59397
rect 263547 59332 263548 59396
rect 263612 59332 263613 59396
rect 263547 59331 263613 59332
rect 265206 58173 265266 59470
rect 265203 58172 265269 58173
rect 265203 58108 265204 58172
rect 265268 58108 265269 58172
rect 265203 58107 265269 58108
rect 260971 57220 261037 57221
rect 260971 57156 260972 57220
rect 261036 57156 261037 57220
rect 260971 57155 261037 57156
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 46894 261854 58000
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 50614 265574 58000
rect 265942 57901 266002 59470
rect 266310 57901 266370 59470
rect 265939 57900 266005 57901
rect 265939 57836 265940 57900
rect 266004 57836 266005 57900
rect 265939 57835 266005 57836
rect 266307 57900 266373 57901
rect 266307 57836 266308 57900
rect 266372 57836 266373 57900
rect 266307 57835 266373 57836
rect 267598 57629 267658 59470
rect 267595 57628 267661 57629
rect 267595 57564 267596 57628
rect 267660 57564 267661 57628
rect 267595 57563 267661 57564
rect 268334 56405 268394 59470
rect 268702 57901 268762 59470
rect 268699 57900 268765 57901
rect 268699 57836 268700 57900
rect 268764 57836 268765 57900
rect 268699 57835 268765 57836
rect 269806 57629 269866 59470
rect 270910 59470 271068 59530
rect 271144 59530 271204 60106
rect 272232 59530 272292 60106
rect 273320 59530 273380 60106
rect 273592 59530 273652 60106
rect 274408 59530 274468 60106
rect 275768 59530 275828 60106
rect 271144 59470 271338 59530
rect 269803 57628 269869 57629
rect 269803 57564 269804 57628
rect 269868 57564 269869 57628
rect 269803 57563 269869 57564
rect 270910 57493 270970 59470
rect 271278 57901 271338 59470
rect 272198 59470 272292 59530
rect 273302 59470 273380 59530
rect 273486 59470 273652 59530
rect 274406 59470 274468 59530
rect 275694 59470 275828 59530
rect 276040 59530 276100 60106
rect 276992 59530 277052 60106
rect 278080 59530 278140 60106
rect 278488 59530 278548 60106
rect 276040 59470 276122 59530
rect 272198 58173 272258 59470
rect 272195 58172 272261 58173
rect 272195 58108 272196 58172
rect 272260 58108 272261 58172
rect 272195 58107 272261 58108
rect 271275 57900 271341 57901
rect 271275 57836 271276 57900
rect 271340 57836 271341 57900
rect 271275 57835 271341 57836
rect 270907 57492 270973 57493
rect 270907 57428 270908 57492
rect 270972 57428 270973 57492
rect 270907 57427 270973 57428
rect 271794 57454 272414 58000
rect 273302 57901 273362 59470
rect 273486 59125 273546 59470
rect 273483 59124 273549 59125
rect 273483 59060 273484 59124
rect 273548 59060 273549 59124
rect 273483 59059 273549 59060
rect 273299 57900 273365 57901
rect 273299 57836 273300 57900
rect 273364 57836 273365 57900
rect 273299 57835 273365 57836
rect 274406 57629 274466 59470
rect 275694 58173 275754 59470
rect 276062 58989 276122 59470
rect 276982 59470 277052 59530
rect 277902 59470 278140 59530
rect 278454 59470 278548 59530
rect 279168 59530 279228 60106
rect 280936 59530 280996 60106
rect 279168 59470 279250 59530
rect 276059 58988 276125 58989
rect 276059 58924 276060 58988
rect 276124 58924 276125 58988
rect 276059 58923 276125 58924
rect 275691 58172 275757 58173
rect 275691 58108 275692 58172
rect 275756 58108 275757 58172
rect 275691 58107 275757 58108
rect 274403 57628 274469 57629
rect 274403 57564 274404 57628
rect 274468 57564 274469 57628
rect 274403 57563 274469 57564
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 268331 56404 268397 56405
rect 268331 56340 268332 56404
rect 268396 56340 268397 56404
rect 268331 56339 268397 56340
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 25174 276134 58000
rect 276982 57629 277042 59470
rect 277902 57990 277962 59470
rect 278454 58853 278514 59470
rect 279190 59261 279250 59470
rect 280846 59470 280996 59530
rect 283520 59530 283580 60106
rect 285968 59530 286028 60106
rect 288280 59530 288340 60106
rect 291000 59530 291060 60106
rect 293448 59530 293508 60106
rect 283520 59470 283850 59530
rect 285968 59470 286058 59530
rect 279187 59260 279253 59261
rect 279187 59196 279188 59260
rect 279252 59196 279253 59260
rect 279187 59195 279253 59196
rect 278451 58852 278517 58853
rect 278451 58788 278452 58852
rect 278516 58788 278517 58852
rect 278451 58787 278517 58788
rect 277166 57930 277962 57990
rect 276979 57628 277045 57629
rect 276979 57564 276980 57628
rect 277044 57564 277045 57628
rect 276979 57563 277045 57564
rect 277166 56269 277226 57930
rect 277163 56268 277229 56269
rect 277163 56204 277164 56268
rect 277228 56204 277229 56268
rect 277163 56203 277229 56204
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 28894 279854 58000
rect 280846 57765 280906 59470
rect 280843 57764 280909 57765
rect 280843 57700 280844 57764
rect 280908 57700 280909 57764
rect 280843 57699 280909 57700
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 32614 283574 58000
rect 283790 56677 283850 59470
rect 285998 59125 286058 59470
rect 288206 59470 288340 59530
rect 290966 59470 291060 59530
rect 293358 59470 293508 59530
rect 295896 59530 295956 60106
rect 298480 59530 298540 60106
rect 300928 59530 300988 60106
rect 303512 59530 303572 60106
rect 305960 59669 306020 60106
rect 305957 59668 306023 59669
rect 305957 59604 305958 59668
rect 306022 59604 306023 59668
rect 305957 59603 306023 59604
rect 295896 59470 295994 59530
rect 298480 59470 298570 59530
rect 285995 59124 286061 59125
rect 285995 59060 285996 59124
rect 286060 59060 286061 59124
rect 285995 59059 286061 59060
rect 288206 57901 288266 59470
rect 290966 59261 291026 59470
rect 290963 59260 291029 59261
rect 290963 59196 290964 59260
rect 291028 59196 291029 59260
rect 290963 59195 291029 59196
rect 288203 57900 288269 57901
rect 288203 57836 288204 57900
rect 288268 57836 288269 57900
rect 288203 57835 288269 57836
rect 283787 56676 283853 56677
rect 283787 56612 283788 56676
rect 283852 56612 283853 56676
rect 283787 56611 283853 56612
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 39454 290414 58000
rect 293358 57901 293418 59470
rect 293355 57900 293421 57901
rect 293355 57836 293356 57900
rect 293420 57836 293421 57900
rect 293355 57835 293421 57836
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 43174 294134 58000
rect 295934 57901 295994 59470
rect 298510 59261 298570 59470
rect 300902 59470 300988 59530
rect 303478 59470 303572 59530
rect 308544 59530 308604 60106
rect 310992 59530 311052 60106
rect 313440 59530 313500 60106
rect 315888 59530 315948 60106
rect 318472 59669 318532 60106
rect 318469 59668 318535 59669
rect 318469 59604 318470 59668
rect 318534 59604 318535 59668
rect 318469 59603 318535 59604
rect 308544 59470 308690 59530
rect 310992 59470 311082 59530
rect 298507 59260 298573 59261
rect 298507 59196 298508 59260
rect 298572 59196 298573 59260
rect 298507 59195 298573 59196
rect 300902 58173 300962 59470
rect 300899 58172 300965 58173
rect 300899 58108 300900 58172
rect 300964 58108 300965 58172
rect 300899 58107 300965 58108
rect 295931 57900 295997 57901
rect 295931 57836 295932 57900
rect 295996 57836 295997 57900
rect 295931 57835 295997 57836
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 46894 297854 58000
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 50614 301574 58000
rect 303478 57901 303538 59470
rect 303475 57900 303541 57901
rect 303475 57836 303476 57900
rect 303540 57836 303541 57900
rect 303475 57835 303541 57836
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 57454 308414 58000
rect 308630 57901 308690 59470
rect 311022 57901 311082 59470
rect 313414 59470 313500 59530
rect 315806 59470 315948 59530
rect 320920 59530 320980 60106
rect 323368 59530 323428 60106
rect 325952 59530 326012 60106
rect 343224 59530 343284 60106
rect 320920 59470 321018 59530
rect 313414 59261 313474 59470
rect 313411 59260 313477 59261
rect 313411 59196 313412 59260
rect 313476 59196 313477 59260
rect 313411 59195 313477 59196
rect 315806 58173 315866 59470
rect 315803 58172 315869 58173
rect 315803 58108 315804 58172
rect 315868 58108 315869 58172
rect 315803 58107 315869 58108
rect 308627 57900 308693 57901
rect 308627 57836 308628 57900
rect 308692 57836 308693 57900
rect 308627 57835 308693 57836
rect 311019 57900 311085 57901
rect 311019 57836 311020 57900
rect 311084 57836 311085 57900
rect 311019 57835 311085 57836
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 25174 312134 58000
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 28894 315854 58000
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 32614 319574 58000
rect 320958 57901 321018 59470
rect 323350 59470 323428 59530
rect 325926 59470 326012 59530
rect 343222 59470 343284 59530
rect 343360 59530 343420 60106
rect 343360 59470 343466 59530
rect 323350 57901 323410 59470
rect 325926 59261 325986 59470
rect 325923 59260 325989 59261
rect 325923 59196 325924 59260
rect 325988 59196 325989 59260
rect 325923 59195 325989 59196
rect 320955 57900 321021 57901
rect 320955 57836 320956 57900
rect 321020 57836 321021 57900
rect 320955 57835 321021 57836
rect 323347 57900 323413 57901
rect 323347 57836 323348 57900
rect 323412 57836 323413 57900
rect 323347 57835 323413 57836
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 39454 326414 58000
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 43174 330134 58000
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 46894 333854 58000
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 50614 337574 58000
rect 343222 57901 343282 59470
rect 343406 57901 343466 59470
rect 357942 59125 358002 477939
rect 358123 477868 358189 477869
rect 358123 477804 358124 477868
rect 358188 477804 358189 477868
rect 358123 477803 358189 477804
rect 358126 407829 358186 477803
rect 359411 476916 359477 476917
rect 359411 476852 359412 476916
rect 359476 476852 359477 476916
rect 359411 476851 359477 476852
rect 358123 407828 358189 407829
rect 358123 407764 358124 407828
rect 358188 407764 358189 407828
rect 358123 407763 358189 407764
rect 359414 268973 359474 476851
rect 359595 469844 359661 469845
rect 359595 469780 359596 469844
rect 359660 469780 359661 469844
rect 359595 469779 359661 469780
rect 359598 269245 359658 469779
rect 359779 461548 359845 461549
rect 359779 461484 359780 461548
rect 359844 461484 359845 461548
rect 359779 461483 359845 461484
rect 359782 279989 359842 461483
rect 359963 460324 360029 460325
rect 359963 460260 359964 460324
rect 360028 460260 360029 460324
rect 359963 460259 360029 460260
rect 359966 374645 360026 460259
rect 359963 374644 360029 374645
rect 359963 374580 359964 374644
rect 360028 374580 360029 374644
rect 359963 374579 360029 374580
rect 359779 279988 359845 279989
rect 359779 279924 359780 279988
rect 359844 279924 359845 279988
rect 359779 279923 359845 279924
rect 359595 269244 359661 269245
rect 359595 269180 359596 269244
rect 359660 269180 359661 269244
rect 359595 269179 359661 269180
rect 359411 268972 359477 268973
rect 359411 268908 359412 268972
rect 359476 268908 359477 268972
rect 359411 268907 359477 268908
rect 360702 59261 360762 478755
rect 360886 149157 360946 485011
rect 361794 471454 362414 506898
rect 365514 511174 366134 518000
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 363459 483716 363525 483717
rect 363459 483652 363460 483716
rect 363524 483652 363525 483716
rect 363459 483651 363525 483652
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 360883 149156 360949 149157
rect 360883 149092 360884 149156
rect 360948 149092 360949 149156
rect 360883 149091 360949 149092
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 360699 59260 360765 59261
rect 360699 59196 360700 59260
rect 360764 59196 360765 59260
rect 360699 59195 360765 59196
rect 357939 59124 358005 59125
rect 357939 59060 357940 59124
rect 358004 59060 358005 59124
rect 357939 59059 358005 59060
rect 343219 57900 343285 57901
rect 343219 57836 343220 57900
rect 343284 57836 343285 57900
rect 343219 57835 343285 57836
rect 343403 57900 343469 57901
rect 343403 57836 343404 57900
rect 343468 57836 343469 57900
rect 343403 57835 343469 57836
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 57454 344414 58000
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 25174 348134 58000
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 28894 351854 58000
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 32614 355574 58000
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 363462 3637 363522 483651
rect 364931 482220 364997 482221
rect 364931 482156 364932 482220
rect 364996 482156 364997 482220
rect 364931 482155 364997 482156
rect 363643 474196 363709 474197
rect 363643 474132 363644 474196
rect 363708 474132 363709 474196
rect 363643 474131 363709 474132
rect 363646 56677 363706 474131
rect 363643 56676 363709 56677
rect 363643 56612 363644 56676
rect 363708 56612 363709 56676
rect 363643 56611 363709 56612
rect 363459 3636 363525 3637
rect 363459 3572 363460 3636
rect 363524 3572 363525 3636
rect 363459 3571 363525 3572
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 364934 3365 364994 482155
rect 365115 479772 365181 479773
rect 365115 479708 365116 479772
rect 365180 479708 365181 479772
rect 365115 479707 365181 479708
rect 365118 3773 365178 479707
rect 365514 475174 366134 510618
rect 369234 514894 369854 518000
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 372954 482614 373574 518000
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 369234 478574 369854 478658
rect 371739 478684 371805 478685
rect 371739 478620 371740 478684
rect 371804 478620 371805 478684
rect 371739 478619 371805 478620
rect 367691 478548 367757 478549
rect 367691 478484 367692 478548
rect 367756 478484 367757 478548
rect 367691 478483 367757 478484
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 367694 58445 367754 478483
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 370451 478412 370517 478413
rect 370451 478348 370452 478412
rect 370516 478348 370517 478412
rect 370451 478347 370517 478348
rect 367875 476780 367941 476781
rect 367875 476716 367876 476780
rect 367940 476716 367941 476780
rect 367875 476715 367941 476716
rect 367878 68101 367938 476715
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 367875 68100 367941 68101
rect 367875 68036 367876 68100
rect 367940 68036 367941 68100
rect 367875 68035 367941 68036
rect 367691 58444 367757 58445
rect 367691 58380 367692 58444
rect 367756 58380 367757 58444
rect 367691 58379 367757 58380
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365115 3772 365181 3773
rect 365115 3708 365116 3772
rect 365180 3708 365181 3772
rect 365115 3707 365181 3708
rect 364931 3364 364997 3365
rect 364931 3300 364932 3364
rect 364996 3300 364997 3364
rect 364931 3299 364997 3300
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 46894 369854 82338
rect 370454 58717 370514 478347
rect 371742 58989 371802 478619
rect 371923 475556 371989 475557
rect 371923 475492 371924 475556
rect 371988 475492 371989 475556
rect 371923 475491 371989 475492
rect 371739 58988 371805 58989
rect 371739 58924 371740 58988
rect 371804 58924 371805 58988
rect 371739 58923 371805 58924
rect 370451 58716 370517 58717
rect 370451 58652 370452 58716
rect 370516 58652 370517 58716
rect 370451 58651 370517 58652
rect 371926 57629 371986 475491
rect 372954 446614 373574 482058
rect 379794 489454 380414 518000
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 374499 478412 374565 478413
rect 374499 478348 374500 478412
rect 374564 478348 374565 478412
rect 374499 478347 374565 478348
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 357554 373574 374058
rect 372954 357318 372986 357554
rect 373222 357318 373306 357554
rect 373542 357318 373574 357554
rect 372954 357234 373574 357318
rect 372954 356998 372986 357234
rect 373222 356998 373306 357234
rect 373542 356998 373574 357234
rect 372954 338614 373574 356998
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 371923 57628 371989 57629
rect 371923 57564 371924 57628
rect 371988 57564 371989 57628
rect 371923 57563 371989 57564
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 374502 3501 374562 478347
rect 375971 478276 376037 478277
rect 375971 478212 375972 478276
rect 376036 478212 376037 478276
rect 375971 478211 376037 478212
rect 374683 478140 374749 478141
rect 374683 478076 374684 478140
rect 374748 478076 374749 478140
rect 374683 478075 374749 478076
rect 374686 58581 374746 478075
rect 375974 58853 376034 478211
rect 377259 474332 377325 474333
rect 377259 474268 377260 474332
rect 377324 474268 377325 474332
rect 377259 474267 377325 474268
rect 376155 465764 376221 465765
rect 376155 465700 376156 465764
rect 376220 465700 376221 465764
rect 376155 465699 376221 465700
rect 375971 58852 376037 58853
rect 375971 58788 375972 58852
rect 376036 58788 376037 58852
rect 375971 58787 376037 58788
rect 374683 58580 374749 58581
rect 374683 58516 374684 58580
rect 374748 58516 374749 58580
rect 374683 58515 374749 58516
rect 376158 57357 376218 465699
rect 376891 462908 376957 462909
rect 376891 462844 376892 462908
rect 376956 462844 376957 462908
rect 376891 462843 376957 462844
rect 376894 372741 376954 462843
rect 376891 372740 376957 372741
rect 376891 372676 376892 372740
rect 376956 372676 376957 372740
rect 376891 372675 376957 372676
rect 376891 368524 376957 368525
rect 376891 368460 376892 368524
rect 376956 368460 376957 368524
rect 376891 368459 376957 368460
rect 376894 269381 376954 368459
rect 376891 269380 376957 269381
rect 376891 269316 376892 269380
rect 376956 269316 376957 269380
rect 376891 269315 376957 269316
rect 377262 267341 377322 474267
rect 379467 472564 379533 472565
rect 379467 472500 379468 472564
rect 379532 472500 379533 472564
rect 379467 472499 379533 472500
rect 378731 471204 378797 471205
rect 378731 471140 378732 471204
rect 378796 471140 378797 471204
rect 378731 471139 378797 471140
rect 377443 465900 377509 465901
rect 377443 465836 377444 465900
rect 377508 465836 377509 465900
rect 377443 465835 377509 465836
rect 377446 371925 377506 465835
rect 377627 460188 377693 460189
rect 377627 460124 377628 460188
rect 377692 460124 377693 460188
rect 377627 460123 377693 460124
rect 377630 373965 377690 460123
rect 377627 373964 377693 373965
rect 377627 373900 377628 373964
rect 377692 373900 377693 373964
rect 377627 373899 377693 373900
rect 377443 371924 377509 371925
rect 377443 371860 377444 371924
rect 377508 371860 377509 371924
rect 377443 371859 377509 371860
rect 377995 269380 378061 269381
rect 377995 269316 377996 269380
rect 378060 269316 378061 269380
rect 377995 269315 378061 269316
rect 377998 268837 378058 269315
rect 377995 268836 378061 268837
rect 377995 268772 377996 268836
rect 378060 268772 378061 268836
rect 377995 268771 378061 268772
rect 377259 267340 377325 267341
rect 377259 267276 377260 267340
rect 377324 267276 377325 267340
rect 377259 267275 377325 267276
rect 377995 251020 378061 251021
rect 377995 250956 377996 251020
rect 378060 250956 378061 251020
rect 377995 250955 378061 250956
rect 377627 148340 377693 148341
rect 377627 148276 377628 148340
rect 377692 148276 377693 148340
rect 377627 148275 377693 148276
rect 376155 57356 376221 57357
rect 376155 57292 376156 57356
rect 376220 57292 376221 57356
rect 376155 57291 376221 57292
rect 377630 55181 377690 148275
rect 377998 146301 378058 250955
rect 377995 146300 378061 146301
rect 377995 146236 377996 146300
rect 378060 146236 378061 146300
rect 377995 146235 378061 146236
rect 377811 145620 377877 145621
rect 377811 145556 377812 145620
rect 377876 145556 377877 145620
rect 377811 145555 377877 145556
rect 377814 59397 377874 145555
rect 377811 59396 377877 59397
rect 377811 59332 377812 59396
rect 377876 59332 377877 59396
rect 377811 59331 377877 59332
rect 378734 57765 378794 471139
rect 379470 470610 379530 472499
rect 379470 470550 379714 470610
rect 378915 468484 378981 468485
rect 378915 468420 378916 468484
rect 378980 468420 378981 468484
rect 378915 468419 378981 468420
rect 378731 57764 378797 57765
rect 378731 57700 378732 57764
rect 378796 57700 378797 57764
rect 378731 57699 378797 57700
rect 378918 57493 378978 468419
rect 379099 458964 379165 458965
rect 379099 458900 379100 458964
rect 379164 458900 379165 458964
rect 379099 458899 379165 458900
rect 378915 57492 378981 57493
rect 378915 57428 378916 57492
rect 378980 57428 378981 57492
rect 378915 57427 378981 57428
rect 379102 57085 379162 458899
rect 379283 458828 379349 458829
rect 379283 458764 379284 458828
rect 379348 458764 379349 458828
rect 379283 458763 379349 458764
rect 379286 57221 379346 458763
rect 379654 267750 379714 470550
rect 379794 460308 380414 488898
rect 383514 493174 384134 518000
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 460308 384134 492618
rect 387234 496894 387854 518000
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460308 387854 496338
rect 390954 500614 391574 518000
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 460308 391574 464058
rect 397794 507454 398414 518000
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 460308 398414 470898
rect 401514 511174 402134 518000
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 460308 402134 474618
rect 405234 514894 405854 518000
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 460308 405854 478338
rect 408954 482614 409574 518000
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 460308 409574 482058
rect 415794 489454 416414 518000
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 460308 416414 488898
rect 419514 493174 420134 518000
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 460308 420134 492618
rect 423234 496894 423854 518000
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460308 423854 496338
rect 426954 500614 427574 518000
rect 430990 517309 431050 592179
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 430987 517308 431053 517309
rect 430987 517244 430988 517308
rect 431052 517244 431053 517308
rect 430987 517243 431053 517244
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 460308 427574 464058
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 460308 434414 470898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 460308 438134 474618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 460308 441854 478338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 460308 445574 482058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 460308 452414 488898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 622000 459854 640338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 622000 463574 644058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 622000 470414 650898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 622000 474134 654618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 622000 477854 622338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 622000 481574 626058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 622000 488414 632898
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 622000 492134 636618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 622000 495854 640338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 622000 499574 644058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 622000 506414 650898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 622000 510134 654618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 476067 619988 476133 619989
rect 476067 619924 476068 619988
rect 476132 619924 476133 619988
rect 476067 619923 476133 619924
rect 488579 619988 488645 619989
rect 488579 619924 488580 619988
rect 488644 619924 488645 619988
rect 488579 619923 488645 619924
rect 506611 619988 506677 619989
rect 506611 619924 506612 619988
rect 506676 619924 506677 619988
rect 506611 619923 506677 619924
rect 464208 615454 464528 615486
rect 464208 615218 464250 615454
rect 464486 615218 464528 615454
rect 464208 615134 464528 615218
rect 464208 614898 464250 615134
rect 464486 614898 464528 615134
rect 464208 614866 464528 614898
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 464208 579454 464528 579486
rect 464208 579218 464250 579454
rect 464486 579218 464528 579454
rect 464208 579134 464528 579218
rect 464208 578898 464250 579134
rect 464486 578898 464528 579134
rect 464208 578866 464528 578898
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 460308 456134 492618
rect 459234 532894 459854 568000
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460308 459854 496338
rect 462954 536614 463574 568000
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 460308 463574 464058
rect 469794 543454 470414 568000
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 460308 470414 470898
rect 473514 547174 474134 568000
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 476070 479501 476130 619923
rect 479568 597454 479888 597486
rect 479568 597218 479610 597454
rect 479846 597218 479888 597454
rect 479568 597134 479888 597218
rect 479568 596898 479610 597134
rect 479846 596898 479888 597134
rect 479568 596866 479888 596898
rect 477234 550894 477854 568000
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 476067 479500 476133 479501
rect 476067 479436 476068 479500
rect 476132 479436 476133 479500
rect 476067 479435 476133 479436
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 460308 474134 474618
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 460308 477854 478338
rect 480954 554614 481574 568000
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 460308 481574 482058
rect 487794 561454 488414 568000
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 460308 488414 488898
rect 488582 483717 488642 619923
rect 494928 615454 495248 615486
rect 494928 615218 494970 615454
rect 495206 615218 495248 615454
rect 494928 615134 495248 615218
rect 494928 614898 494970 615134
rect 495206 614898 495248 615134
rect 494928 614866 495248 614898
rect 494928 579454 495248 579486
rect 494928 579218 494970 579454
rect 495206 579218 495248 579454
rect 494928 579134 495248 579218
rect 494928 578898 494970 579134
rect 495206 578898 495248 579134
rect 494928 578866 495248 578898
rect 491514 565174 492134 568000
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 488579 483716 488645 483717
rect 488579 483652 488580 483716
rect 488644 483652 488645 483716
rect 488579 483651 488645 483652
rect 491514 460308 492134 492618
rect 495234 532894 495854 568000
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460308 495854 496338
rect 498954 536614 499574 568000
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498515 461004 498581 461005
rect 498515 460940 498516 461004
rect 498580 460940 498581 461004
rect 498515 460939 498581 460940
rect 498518 458690 498578 460939
rect 498954 460308 499574 464058
rect 505794 543454 506414 568000
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 506614 480861 506674 619923
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 509514 547174 510134 568000
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 506611 480860 506677 480861
rect 506611 480796 506612 480860
rect 506676 480796 506677 480860
rect 506611 480795 506677 480796
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 499803 461004 499869 461005
rect 499803 460940 499804 461004
rect 499868 460940 499869 461004
rect 499803 460939 499869 460940
rect 499806 458690 499866 460939
rect 505794 460308 506414 470898
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 460308 510134 474618
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 510843 461004 510909 461005
rect 510843 460940 510844 461004
rect 510908 460940 510909 461004
rect 510843 460939 510909 460940
rect 510846 458690 510906 460939
rect 513234 460308 513854 478338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 460308 517574 482058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 498464 458630 498578 458690
rect 499688 458630 499866 458690
rect 510840 458630 510906 458690
rect 498464 458202 498524 458630
rect 499688 458202 499748 458630
rect 510840 458202 510900 458630
rect 380272 453454 380620 453486
rect 380272 453218 380328 453454
rect 380564 453218 380620 453454
rect 380272 453134 380620 453218
rect 380272 452898 380328 453134
rect 380564 452898 380620 453134
rect 380272 452866 380620 452898
rect 516000 453454 516348 453486
rect 516000 453218 516056 453454
rect 516292 453218 516348 453454
rect 516000 453134 516348 453218
rect 516000 452898 516056 453134
rect 516292 452898 516348 453134
rect 516000 452866 516348 452898
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 380952 435454 381300 435486
rect 380952 435218 381008 435454
rect 381244 435218 381300 435454
rect 380952 435134 381300 435218
rect 380952 434898 381008 435134
rect 381244 434898 381300 435134
rect 380952 434866 381300 434898
rect 515320 435454 515668 435486
rect 515320 435218 515376 435454
rect 515612 435218 515668 435454
rect 515320 435134 515668 435218
rect 515320 434898 515376 435134
rect 515612 434898 515668 435134
rect 515320 434866 515668 434898
rect 380272 417454 380620 417486
rect 380272 417218 380328 417454
rect 380564 417218 380620 417454
rect 380272 417134 380620 417218
rect 380272 416898 380328 417134
rect 380564 416898 380620 417134
rect 380272 416866 380620 416898
rect 516000 417454 516348 417486
rect 516000 417218 516056 417454
rect 516292 417218 516348 417454
rect 516000 417134 516348 417218
rect 516000 416898 516056 417134
rect 516292 416898 516348 417134
rect 516000 416866 516348 416898
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 380952 399454 381300 399486
rect 380952 399218 381008 399454
rect 381244 399218 381300 399454
rect 380952 399134 381300 399218
rect 380952 398898 381008 399134
rect 381244 398898 381300 399134
rect 380952 398866 381300 398898
rect 515320 399454 515668 399486
rect 515320 399218 515376 399454
rect 515612 399218 515668 399454
rect 515320 399134 515668 399218
rect 515320 398898 515376 399134
rect 515612 398898 515668 399134
rect 515320 398866 515668 398898
rect 380272 381454 380620 381486
rect 380272 381218 380328 381454
rect 380564 381218 380620 381454
rect 380272 381134 380620 381218
rect 380272 380898 380328 381134
rect 380564 380898 380620 381134
rect 380272 380866 380620 380898
rect 516000 381454 516348 381486
rect 516000 381218 516056 381454
rect 516292 381218 516348 381454
rect 516000 381134 516348 381218
rect 516000 380898 516056 381134
rect 516292 380898 516348 381134
rect 516000 380866 516348 380898
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 407803 375052 407869 375053
rect 396086 374990 396274 375050
rect 379794 364394 380414 373000
rect 379794 364158 379826 364394
rect 380062 364158 380146 364394
rect 380382 364158 380414 364394
rect 379794 364074 380414 364158
rect 379794 363838 379826 364074
rect 380062 363838 380146 364074
rect 380382 363838 380414 364074
rect 379794 355308 380414 363838
rect 383514 366234 384134 373000
rect 383514 365998 383546 366234
rect 383782 365998 383866 366234
rect 384102 365998 384134 366234
rect 383514 365914 384134 365998
rect 383514 365678 383546 365914
rect 383782 365678 383866 365914
rect 384102 365678 384134 365914
rect 383514 355308 384134 365678
rect 387234 369954 387854 373000
rect 387234 369718 387266 369954
rect 387502 369718 387586 369954
rect 387822 369718 387854 369954
rect 387234 369634 387854 369718
rect 387234 369398 387266 369634
rect 387502 369398 387586 369634
rect 387822 369398 387854 369634
rect 387234 355308 387854 369398
rect 390954 356614 391574 373000
rect 396214 372061 396274 374990
rect 396582 374990 397174 375050
rect 397502 374990 398262 375050
rect 398974 374990 399622 375050
rect 400262 374990 400574 375050
rect 401798 374990 402346 375050
rect 396211 372060 396277 372061
rect 396211 371996 396212 372060
rect 396276 371996 396277 372060
rect 396211 371995 396277 371996
rect 396582 371381 396642 374990
rect 397502 372061 397562 374990
rect 397499 372060 397565 372061
rect 397499 371996 397500 372060
rect 397564 371996 397565 372060
rect 397499 371995 397565 371996
rect 396579 371380 396645 371381
rect 396579 371316 396580 371380
rect 396644 371316 396645 371380
rect 396579 371315 396645 371316
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 355308 391574 356058
rect 397794 363454 398414 373000
rect 398974 372061 399034 374990
rect 400262 372061 400322 374990
rect 398971 372060 399037 372061
rect 398971 371996 398972 372060
rect 399036 371996 399037 372060
rect 398971 371995 399037 371996
rect 400259 372060 400325 372061
rect 400259 371996 400260 372060
rect 400324 371996 400325 372060
rect 400259 371995 400325 371996
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 355308 398414 362898
rect 401514 367174 402134 373000
rect 402286 371653 402346 374990
rect 403022 374990 403158 375050
rect 402283 371652 402349 371653
rect 402283 371588 402284 371652
rect 402348 371588 402349 371652
rect 402283 371587 402349 371588
rect 403022 371381 403082 374990
rect 404216 374781 404276 375020
rect 404862 374990 405470 375050
rect 406150 374990 406558 375050
rect 407254 374990 407646 375050
rect 404213 374780 404279 374781
rect 404213 374716 404214 374780
rect 404278 374716 404279 374780
rect 404213 374715 404279 374716
rect 404862 372197 404922 374990
rect 404859 372196 404925 372197
rect 404859 372132 404860 372196
rect 404924 372132 404925 372196
rect 404859 372131 404925 372132
rect 403019 371380 403085 371381
rect 403019 371316 403020 371380
rect 403084 371316 403085 371380
rect 403019 371315 403085 371316
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 355308 402134 366618
rect 405234 370894 405854 373000
rect 406150 371381 406210 374990
rect 407254 371517 407314 374990
rect 407803 374988 407804 375052
rect 407868 375050 407869 375052
rect 425099 375052 425165 375053
rect 407868 374990 408326 375050
rect 408542 374990 408734 375050
rect 410014 374990 410094 375050
rect 407868 374988 407869 374990
rect 407803 374987 407869 374988
rect 408542 372605 408602 374990
rect 408539 372604 408605 372605
rect 408539 372540 408540 372604
rect 408604 372540 408605 372604
rect 408539 372539 408605 372540
rect 407251 371516 407317 371517
rect 407251 371452 407252 371516
rect 407316 371452 407317 371516
rect 407251 371451 407317 371452
rect 406147 371380 406213 371381
rect 406147 371316 406148 371380
rect 406212 371316 406213 371380
rect 406147 371315 406213 371316
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 355308 405854 370338
rect 408954 357554 409574 373000
rect 410014 372061 410074 374990
rect 410744 374645 410804 375020
rect 410741 374644 410807 374645
rect 410741 374580 410742 374644
rect 410806 374580 410807 374644
rect 410741 374579 410807 374580
rect 410011 372060 410077 372061
rect 410011 371996 410012 372060
rect 410076 371996 410077 372060
rect 410011 371995 410077 371996
rect 411302 371653 411362 375050
rect 411854 374990 412406 375050
rect 412774 374990 413494 375050
rect 413630 374990 413754 375050
rect 411299 371652 411365 371653
rect 411299 371588 411300 371652
rect 411364 371588 411365 371652
rect 411299 371587 411365 371588
rect 411854 371517 411914 374990
rect 411851 371516 411917 371517
rect 411851 371452 411852 371516
rect 411916 371452 411917 371516
rect 411851 371451 411917 371452
rect 412774 371381 412834 374990
rect 413694 371381 413754 374990
rect 414062 374990 414582 375050
rect 415534 374990 415942 375050
rect 416078 374990 416146 375050
rect 414062 371381 414122 374990
rect 415534 371381 415594 374990
rect 416086 373829 416146 374990
rect 416822 374990 417030 375050
rect 416083 373828 416149 373829
rect 416083 373764 416084 373828
rect 416148 373764 416149 373828
rect 416083 373763 416149 373764
rect 412771 371380 412837 371381
rect 412771 371316 412772 371380
rect 412836 371316 412837 371380
rect 412771 371315 412837 371316
rect 413691 371380 413757 371381
rect 413691 371316 413692 371380
rect 413756 371316 413757 371380
rect 413691 371315 413757 371316
rect 414059 371380 414125 371381
rect 414059 371316 414060 371380
rect 414124 371316 414125 371380
rect 414059 371315 414125 371316
rect 415531 371380 415597 371381
rect 415531 371316 415532 371380
rect 415596 371316 415597 371380
rect 415531 371315 415597 371316
rect 408954 357318 408986 357554
rect 409222 357318 409306 357554
rect 409542 357318 409574 357554
rect 408954 357234 409574 357318
rect 408954 356998 408986 357234
rect 409222 356998 409306 357234
rect 409542 356998 409574 357234
rect 408954 355308 409574 356998
rect 415794 364394 416414 373000
rect 416822 371381 416882 374990
rect 418110 371517 418170 375050
rect 418294 374990 418526 375050
rect 418846 374990 419478 375050
rect 420318 374990 420702 375050
rect 418107 371516 418173 371517
rect 418107 371452 418108 371516
rect 418172 371452 418173 371516
rect 418107 371451 418173 371452
rect 418294 371381 418354 374990
rect 418846 371653 418906 374990
rect 418843 371652 418909 371653
rect 418843 371588 418844 371652
rect 418908 371588 418909 371652
rect 418843 371587 418909 371588
rect 416819 371380 416885 371381
rect 416819 371316 416820 371380
rect 416884 371316 416885 371380
rect 416819 371315 416885 371316
rect 418291 371380 418357 371381
rect 418291 371316 418292 371380
rect 418356 371316 418357 371380
rect 418291 371315 418357 371316
rect 415794 364158 415826 364394
rect 416062 364158 416146 364394
rect 416382 364158 416414 364394
rect 415794 364074 416414 364158
rect 415794 363838 415826 364074
rect 416062 363838 416146 364074
rect 416382 363838 416414 364074
rect 415794 355308 416414 363838
rect 419514 366234 420134 373000
rect 420318 371381 420378 374990
rect 421054 373829 421114 375050
rect 421238 374990 421790 375050
rect 422342 374990 422878 375050
rect 423078 374990 423558 375050
rect 423966 374990 424058 375050
rect 421051 373828 421117 373829
rect 421051 373764 421052 373828
rect 421116 373764 421117 373828
rect 421051 373763 421117 373764
rect 421238 371517 421298 374990
rect 421235 371516 421301 371517
rect 421235 371452 421236 371516
rect 421300 371452 421301 371516
rect 421235 371451 421301 371452
rect 422342 371381 422402 374990
rect 423078 373829 423138 374990
rect 423075 373828 423141 373829
rect 423075 373764 423076 373828
rect 423140 373764 423141 373828
rect 423075 373763 423141 373764
rect 420315 371380 420381 371381
rect 420315 371316 420316 371380
rect 420380 371316 420381 371380
rect 420315 371315 420381 371316
rect 422339 371380 422405 371381
rect 422339 371316 422340 371380
rect 422404 371316 422405 371380
rect 422339 371315 422405 371316
rect 419514 365998 419546 366234
rect 419782 365998 419866 366234
rect 420102 365998 420134 366234
rect 419514 365914 420134 365998
rect 419514 365678 419546 365914
rect 419782 365678 419866 365914
rect 420102 365678 420134 365914
rect 419514 355308 420134 365678
rect 423234 369954 423854 373000
rect 423998 371653 424058 374990
rect 425099 374988 425100 375052
rect 425164 375050 425165 375052
rect 440371 375052 440437 375053
rect 425164 374990 425326 375050
rect 425654 374990 426006 375050
rect 425164 374988 425165 374990
rect 425099 374987 425165 374988
rect 423995 371652 424061 371653
rect 423995 371588 423996 371652
rect 424060 371588 424061 371652
rect 423995 371587 424061 371588
rect 425654 371381 425714 374990
rect 426390 372605 426450 375050
rect 426942 374990 427638 375050
rect 427862 374990 428318 375050
rect 428598 374990 428726 375050
rect 429150 374990 429814 375050
rect 430622 374990 431038 375050
rect 426942 373829 427002 374990
rect 426939 373828 427005 373829
rect 426939 373764 426940 373828
rect 427004 373764 427005 373828
rect 426939 373763 427005 373764
rect 426387 372604 426453 372605
rect 426387 372540 426388 372604
rect 426452 372540 426453 372604
rect 426387 372539 426453 372540
rect 425651 371380 425717 371381
rect 425651 371316 425652 371380
rect 425716 371316 425717 371380
rect 425651 371315 425717 371316
rect 423234 369718 423266 369954
rect 423502 369718 423586 369954
rect 423822 369718 423854 369954
rect 423234 369634 423854 369718
rect 423234 369398 423266 369634
rect 423502 369398 423586 369634
rect 423822 369398 423854 369634
rect 423234 355308 423854 369398
rect 426954 356614 427574 373000
rect 427862 371653 427922 374990
rect 427859 371652 427925 371653
rect 427859 371588 427860 371652
rect 427924 371588 427925 371652
rect 427859 371587 427925 371588
rect 428598 371381 428658 374990
rect 429150 374101 429210 374990
rect 429147 374100 429213 374101
rect 429147 374036 429148 374100
rect 429212 374036 429213 374100
rect 429147 374035 429213 374036
rect 430622 373829 430682 374990
rect 430619 373828 430685 373829
rect 430619 373764 430620 373828
rect 430684 373764 430685 373828
rect 430619 373763 430685 373764
rect 431174 372469 431234 375050
rect 432094 374990 432262 375050
rect 431171 372468 431237 372469
rect 431171 372404 431172 372468
rect 431236 372404 431237 372468
rect 431171 372403 431237 372404
rect 432094 371381 432154 374990
rect 433320 374370 433380 375020
rect 433592 374509 433652 375020
rect 433750 374990 434438 375050
rect 434854 374990 435798 375050
rect 433589 374508 433655 374509
rect 433589 374444 433590 374508
rect 433654 374444 433655 374508
rect 433589 374443 433655 374444
rect 433320 374310 433442 374370
rect 433382 371925 433442 374310
rect 433750 374010 433810 374990
rect 433566 373950 433810 374010
rect 433566 372605 433626 373950
rect 433563 372604 433629 372605
rect 433563 372540 433564 372604
rect 433628 372540 433629 372604
rect 433563 372539 433629 372540
rect 433379 371924 433445 371925
rect 433379 371860 433380 371924
rect 433444 371860 433445 371924
rect 433379 371859 433445 371860
rect 428595 371380 428661 371381
rect 428595 371316 428596 371380
rect 428660 371316 428661 371380
rect 428595 371315 428661 371316
rect 432091 371380 432157 371381
rect 432091 371316 432092 371380
rect 432156 371316 432157 371380
rect 432091 371315 432157 371316
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 355308 427574 356058
rect 433794 363454 434414 373000
rect 434854 371381 434914 374990
rect 436040 374509 436100 375020
rect 436326 374990 437022 375050
rect 438110 374990 438410 375050
rect 436037 374508 436103 374509
rect 436037 374444 436038 374508
rect 436102 374444 436103 374508
rect 436037 374443 436103 374444
rect 436326 371381 436386 374990
rect 434851 371380 434917 371381
rect 434851 371316 434852 371380
rect 434916 371316 434917 371380
rect 434851 371315 434917 371316
rect 436323 371380 436389 371381
rect 436323 371316 436324 371380
rect 436388 371316 436389 371380
rect 436323 371315 436389 371316
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 355308 434414 362898
rect 437514 367174 438134 373000
rect 438350 372605 438410 374990
rect 438488 374509 438548 375020
rect 439198 374990 439514 375050
rect 438485 374508 438551 374509
rect 438485 374444 438486 374508
rect 438550 374444 438551 374508
rect 438485 374443 438551 374444
rect 438347 372604 438413 372605
rect 438347 372540 438348 372604
rect 438412 372540 438413 372604
rect 438347 372539 438413 372540
rect 439454 371789 439514 374990
rect 440371 374988 440372 375052
rect 440436 375050 440437 375052
rect 443131 375052 443197 375053
rect 440436 374990 440966 375050
rect 440436 374988 440437 374990
rect 440371 374987 440437 374988
rect 443131 374988 443132 375052
rect 443196 375050 443197 375052
rect 443196 374990 443550 375050
rect 445894 374990 445998 375050
rect 447734 374990 448310 375050
rect 443196 374988 443197 374990
rect 443131 374987 443197 374988
rect 445894 373693 445954 374990
rect 445891 373692 445957 373693
rect 445891 373628 445892 373692
rect 445956 373628 445957 373692
rect 445891 373627 445957 373628
rect 447734 373557 447794 374990
rect 451000 374645 451060 375020
rect 452886 374990 453478 375050
rect 455462 374990 455926 375050
rect 458222 374990 458510 375050
rect 460958 374990 461042 375050
rect 450997 374644 451063 374645
rect 450997 374580 450998 374644
rect 451062 374580 451063 374644
rect 450997 374579 451063 374580
rect 447731 373556 447797 373557
rect 447731 373492 447732 373556
rect 447796 373492 447797 373556
rect 447731 373491 447797 373492
rect 452886 373421 452946 374990
rect 455462 373693 455522 374990
rect 455459 373692 455525 373693
rect 455459 373628 455460 373692
rect 455524 373628 455525 373692
rect 455459 373627 455525 373628
rect 458222 373557 458282 374990
rect 458219 373556 458285 373557
rect 458219 373492 458220 373556
rect 458284 373492 458285 373556
rect 458219 373491 458285 373492
rect 452883 373420 452949 373421
rect 452883 373356 452884 373420
rect 452948 373356 452949 373420
rect 452883 373355 452949 373356
rect 439451 371788 439517 371789
rect 439451 371724 439452 371788
rect 439516 371724 439517 371788
rect 439451 371723 439517 371724
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 355308 438134 366618
rect 441234 370894 441854 373000
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 355308 441854 370338
rect 444954 357554 445574 373000
rect 444954 357318 444986 357554
rect 445222 357318 445306 357554
rect 445542 357318 445574 357554
rect 444954 357234 445574 357318
rect 444954 356998 444986 357234
rect 445222 356998 445306 357234
rect 445542 356998 445574 357234
rect 444954 355308 445574 356998
rect 451794 364394 452414 373000
rect 451794 364158 451826 364394
rect 452062 364158 452146 364394
rect 452382 364158 452414 364394
rect 451794 364074 452414 364158
rect 451794 363838 451826 364074
rect 452062 363838 452146 364074
rect 452382 363838 452414 364074
rect 451794 355308 452414 363838
rect 455514 366234 456134 373000
rect 455514 365998 455546 366234
rect 455782 365998 455866 366234
rect 456102 365998 456134 366234
rect 455514 365914 456134 365998
rect 455514 365678 455546 365914
rect 455782 365678 455866 365914
rect 456102 365678 456134 365914
rect 455514 355308 456134 365678
rect 459234 369954 459854 373000
rect 460982 371381 461042 374990
rect 462638 374990 463542 375050
rect 465398 374990 465990 375050
rect 467974 374990 468574 375050
rect 470734 374990 471022 375050
rect 473310 374990 473470 375050
rect 475334 374990 475918 375050
rect 478094 374990 478502 375050
rect 480302 374990 480950 375050
rect 483246 374990 483398 375050
rect 485822 374990 485982 375050
rect 503118 374990 503254 375050
rect 503390 374990 503546 375050
rect 462638 371653 462698 374990
rect 462635 371652 462701 371653
rect 462635 371588 462636 371652
rect 462700 371588 462701 371652
rect 462635 371587 462701 371588
rect 460979 371380 461045 371381
rect 460979 371316 460980 371380
rect 461044 371316 461045 371380
rect 460979 371315 461045 371316
rect 459234 369718 459266 369954
rect 459502 369718 459586 369954
rect 459822 369718 459854 369954
rect 459234 369634 459854 369718
rect 459234 369398 459266 369634
rect 459502 369398 459586 369634
rect 459822 369398 459854 369634
rect 459234 355308 459854 369398
rect 462954 356614 463574 373000
rect 465398 371653 465458 374990
rect 465395 371652 465461 371653
rect 465395 371588 465396 371652
rect 465460 371588 465461 371652
rect 465395 371587 465461 371588
rect 467974 371381 468034 374990
rect 467971 371380 468037 371381
rect 467971 371316 467972 371380
rect 468036 371316 468037 371380
rect 467971 371315 468037 371316
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 355308 463574 356058
rect 469794 363454 470414 373000
rect 470734 372333 470794 374990
rect 470731 372332 470797 372333
rect 470731 372268 470732 372332
rect 470796 372268 470797 372332
rect 470731 372267 470797 372268
rect 473310 371381 473370 374990
rect 475334 373965 475394 374990
rect 475331 373964 475397 373965
rect 475331 373900 475332 373964
rect 475396 373900 475397 373964
rect 475331 373899 475397 373900
rect 473307 371380 473373 371381
rect 473307 371316 473308 371380
rect 473372 371316 473373 371380
rect 473307 371315 473373 371316
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 355308 470414 362898
rect 473514 367174 474134 373000
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 355308 474134 366618
rect 477234 370894 477854 373000
rect 478094 371653 478154 374990
rect 478091 371652 478157 371653
rect 478091 371588 478092 371652
rect 478156 371588 478157 371652
rect 478091 371587 478157 371588
rect 480302 371517 480362 374990
rect 480299 371516 480365 371517
rect 480299 371452 480300 371516
rect 480364 371452 480365 371516
rect 480299 371451 480365 371452
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 355308 477854 370338
rect 480954 357554 481574 373000
rect 483246 371381 483306 374990
rect 485822 373421 485882 374990
rect 485819 373420 485885 373421
rect 485819 373356 485820 373420
rect 485884 373356 485885 373420
rect 485819 373355 485885 373356
rect 483243 371380 483309 371381
rect 483243 371316 483244 371380
rect 483308 371316 483309 371380
rect 483243 371315 483309 371316
rect 480954 357318 480986 357554
rect 481222 357318 481306 357554
rect 481542 357318 481574 357554
rect 480954 357234 481574 357318
rect 480954 356998 480986 357234
rect 481222 356998 481306 357234
rect 481542 356998 481574 357234
rect 480954 355308 481574 356998
rect 487794 364394 488414 373000
rect 487794 364158 487826 364394
rect 488062 364158 488146 364394
rect 488382 364158 488414 364394
rect 487794 364074 488414 364158
rect 487794 363838 487826 364074
rect 488062 363838 488146 364074
rect 488382 363838 488414 364074
rect 487794 355308 488414 363838
rect 491514 366234 492134 373000
rect 491514 365998 491546 366234
rect 491782 365998 491866 366234
rect 492102 365998 492134 366234
rect 491514 365914 492134 365998
rect 491514 365678 491546 365914
rect 491782 365678 491866 365914
rect 492102 365678 492134 365914
rect 491514 355308 492134 365678
rect 495234 369954 495854 373000
rect 495234 369718 495266 369954
rect 495502 369718 495586 369954
rect 495822 369718 495854 369954
rect 495234 369634 495854 369718
rect 495234 369398 495266 369634
rect 495502 369398 495586 369634
rect 495822 369398 495854 369634
rect 495234 355308 495854 369398
rect 498954 356614 499574 373000
rect 503118 372197 503178 374990
rect 503486 372197 503546 374990
rect 503115 372196 503181 372197
rect 503115 372132 503116 372196
rect 503180 372132 503181 372196
rect 503115 372131 503181 372132
rect 503483 372196 503549 372197
rect 503483 372132 503484 372196
rect 503548 372132 503549 372196
rect 503483 372131 503549 372132
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 355308 499574 356058
rect 505794 363454 506414 373000
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 355308 506414 362898
rect 509514 367174 510134 373000
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 355308 510134 366618
rect 513234 370894 513854 373000
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 355308 513854 370338
rect 516954 357554 517574 373000
rect 516954 357318 516986 357554
rect 517222 357318 517306 357554
rect 517542 357318 517574 357554
rect 516954 357234 517574 357318
rect 516954 356998 516986 357234
rect 517222 356998 517306 357234
rect 517542 356998 517574 357234
rect 516954 355308 517574 356998
rect 498515 355060 498581 355061
rect 498515 354996 498516 355060
rect 498580 354996 498581 355060
rect 498515 354995 498581 354996
rect 498518 353970 498578 354995
rect 499803 354924 499869 354925
rect 499803 354860 499804 354924
rect 499868 354860 499869 354924
rect 499803 354859 499869 354860
rect 499806 353970 499866 354859
rect 510843 354788 510909 354789
rect 510843 354724 510844 354788
rect 510908 354724 510909 354788
rect 510843 354723 510909 354724
rect 510846 353970 510906 354723
rect 498464 353910 498578 353970
rect 499688 353910 499866 353970
rect 510840 353910 510906 353970
rect 498464 353260 498524 353910
rect 499688 353260 499748 353910
rect 510840 353260 510900 353910
rect 380272 345454 380620 345486
rect 380272 345218 380328 345454
rect 380564 345218 380620 345454
rect 380272 345134 380620 345218
rect 380272 344898 380328 345134
rect 380564 344898 380620 345134
rect 380272 344866 380620 344898
rect 516000 345454 516348 345486
rect 516000 345218 516056 345454
rect 516292 345218 516348 345454
rect 516000 345134 516348 345218
rect 516000 344898 516056 345134
rect 516292 344898 516348 345134
rect 516000 344866 516348 344898
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 380952 327454 381300 327486
rect 380952 327218 381008 327454
rect 381244 327218 381300 327454
rect 380952 327134 381300 327218
rect 380952 326898 381008 327134
rect 381244 326898 381300 327134
rect 380952 326866 381300 326898
rect 515320 327454 515668 327486
rect 515320 327218 515376 327454
rect 515612 327218 515668 327454
rect 515320 327134 515668 327218
rect 515320 326898 515376 327134
rect 515612 326898 515668 327134
rect 515320 326866 515668 326898
rect 380272 309454 380620 309486
rect 380272 309218 380328 309454
rect 380564 309218 380620 309454
rect 380272 309134 380620 309218
rect 380272 308898 380328 309134
rect 380564 308898 380620 309134
rect 380272 308866 380620 308898
rect 516000 309454 516348 309486
rect 516000 309218 516056 309454
rect 516292 309218 516348 309454
rect 516000 309134 516348 309218
rect 516000 308898 516056 309134
rect 516292 308898 516348 309134
rect 516000 308866 516348 308898
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 380952 291454 381300 291486
rect 380952 291218 381008 291454
rect 381244 291218 381300 291454
rect 380952 291134 381300 291218
rect 380952 290898 381008 291134
rect 381244 290898 381300 291134
rect 380952 290866 381300 290898
rect 515320 291454 515668 291486
rect 515320 291218 515376 291454
rect 515612 291218 515668 291454
rect 515320 291134 515668 291218
rect 515320 290898 515376 291134
rect 515612 290898 515668 291134
rect 515320 290866 515668 290898
rect 380272 273454 380620 273486
rect 380272 273218 380328 273454
rect 380564 273218 380620 273454
rect 380272 273134 380620 273218
rect 380272 272898 380328 273134
rect 380564 272898 380620 273134
rect 380272 272866 380620 272898
rect 516000 273454 516348 273486
rect 516000 273218 516056 273454
rect 516292 273218 516348 273454
rect 516000 273134 516348 273218
rect 516000 272898 516056 273134
rect 516292 272898 516348 273134
rect 516000 272866 516348 272898
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 396056 269650 396116 270106
rect 397144 269650 397204 270106
rect 396030 269590 396116 269650
rect 397134 269590 397204 269650
rect 398232 269650 398292 270106
rect 399592 269650 399652 270106
rect 400544 269650 400604 270106
rect 401768 269650 401828 270106
rect 403128 269650 403188 270106
rect 404216 269650 404276 270106
rect 405440 269650 405500 270106
rect 406528 269650 406588 270106
rect 398232 269590 398298 269650
rect 379470 267690 379714 267750
rect 379470 267477 379530 267690
rect 379467 267476 379533 267477
rect 379467 267412 379468 267476
rect 379532 267412 379533 267476
rect 379467 267411 379533 267412
rect 379794 256394 380414 268000
rect 379794 256158 379826 256394
rect 380062 256158 380146 256394
rect 380382 256158 380414 256394
rect 379794 256074 380414 256158
rect 379794 255838 379826 256074
rect 380062 255838 380146 256074
rect 380382 255838 380414 256074
rect 379794 250308 380414 255838
rect 383514 260114 384134 268000
rect 383514 259878 383546 260114
rect 383782 259878 383866 260114
rect 384102 259878 384134 260114
rect 383514 259794 384134 259878
rect 383514 259558 383546 259794
rect 383782 259558 383866 259794
rect 384102 259558 384134 259794
rect 383514 250308 384134 259558
rect 387234 261954 387854 268000
rect 387234 261718 387266 261954
rect 387502 261718 387586 261954
rect 387822 261718 387854 261954
rect 387234 261634 387854 261718
rect 387234 261398 387266 261634
rect 387502 261398 387586 261634
rect 387822 261398 387854 261634
rect 387234 250308 387854 261398
rect 390954 265674 391574 268000
rect 396030 266389 396090 269590
rect 397134 267205 397194 269590
rect 398238 268157 398298 269590
rect 399526 269590 399652 269650
rect 400446 269590 400604 269650
rect 401734 269590 401828 269650
rect 403022 269590 403188 269650
rect 404126 269590 404276 269650
rect 405046 269590 405500 269650
rect 406518 269590 406588 269650
rect 407616 269650 407676 270106
rect 408296 269650 408356 270106
rect 407616 269590 407682 269650
rect 398235 268156 398301 268157
rect 398235 268092 398236 268156
rect 398300 268092 398301 268156
rect 398235 268091 398301 268092
rect 397131 267204 397197 267205
rect 397131 267140 397132 267204
rect 397196 267140 397197 267204
rect 397131 267139 397197 267140
rect 396027 266388 396093 266389
rect 396027 266324 396028 266388
rect 396092 266324 396093 266388
rect 396027 266323 396093 266324
rect 390954 265438 390986 265674
rect 391222 265438 391306 265674
rect 391542 265438 391574 265674
rect 390954 265354 391574 265438
rect 390954 265118 390986 265354
rect 391222 265118 391306 265354
rect 391542 265118 391574 265354
rect 390954 250308 391574 265118
rect 397794 255454 398414 268000
rect 399526 266389 399586 269590
rect 400446 266389 400506 269590
rect 401734 268157 401794 269590
rect 401731 268156 401797 268157
rect 401731 268092 401732 268156
rect 401796 268092 401797 268156
rect 401731 268091 401797 268092
rect 399523 266388 399589 266389
rect 399523 266324 399524 266388
rect 399588 266324 399589 266388
rect 399523 266323 399589 266324
rect 400443 266388 400509 266389
rect 400443 266324 400444 266388
rect 400508 266324 400509 266388
rect 400443 266323 400509 266324
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 250308 398414 254898
rect 401514 259174 402134 268000
rect 403022 267749 403082 269590
rect 403019 267748 403085 267749
rect 403019 267684 403020 267748
rect 403084 267684 403085 267748
rect 403019 267683 403085 267684
rect 404126 266389 404186 269590
rect 405046 266389 405106 269590
rect 404123 266388 404189 266389
rect 404123 266324 404124 266388
rect 404188 266324 404189 266388
rect 404123 266323 404189 266324
rect 405043 266388 405109 266389
rect 405043 266324 405044 266388
rect 405108 266324 405109 266388
rect 405043 266323 405109 266324
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 250308 402134 258618
rect 405234 262894 405854 268000
rect 406518 266389 406578 269590
rect 407622 266389 407682 269590
rect 408174 269590 408356 269650
rect 408704 269650 408764 270106
rect 410064 269650 410124 270106
rect 408704 269590 408786 269650
rect 408174 267341 408234 269590
rect 408171 267340 408237 267341
rect 408171 267276 408172 267340
rect 408236 267276 408237 267340
rect 408171 267275 408237 267276
rect 408726 266661 408786 269590
rect 410014 269590 410124 269650
rect 410744 269650 410804 270106
rect 411288 269650 411348 270106
rect 412376 269650 412436 270106
rect 413464 269650 413524 270106
rect 410744 269590 410810 269650
rect 411288 269590 411362 269650
rect 412376 269590 412466 269650
rect 408723 266660 408789 266661
rect 408723 266596 408724 266660
rect 408788 266596 408789 266660
rect 408723 266595 408789 266596
rect 408954 266614 409574 268000
rect 406515 266388 406581 266389
rect 406515 266324 406516 266388
rect 406580 266324 406581 266388
rect 406515 266323 406581 266324
rect 407619 266388 407685 266389
rect 407619 266324 407620 266388
rect 407684 266324 407685 266388
rect 407619 266323 407685 266324
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 410014 266389 410074 269590
rect 410750 267069 410810 269590
rect 410747 267068 410813 267069
rect 410747 267004 410748 267068
rect 410812 267004 410813 267068
rect 410747 267003 410813 267004
rect 411302 266389 411362 269590
rect 412406 266525 412466 269590
rect 413326 269590 413524 269650
rect 413600 269650 413660 270106
rect 414552 269650 414612 270106
rect 415912 269650 415972 270106
rect 416048 269789 416108 270106
rect 416045 269788 416111 269789
rect 416045 269724 416046 269788
rect 416110 269724 416111 269788
rect 416045 269723 416111 269724
rect 413600 269590 413754 269650
rect 412403 266524 412469 266525
rect 412403 266460 412404 266524
rect 412468 266460 412469 266524
rect 412403 266459 412469 266460
rect 413326 266389 413386 269590
rect 413694 267069 413754 269590
rect 414430 269590 414612 269650
rect 415534 269590 415972 269650
rect 417000 269650 417060 270106
rect 418088 269650 418148 270106
rect 418496 269650 418556 270106
rect 419448 269650 419508 270106
rect 417000 269590 417066 269650
rect 418088 269590 418170 269650
rect 414430 267749 414490 269590
rect 415534 267749 415594 269590
rect 417006 268837 417066 269590
rect 417003 268836 417069 268837
rect 417003 268772 417004 268836
rect 417068 268772 417069 268836
rect 417003 268771 417069 268772
rect 414427 267748 414493 267749
rect 414427 267684 414428 267748
rect 414492 267684 414493 267748
rect 414427 267683 414493 267684
rect 415531 267748 415597 267749
rect 415531 267684 415532 267748
rect 415596 267684 415597 267748
rect 415531 267683 415597 267684
rect 413691 267068 413757 267069
rect 413691 267004 413692 267068
rect 413756 267004 413757 267068
rect 413691 267003 413757 267004
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 250308 405854 262338
rect 408954 266294 409574 266378
rect 410011 266388 410077 266389
rect 410011 266324 410012 266388
rect 410076 266324 410077 266388
rect 410011 266323 410077 266324
rect 411299 266388 411365 266389
rect 411299 266324 411300 266388
rect 411364 266324 411365 266388
rect 411299 266323 411365 266324
rect 413323 266388 413389 266389
rect 413323 266324 413324 266388
rect 413388 266324 413389 266388
rect 413323 266323 413389 266324
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 250308 409574 266058
rect 415794 256394 416414 268000
rect 418110 266389 418170 269590
rect 418478 269590 418556 269650
rect 419214 269590 419508 269650
rect 420672 269650 420732 270106
rect 421080 269650 421140 270106
rect 420672 269590 420746 269650
rect 418478 267205 418538 269590
rect 418475 267204 418541 267205
rect 418475 267140 418476 267204
rect 418540 267140 418541 267204
rect 418475 267139 418541 267140
rect 419214 266525 419274 269590
rect 419211 266524 419277 266525
rect 419211 266460 419212 266524
rect 419276 266460 419277 266524
rect 419211 266459 419277 266460
rect 418107 266388 418173 266389
rect 418107 266324 418108 266388
rect 418172 266324 418173 266388
rect 418107 266323 418173 266324
rect 415794 256158 415826 256394
rect 416062 256158 416146 256394
rect 416382 256158 416414 256394
rect 415794 256074 416414 256158
rect 415794 255838 415826 256074
rect 416062 255838 416146 256074
rect 416382 255838 416414 256074
rect 415794 250308 416414 255838
rect 419514 260114 420134 268000
rect 420686 266389 420746 269590
rect 421054 269590 421140 269650
rect 421760 269650 421820 270106
rect 422848 269650 422908 270106
rect 423528 269650 423588 270106
rect 421760 269590 421850 269650
rect 422848 269590 422954 269650
rect 421054 268837 421114 269590
rect 421051 268836 421117 268837
rect 421051 268772 421052 268836
rect 421116 268772 421117 268836
rect 421051 268771 421117 268772
rect 421790 266389 421850 269590
rect 422894 268973 422954 269590
rect 423446 269590 423588 269650
rect 423936 269650 423996 270106
rect 425296 269789 425356 270106
rect 425293 269788 425359 269789
rect 425293 269724 425294 269788
rect 425358 269724 425359 269788
rect 425293 269723 425359 269724
rect 425976 269650 426036 270106
rect 426384 269650 426444 270106
rect 427608 269650 427668 270106
rect 428288 269650 428348 270106
rect 428696 269650 428756 270106
rect 429784 269653 429844 270106
rect 423936 269590 424058 269650
rect 425976 269590 426082 269650
rect 426384 269590 426450 269650
rect 427608 269590 427738 269650
rect 422891 268972 422957 268973
rect 422891 268908 422892 268972
rect 422956 268908 422957 268972
rect 422891 268907 422957 268908
rect 423446 268837 423506 269590
rect 423443 268836 423509 268837
rect 423443 268772 423444 268836
rect 423508 268772 423509 268836
rect 423443 268771 423509 268772
rect 423998 268701 424058 269590
rect 426022 268973 426082 269590
rect 426019 268972 426085 268973
rect 426019 268908 426020 268972
rect 426084 268908 426085 268972
rect 426019 268907 426085 268908
rect 423995 268700 424061 268701
rect 423995 268636 423996 268700
rect 424060 268636 424061 268700
rect 423995 268635 424061 268636
rect 420683 266388 420749 266389
rect 420683 266324 420684 266388
rect 420748 266324 420749 266388
rect 420683 266323 420749 266324
rect 421787 266388 421853 266389
rect 421787 266324 421788 266388
rect 421852 266324 421853 266388
rect 421787 266323 421853 266324
rect 419514 259878 419546 260114
rect 419782 259878 419866 260114
rect 420102 259878 420134 260114
rect 419514 259794 420134 259878
rect 419514 259558 419546 259794
rect 419782 259558 419866 259794
rect 420102 259558 420134 259794
rect 419514 250308 420134 259558
rect 423234 261954 423854 268000
rect 426390 265709 426450 269590
rect 426387 265708 426453 265709
rect 426387 265644 426388 265708
rect 426452 265644 426453 265708
rect 426387 265643 426453 265644
rect 426954 265674 427574 268000
rect 427678 266389 427738 269590
rect 428230 269590 428348 269650
rect 428598 269590 428756 269650
rect 429781 269652 429847 269653
rect 428230 267477 428290 269590
rect 428598 267749 428658 269590
rect 429781 269588 429782 269652
rect 429846 269588 429847 269652
rect 431008 269650 431068 270106
rect 429781 269587 429847 269588
rect 430990 269590 431068 269650
rect 431144 269650 431204 270106
rect 432232 269650 432292 270106
rect 433320 269789 433380 270106
rect 433317 269788 433383 269789
rect 433317 269724 433318 269788
rect 433382 269724 433383 269788
rect 433317 269723 433383 269724
rect 433592 269650 433652 270106
rect 434408 269789 434468 270106
rect 434405 269788 434471 269789
rect 434405 269724 434406 269788
rect 434470 269724 434471 269788
rect 434405 269723 434471 269724
rect 435768 269650 435828 270106
rect 436040 269653 436100 270106
rect 431144 269590 431234 269650
rect 432232 269590 432338 269650
rect 430990 268973 431050 269590
rect 430987 268972 431053 268973
rect 430987 268908 430988 268972
rect 431052 268908 431053 268972
rect 430987 268907 431053 268908
rect 428595 267748 428661 267749
rect 428595 267684 428596 267748
rect 428660 267684 428661 267748
rect 428595 267683 428661 267684
rect 428227 267476 428293 267477
rect 428227 267412 428228 267476
rect 428292 267412 428293 267476
rect 428227 267411 428293 267412
rect 427675 266388 427741 266389
rect 427675 266324 427676 266388
rect 427740 266324 427741 266388
rect 427675 266323 427741 266324
rect 423234 261718 423266 261954
rect 423502 261718 423586 261954
rect 423822 261718 423854 261954
rect 423234 261634 423854 261718
rect 423234 261398 423266 261634
rect 423502 261398 423586 261634
rect 423822 261398 423854 261634
rect 423234 250308 423854 261398
rect 426954 265438 426986 265674
rect 427222 265438 427306 265674
rect 427542 265438 427574 265674
rect 431174 265573 431234 269590
rect 432278 268973 432338 269590
rect 433566 269590 433652 269650
rect 435590 269590 435828 269650
rect 436037 269652 436103 269653
rect 432275 268972 432341 268973
rect 432275 268908 432276 268972
rect 432340 268908 432341 268972
rect 432275 268907 432341 268908
rect 433566 267069 433626 269590
rect 433563 267068 433629 267069
rect 433563 267004 433564 267068
rect 433628 267004 433629 267068
rect 433563 267003 433629 267004
rect 431171 265572 431237 265573
rect 431171 265508 431172 265572
rect 431236 265508 431237 265572
rect 431171 265507 431237 265508
rect 426954 265354 427574 265438
rect 426954 265118 426986 265354
rect 427222 265118 427306 265354
rect 427542 265118 427574 265354
rect 426954 250308 427574 265118
rect 433794 255454 434414 268000
rect 435590 267749 435650 269590
rect 436037 269588 436038 269652
rect 436102 269588 436103 269652
rect 436992 269650 437052 270106
rect 436037 269587 436103 269588
rect 436878 269590 437052 269650
rect 438080 269650 438140 270106
rect 438488 269650 438548 270106
rect 439168 269650 439228 270106
rect 440936 269650 440996 270106
rect 443520 269650 443580 270106
rect 445968 269650 446028 270106
rect 438080 269590 438410 269650
rect 438488 269590 438594 269650
rect 439168 269590 439330 269650
rect 435587 267748 435653 267749
rect 435587 267684 435588 267748
rect 435652 267684 435653 267748
rect 435587 267683 435653 267684
rect 436878 266389 436938 269590
rect 436875 266388 436941 266389
rect 436875 266324 436876 266388
rect 436940 266324 436941 266388
rect 436875 266323 436941 266324
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 250308 434414 254898
rect 437514 259174 438134 268000
rect 438350 266661 438410 269590
rect 438534 267205 438594 269590
rect 439270 267341 439330 269590
rect 440926 269590 440996 269650
rect 443502 269590 443580 269650
rect 445894 269590 446028 269650
rect 448280 269650 448340 270106
rect 451000 269650 451060 270106
rect 453448 269650 453508 270106
rect 455896 269650 455956 270106
rect 458480 269650 458540 270106
rect 448280 269590 448346 269650
rect 451000 269590 451106 269650
rect 440926 267341 440986 269590
rect 439267 267340 439333 267341
rect 439267 267276 439268 267340
rect 439332 267276 439333 267340
rect 439267 267275 439333 267276
rect 440923 267340 440989 267341
rect 440923 267276 440924 267340
rect 440988 267276 440989 267340
rect 440923 267275 440989 267276
rect 438531 267204 438597 267205
rect 438531 267140 438532 267204
rect 438596 267140 438597 267204
rect 438531 267139 438597 267140
rect 438347 266660 438413 266661
rect 438347 266596 438348 266660
rect 438412 266596 438413 266660
rect 438347 266595 438413 266596
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 250308 438134 258618
rect 441234 262894 441854 268000
rect 443502 267477 443562 269590
rect 443499 267476 443565 267477
rect 443499 267412 443500 267476
rect 443564 267412 443565 267476
rect 443499 267411 443565 267412
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 250308 441854 262338
rect 444954 266614 445574 268000
rect 445894 267205 445954 269590
rect 448286 267341 448346 269590
rect 451046 267749 451106 269590
rect 453438 269590 453508 269650
rect 455830 269590 455956 269650
rect 458406 269590 458540 269650
rect 460928 269650 460988 270106
rect 463512 269650 463572 270106
rect 465960 269650 466020 270106
rect 468544 269653 468604 270106
rect 470992 269653 471052 270106
rect 460928 269590 461042 269650
rect 463512 269590 463618 269650
rect 451043 267748 451109 267749
rect 451043 267684 451044 267748
rect 451108 267684 451109 267748
rect 451043 267683 451109 267684
rect 448283 267340 448349 267341
rect 448283 267276 448284 267340
rect 448348 267276 448349 267340
rect 448283 267275 448349 267276
rect 445891 267204 445957 267205
rect 445891 267140 445892 267204
rect 445956 267140 445957 267204
rect 445891 267139 445957 267140
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 250308 445574 266058
rect 451794 256394 452414 268000
rect 453438 267749 453498 269590
rect 455830 268157 455890 269590
rect 455827 268156 455893 268157
rect 455827 268092 455828 268156
rect 455892 268092 455893 268156
rect 455827 268091 455893 268092
rect 453435 267748 453501 267749
rect 453435 267684 453436 267748
rect 453500 267684 453501 267748
rect 453435 267683 453501 267684
rect 451794 256158 451826 256394
rect 452062 256158 452146 256394
rect 452382 256158 452414 256394
rect 451794 256074 452414 256158
rect 451794 255838 451826 256074
rect 452062 255838 452146 256074
rect 452382 255838 452414 256074
rect 451794 250308 452414 255838
rect 455514 260114 456134 268000
rect 458406 267749 458466 269590
rect 458403 267748 458469 267749
rect 458403 267684 458404 267748
rect 458468 267684 458469 267748
rect 458403 267683 458469 267684
rect 455514 259878 455546 260114
rect 455782 259878 455866 260114
rect 456102 259878 456134 260114
rect 455514 259794 456134 259878
rect 455514 259558 455546 259794
rect 455782 259558 455866 259794
rect 456102 259558 456134 259794
rect 455514 250308 456134 259558
rect 459234 261954 459854 268000
rect 460982 267749 461042 269590
rect 463558 268157 463618 269590
rect 465950 269590 466020 269650
rect 468541 269652 468607 269653
rect 463555 268156 463621 268157
rect 463555 268092 463556 268156
rect 463620 268092 463621 268156
rect 463555 268091 463621 268092
rect 460979 267748 461045 267749
rect 460979 267684 460980 267748
rect 461044 267684 461045 267748
rect 460979 267683 461045 267684
rect 459234 261718 459266 261954
rect 459502 261718 459586 261954
rect 459822 261718 459854 261954
rect 459234 261634 459854 261718
rect 459234 261398 459266 261634
rect 459502 261398 459586 261634
rect 459822 261398 459854 261634
rect 459234 250308 459854 261398
rect 462954 265674 463574 268000
rect 465950 266933 466010 269590
rect 468541 269588 468542 269652
rect 468606 269588 468607 269652
rect 468541 269587 468607 269588
rect 470989 269652 471055 269653
rect 470989 269588 470990 269652
rect 471054 269588 471055 269652
rect 473440 269650 473500 270106
rect 475888 269650 475948 270106
rect 478472 269650 478532 270106
rect 480920 269653 480980 270106
rect 473440 269590 473554 269650
rect 470989 269587 471055 269588
rect 473494 269245 473554 269590
rect 475886 269590 475948 269650
rect 478462 269590 478532 269650
rect 480917 269652 480983 269653
rect 473491 269244 473557 269245
rect 473491 269180 473492 269244
rect 473556 269180 473557 269244
rect 473491 269179 473557 269180
rect 475886 268973 475946 269590
rect 478462 268973 478522 269590
rect 480917 269588 480918 269652
rect 480982 269588 480983 269652
rect 483368 269650 483428 270106
rect 485952 269650 486012 270106
rect 503224 269650 503284 270106
rect 483368 269590 483490 269650
rect 485952 269590 486066 269650
rect 480917 269587 480983 269588
rect 483430 268973 483490 269590
rect 486006 269109 486066 269590
rect 503118 269590 503284 269650
rect 503360 269650 503420 270106
rect 503360 269590 503546 269650
rect 486003 269108 486069 269109
rect 486003 269044 486004 269108
rect 486068 269044 486069 269108
rect 486003 269043 486069 269044
rect 475883 268972 475949 268973
rect 475883 268908 475884 268972
rect 475948 268908 475949 268972
rect 475883 268907 475949 268908
rect 478459 268972 478525 268973
rect 478459 268908 478460 268972
rect 478524 268908 478525 268972
rect 478459 268907 478525 268908
rect 483427 268972 483493 268973
rect 483427 268908 483428 268972
rect 483492 268908 483493 268972
rect 483427 268907 483493 268908
rect 465947 266932 466013 266933
rect 465947 266868 465948 266932
rect 466012 266868 466013 266932
rect 465947 266867 466013 266868
rect 462954 265438 462986 265674
rect 463222 265438 463306 265674
rect 463542 265438 463574 265674
rect 462954 265354 463574 265438
rect 462954 265118 462986 265354
rect 463222 265118 463306 265354
rect 463542 265118 463574 265354
rect 462954 250308 463574 265118
rect 469794 255454 470414 268000
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 250308 470414 254898
rect 473514 259174 474134 268000
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 250308 474134 258618
rect 477234 262894 477854 268000
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 250308 477854 262338
rect 480954 266614 481574 268000
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 250308 481574 266058
rect 487794 256394 488414 268000
rect 487794 256158 487826 256394
rect 488062 256158 488146 256394
rect 488382 256158 488414 256394
rect 487794 256074 488414 256158
rect 487794 255838 487826 256074
rect 488062 255838 488146 256074
rect 488382 255838 488414 256074
rect 487794 250308 488414 255838
rect 491514 260114 492134 268000
rect 491514 259878 491546 260114
rect 491782 259878 491866 260114
rect 492102 259878 492134 260114
rect 491514 259794 492134 259878
rect 491514 259558 491546 259794
rect 491782 259558 491866 259794
rect 492102 259558 492134 259794
rect 491514 250308 492134 259558
rect 495234 261954 495854 268000
rect 495234 261718 495266 261954
rect 495502 261718 495586 261954
rect 495822 261718 495854 261954
rect 495234 261634 495854 261718
rect 495234 261398 495266 261634
rect 495502 261398 495586 261634
rect 495822 261398 495854 261634
rect 495234 250308 495854 261398
rect 498954 265674 499574 268000
rect 503118 267477 503178 269590
rect 503486 267477 503546 269590
rect 503115 267476 503181 267477
rect 503115 267412 503116 267476
rect 503180 267412 503181 267476
rect 503115 267411 503181 267412
rect 503483 267476 503549 267477
rect 503483 267412 503484 267476
rect 503548 267412 503549 267476
rect 503483 267411 503549 267412
rect 498954 265438 498986 265674
rect 499222 265438 499306 265674
rect 499542 265438 499574 265674
rect 498954 265354 499574 265438
rect 498954 265118 498986 265354
rect 499222 265118 499306 265354
rect 499542 265118 499574 265354
rect 498954 250308 499574 265118
rect 505794 255454 506414 268000
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 250308 506414 254898
rect 509514 259174 510134 268000
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 250308 510134 258618
rect 513234 262894 513854 268000
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 250308 513854 262338
rect 516954 266614 517574 268000
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 250308 517574 266058
rect 498515 249932 498581 249933
rect 498515 249868 498516 249932
rect 498580 249868 498581 249932
rect 498515 249867 498581 249868
rect 499803 249932 499869 249933
rect 499803 249868 499804 249932
rect 499868 249868 499869 249932
rect 499803 249867 499869 249868
rect 510843 249932 510909 249933
rect 510843 249868 510844 249932
rect 510908 249868 510909 249932
rect 510843 249867 510909 249868
rect 498518 248430 498578 249867
rect 499806 248430 499866 249867
rect 510846 248430 510906 249867
rect 498464 248370 498578 248430
rect 499688 248370 499866 248430
rect 510840 248370 510906 248430
rect 498464 248202 498524 248370
rect 499688 248202 499748 248370
rect 510840 248202 510900 248370
rect 380272 237454 380620 237486
rect 380272 237218 380328 237454
rect 380564 237218 380620 237454
rect 380272 237134 380620 237218
rect 380272 236898 380328 237134
rect 380564 236898 380620 237134
rect 380272 236866 380620 236898
rect 516000 237454 516348 237486
rect 516000 237218 516056 237454
rect 516292 237218 516348 237454
rect 516000 237134 516348 237218
rect 516000 236898 516056 237134
rect 516292 236898 516348 237134
rect 516000 236866 516348 236898
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 380952 219454 381300 219486
rect 380952 219218 381008 219454
rect 381244 219218 381300 219454
rect 380952 219134 381300 219218
rect 380952 218898 381008 219134
rect 381244 218898 381300 219134
rect 380952 218866 381300 218898
rect 515320 219454 515668 219486
rect 515320 219218 515376 219454
rect 515612 219218 515668 219454
rect 515320 219134 515668 219218
rect 515320 218898 515376 219134
rect 515612 218898 515668 219134
rect 515320 218866 515668 218898
rect 380272 201454 380620 201486
rect 380272 201218 380328 201454
rect 380564 201218 380620 201454
rect 380272 201134 380620 201218
rect 380272 200898 380328 201134
rect 380564 200898 380620 201134
rect 380272 200866 380620 200898
rect 516000 201454 516348 201486
rect 516000 201218 516056 201454
rect 516292 201218 516348 201454
rect 516000 201134 516348 201218
rect 516000 200898 516056 201134
rect 516292 200898 516348 201134
rect 516000 200866 516348 200898
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 380952 183454 381300 183486
rect 380952 183218 381008 183454
rect 381244 183218 381300 183454
rect 380952 183134 381300 183218
rect 380952 182898 381008 183134
rect 381244 182898 381300 183134
rect 380952 182866 381300 182898
rect 515320 183454 515668 183486
rect 515320 183218 515376 183454
rect 515612 183218 515668 183454
rect 515320 183134 515668 183218
rect 515320 182898 515376 183134
rect 515612 182898 515668 183134
rect 515320 182866 515668 182898
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 396056 164930 396116 165106
rect 397144 164930 397204 165106
rect 396030 164870 396116 164930
rect 397134 164870 397204 164930
rect 398232 164930 398292 165106
rect 399592 164930 399652 165106
rect 400544 164930 400604 165106
rect 401768 164930 401828 165106
rect 403128 164930 403188 165106
rect 404216 164930 404276 165106
rect 405440 164930 405500 165106
rect 406528 164930 406588 165106
rect 398232 164870 398298 164930
rect 379467 148476 379533 148477
rect 379467 148412 379468 148476
rect 379532 148412 379533 148476
rect 379467 148411 379533 148412
rect 379470 142170 379530 148411
rect 379794 148394 380414 163000
rect 379794 148158 379826 148394
rect 380062 148158 380146 148394
rect 380382 148158 380414 148394
rect 379794 148074 380414 148158
rect 379794 147838 379826 148074
rect 380062 147838 380146 148074
rect 380382 147838 380414 148074
rect 379794 145308 380414 147838
rect 383514 152114 384134 163000
rect 383514 151878 383546 152114
rect 383782 151878 383866 152114
rect 384102 151878 384134 152114
rect 383514 151794 384134 151878
rect 383514 151558 383546 151794
rect 383782 151558 383866 151794
rect 384102 151558 384134 151794
rect 383514 145308 384134 151558
rect 387234 153954 387854 163000
rect 387234 153718 387266 153954
rect 387502 153718 387586 153954
rect 387822 153718 387854 153954
rect 387234 153634 387854 153718
rect 387234 153398 387266 153634
rect 387502 153398 387586 153634
rect 387822 153398 387854 153634
rect 387234 145308 387854 153398
rect 390954 157674 391574 163000
rect 396030 162757 396090 164870
rect 396027 162756 396093 162757
rect 396027 162692 396028 162756
rect 396092 162692 396093 162756
rect 396027 162691 396093 162692
rect 397134 162213 397194 164870
rect 398238 163165 398298 164870
rect 399526 164870 399652 164930
rect 400446 164870 400604 164930
rect 401734 164870 401828 164930
rect 403022 164870 403188 164930
rect 404126 164870 404276 164930
rect 405046 164870 405500 164930
rect 406518 164870 406588 164930
rect 407616 164930 407676 165106
rect 408296 164930 408356 165106
rect 408704 164930 408764 165106
rect 410064 164930 410124 165106
rect 407616 164870 407682 164930
rect 408296 164870 408418 164930
rect 408704 164870 408786 164930
rect 398235 163164 398301 163165
rect 398235 163100 398236 163164
rect 398300 163100 398301 163164
rect 398235 163099 398301 163100
rect 397131 162212 397197 162213
rect 397131 162148 397132 162212
rect 397196 162148 397197 162212
rect 397131 162147 397197 162148
rect 390954 157438 390986 157674
rect 391222 157438 391306 157674
rect 391542 157438 391574 157674
rect 390954 157354 391574 157438
rect 390954 157118 390986 157354
rect 391222 157118 391306 157354
rect 391542 157118 391574 157354
rect 390954 145308 391574 157118
rect 397794 147454 398414 163000
rect 399526 162757 399586 164870
rect 400446 162757 400506 164870
rect 401734 163165 401794 164870
rect 401731 163164 401797 163165
rect 401731 163100 401732 163164
rect 401796 163100 401797 163164
rect 401731 163099 401797 163100
rect 399523 162756 399589 162757
rect 399523 162692 399524 162756
rect 399588 162692 399589 162756
rect 399523 162691 399589 162692
rect 400443 162756 400509 162757
rect 400443 162692 400444 162756
rect 400508 162692 400509 162756
rect 400443 162691 400509 162692
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 145308 398414 146898
rect 401514 151174 402134 163000
rect 403022 162757 403082 164870
rect 403019 162756 403085 162757
rect 403019 162692 403020 162756
rect 403084 162692 403085 162756
rect 403019 162691 403085 162692
rect 404126 162213 404186 164870
rect 405046 162757 405106 164870
rect 405043 162756 405109 162757
rect 405043 162692 405044 162756
rect 405108 162692 405109 162756
rect 405043 162691 405109 162692
rect 404123 162212 404189 162213
rect 404123 162148 404124 162212
rect 404188 162148 404189 162212
rect 404123 162147 404189 162148
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 145308 402134 150618
rect 405234 154894 405854 163000
rect 406518 162757 406578 164870
rect 407622 162757 407682 164870
rect 408358 162757 408418 164870
rect 408726 162757 408786 164870
rect 410014 164870 410124 164930
rect 410744 164930 410804 165106
rect 411288 164930 411348 165106
rect 412376 164930 412436 165106
rect 413464 164933 413524 165106
rect 413461 164932 413527 164933
rect 410744 164870 410810 164930
rect 411288 164870 411362 164930
rect 412376 164870 412466 164930
rect 406515 162756 406581 162757
rect 406515 162692 406516 162756
rect 406580 162692 406581 162756
rect 406515 162691 406581 162692
rect 407619 162756 407685 162757
rect 407619 162692 407620 162756
rect 407684 162692 407685 162756
rect 407619 162691 407685 162692
rect 408355 162756 408421 162757
rect 408355 162692 408356 162756
rect 408420 162692 408421 162756
rect 408355 162691 408421 162692
rect 408723 162756 408789 162757
rect 408723 162692 408724 162756
rect 408788 162692 408789 162756
rect 408723 162691 408789 162692
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 145308 405854 154338
rect 408954 158614 409574 163000
rect 410014 162757 410074 164870
rect 410750 162757 410810 164870
rect 411302 162757 411362 164870
rect 410011 162756 410077 162757
rect 410011 162692 410012 162756
rect 410076 162692 410077 162756
rect 410011 162691 410077 162692
rect 410747 162756 410813 162757
rect 410747 162692 410748 162756
rect 410812 162692 410813 162756
rect 410747 162691 410813 162692
rect 411299 162756 411365 162757
rect 411299 162692 411300 162756
rect 411364 162692 411365 162756
rect 411299 162691 411365 162692
rect 412406 162213 412466 164870
rect 413461 164868 413462 164932
rect 413526 164868 413527 164932
rect 413600 164930 413660 165106
rect 414552 164930 414612 165106
rect 415912 164930 415972 165106
rect 413600 164870 413754 164930
rect 414552 164870 414674 164930
rect 413461 164867 413527 164868
rect 413694 162757 413754 164870
rect 414614 162757 414674 164870
rect 415534 164870 415972 164930
rect 416048 164930 416108 165106
rect 417000 164930 417060 165106
rect 418088 164930 418148 165106
rect 418496 164930 418556 165106
rect 419448 164930 419508 165106
rect 416048 164870 416146 164930
rect 417000 164870 417066 164930
rect 418088 164870 418170 164930
rect 415534 162757 415594 164870
rect 416086 163165 416146 164870
rect 416083 163164 416149 163165
rect 416083 163100 416084 163164
rect 416148 163100 416149 163164
rect 416083 163099 416149 163100
rect 413691 162756 413757 162757
rect 413691 162692 413692 162756
rect 413756 162692 413757 162756
rect 413691 162691 413757 162692
rect 414611 162756 414677 162757
rect 414611 162692 414612 162756
rect 414676 162692 414677 162756
rect 414611 162691 414677 162692
rect 415531 162756 415597 162757
rect 415531 162692 415532 162756
rect 415596 162692 415597 162756
rect 415531 162691 415597 162692
rect 412403 162212 412469 162213
rect 412403 162148 412404 162212
rect 412468 162148 412469 162212
rect 412403 162147 412469 162148
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 145308 409574 158058
rect 415794 148394 416414 163000
rect 417006 162757 417066 164870
rect 417003 162756 417069 162757
rect 417003 162692 417004 162756
rect 417068 162692 417069 162756
rect 417003 162691 417069 162692
rect 418110 162213 418170 164870
rect 418478 164870 418556 164930
rect 419214 164870 419508 164930
rect 420672 164930 420732 165106
rect 421080 164930 421140 165106
rect 420672 164870 420746 164930
rect 418478 164253 418538 164870
rect 418475 164252 418541 164253
rect 418475 164188 418476 164252
rect 418540 164188 418541 164252
rect 418475 164187 418541 164188
rect 419214 162757 419274 164870
rect 419211 162756 419277 162757
rect 419211 162692 419212 162756
rect 419276 162692 419277 162756
rect 419211 162691 419277 162692
rect 418107 162212 418173 162213
rect 418107 162148 418108 162212
rect 418172 162148 418173 162212
rect 418107 162147 418173 162148
rect 415794 148158 415826 148394
rect 416062 148158 416146 148394
rect 416382 148158 416414 148394
rect 415794 148074 416414 148158
rect 415794 147838 415826 148074
rect 416062 147838 416146 148074
rect 416382 147838 416414 148074
rect 415794 145308 416414 147838
rect 419514 152114 420134 163000
rect 420686 162757 420746 164870
rect 421054 164870 421140 164930
rect 421760 164930 421820 165106
rect 422848 164930 422908 165106
rect 421760 164870 421850 164930
rect 422848 164870 422954 164930
rect 421054 164253 421114 164870
rect 421051 164252 421117 164253
rect 421051 164188 421052 164252
rect 421116 164188 421117 164252
rect 421051 164187 421117 164188
rect 421790 162757 421850 164870
rect 422894 162757 422954 164870
rect 423528 164661 423588 165106
rect 423936 164930 423996 165106
rect 425296 164930 425356 165106
rect 423936 164870 424058 164930
rect 423525 164660 423591 164661
rect 423525 164596 423526 164660
rect 423590 164596 423591 164660
rect 423525 164595 423591 164596
rect 420683 162756 420749 162757
rect 420683 162692 420684 162756
rect 420748 162692 420749 162756
rect 420683 162691 420749 162692
rect 421787 162756 421853 162757
rect 421787 162692 421788 162756
rect 421852 162692 421853 162756
rect 421787 162691 421853 162692
rect 422891 162756 422957 162757
rect 422891 162692 422892 162756
rect 422956 162692 422957 162756
rect 422891 162691 422957 162692
rect 419514 151878 419546 152114
rect 419782 151878 419866 152114
rect 420102 151878 420134 152114
rect 419514 151794 420134 151878
rect 419514 151558 419546 151794
rect 419782 151558 419866 151794
rect 420102 151558 420134 151794
rect 419514 145308 420134 151558
rect 423234 153954 423854 163000
rect 423998 162757 424058 164870
rect 425286 164870 425356 164930
rect 425286 162757 425346 164870
rect 425976 164797 426036 165106
rect 426384 164930 426444 165106
rect 427608 164930 427668 165106
rect 428288 164930 428348 165106
rect 426384 164870 426450 164930
rect 427608 164870 427738 164930
rect 425973 164796 426039 164797
rect 425973 164732 425974 164796
rect 426038 164732 426039 164796
rect 425973 164731 426039 164732
rect 426390 162757 426450 164870
rect 423995 162756 424061 162757
rect 423995 162692 423996 162756
rect 424060 162692 424061 162756
rect 423995 162691 424061 162692
rect 425283 162756 425349 162757
rect 425283 162692 425284 162756
rect 425348 162692 425349 162756
rect 425283 162691 425349 162692
rect 426387 162756 426453 162757
rect 426387 162692 426388 162756
rect 426452 162692 426453 162756
rect 426387 162691 426453 162692
rect 423234 153718 423266 153954
rect 423502 153718 423586 153954
rect 423822 153718 423854 153954
rect 423234 153634 423854 153718
rect 423234 153398 423266 153634
rect 423502 153398 423586 153634
rect 423822 153398 423854 153634
rect 423234 145308 423854 153398
rect 426954 157674 427574 163000
rect 427678 162213 427738 164870
rect 428230 164870 428348 164930
rect 428696 164930 428756 165106
rect 428696 164870 428842 164930
rect 428230 164253 428290 164870
rect 428227 164252 428293 164253
rect 428227 164188 428228 164252
rect 428292 164188 428293 164252
rect 428227 164187 428293 164188
rect 428782 162757 428842 164870
rect 429784 164661 429844 165106
rect 431008 164930 431068 165106
rect 430990 164870 431068 164930
rect 431144 164930 431204 165106
rect 432232 164930 432292 165106
rect 431144 164870 431234 164930
rect 429781 164660 429847 164661
rect 429781 164596 429782 164660
rect 429846 164596 429847 164660
rect 429781 164595 429847 164596
rect 430990 164253 431050 164870
rect 430987 164252 431053 164253
rect 430987 164188 430988 164252
rect 431052 164188 431053 164252
rect 430987 164187 431053 164188
rect 431174 162757 431234 164870
rect 432094 164870 432292 164930
rect 433320 164930 433380 165106
rect 433592 164930 433652 165106
rect 433320 164870 433442 164930
rect 432094 164250 432154 164870
rect 431726 164190 432154 164250
rect 431726 162757 431786 164190
rect 428779 162756 428845 162757
rect 428779 162692 428780 162756
rect 428844 162692 428845 162756
rect 428779 162691 428845 162692
rect 431171 162756 431237 162757
rect 431171 162692 431172 162756
rect 431236 162692 431237 162756
rect 431171 162691 431237 162692
rect 431723 162756 431789 162757
rect 431723 162692 431724 162756
rect 431788 162692 431789 162756
rect 431723 162691 431789 162692
rect 433382 162213 433442 164870
rect 433566 164870 433652 164930
rect 434408 164930 434468 165106
rect 435768 164930 435828 165106
rect 436040 164930 436100 165106
rect 434408 164870 434730 164930
rect 435768 164870 435834 164930
rect 427675 162212 427741 162213
rect 427675 162148 427676 162212
rect 427740 162148 427741 162212
rect 427675 162147 427741 162148
rect 433379 162212 433445 162213
rect 433379 162148 433380 162212
rect 433444 162148 433445 162212
rect 433379 162147 433445 162148
rect 433566 162077 433626 164870
rect 433563 162076 433629 162077
rect 433563 162012 433564 162076
rect 433628 162012 433629 162076
rect 433563 162011 433629 162012
rect 426954 157438 426986 157674
rect 427222 157438 427306 157674
rect 427542 157438 427574 157674
rect 426954 157354 427574 157438
rect 426954 157118 426986 157354
rect 427222 157118 427306 157354
rect 427542 157118 427574 157354
rect 426954 145308 427574 157118
rect 433794 147454 434414 163000
rect 434670 162757 434730 164870
rect 435774 162757 435834 164870
rect 435958 164870 436100 164930
rect 435958 162757 436018 164870
rect 436992 164661 437052 165106
rect 438080 164930 438140 165106
rect 438488 164930 438548 165106
rect 439168 164930 439228 165106
rect 440936 164930 440996 165106
rect 443520 164930 443580 165106
rect 445968 164930 446028 165106
rect 438080 164870 438410 164930
rect 438488 164870 438594 164930
rect 436989 164660 437055 164661
rect 436989 164596 436990 164660
rect 437054 164596 437055 164660
rect 436989 164595 437055 164596
rect 434667 162756 434733 162757
rect 434667 162692 434668 162756
rect 434732 162692 434733 162756
rect 434667 162691 434733 162692
rect 435771 162756 435837 162757
rect 435771 162692 435772 162756
rect 435836 162692 435837 162756
rect 435771 162691 435837 162692
rect 435955 162756 436021 162757
rect 435955 162692 435956 162756
rect 436020 162692 436021 162756
rect 435955 162691 436021 162692
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 145308 434414 146898
rect 437514 151174 438134 163000
rect 438350 162757 438410 164870
rect 438534 162757 438594 164870
rect 439086 164870 439228 164930
rect 440926 164870 440996 164930
rect 443502 164870 443580 164930
rect 445894 164870 446028 164930
rect 448280 164930 448340 165106
rect 448280 164870 448346 164930
rect 439086 162757 439146 164870
rect 440926 162757 440986 164870
rect 438347 162756 438413 162757
rect 438347 162692 438348 162756
rect 438412 162692 438413 162756
rect 438347 162691 438413 162692
rect 438531 162756 438597 162757
rect 438531 162692 438532 162756
rect 438596 162692 438597 162756
rect 438531 162691 438597 162692
rect 439083 162756 439149 162757
rect 439083 162692 439084 162756
rect 439148 162692 439149 162756
rect 439083 162691 439149 162692
rect 440923 162756 440989 162757
rect 440923 162692 440924 162756
rect 440988 162692 440989 162756
rect 440923 162691 440989 162692
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 145308 438134 150618
rect 441234 154894 441854 163000
rect 443502 162757 443562 164870
rect 443499 162756 443565 162757
rect 443499 162692 443500 162756
rect 443564 162692 443565 162756
rect 443499 162691 443565 162692
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 145308 441854 154338
rect 444954 158614 445574 163000
rect 445894 162757 445954 164870
rect 448286 162757 448346 164870
rect 451000 164797 451060 165106
rect 450997 164796 451063 164797
rect 450997 164732 450998 164796
rect 451062 164732 451063 164796
rect 453448 164794 453508 165106
rect 455896 164930 455956 165106
rect 458480 164930 458540 165106
rect 450997 164731 451063 164732
rect 453438 164734 453508 164794
rect 455830 164870 455956 164930
rect 458406 164870 458540 164930
rect 460928 164930 460988 165106
rect 463512 164930 463572 165106
rect 465960 164930 466020 165106
rect 468544 164930 468604 165106
rect 460928 164870 461042 164930
rect 445891 162756 445957 162757
rect 445891 162692 445892 162756
rect 445956 162692 445957 162756
rect 445891 162691 445957 162692
rect 448283 162756 448349 162757
rect 448283 162692 448284 162756
rect 448348 162692 448349 162756
rect 448283 162691 448349 162692
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 145308 445574 158058
rect 451794 148394 452414 163000
rect 453438 162757 453498 164734
rect 455830 163165 455890 164870
rect 455827 163164 455893 163165
rect 455827 163100 455828 163164
rect 455892 163100 455893 163164
rect 455827 163099 455893 163100
rect 453435 162756 453501 162757
rect 453435 162692 453436 162756
rect 453500 162692 453501 162756
rect 453435 162691 453501 162692
rect 451794 148158 451826 148394
rect 452062 148158 452146 148394
rect 452382 148158 452414 148394
rect 451794 148074 452414 148158
rect 451794 147838 451826 148074
rect 452062 147838 452146 148074
rect 452382 147838 452414 148074
rect 451794 145308 452414 147838
rect 455514 152114 456134 163000
rect 458406 162757 458466 164870
rect 458403 162756 458469 162757
rect 458403 162692 458404 162756
rect 458468 162692 458469 162756
rect 458403 162691 458469 162692
rect 455514 151878 455546 152114
rect 455782 151878 455866 152114
rect 456102 151878 456134 152114
rect 455514 151794 456134 151878
rect 455514 151558 455546 151794
rect 455782 151558 455866 151794
rect 456102 151558 456134 151794
rect 455514 145308 456134 151558
rect 459234 153954 459854 163000
rect 460982 162349 461042 164870
rect 462638 164870 463572 164930
rect 465950 164870 466020 164930
rect 468526 164870 468604 164930
rect 462638 162485 462698 164870
rect 462635 162484 462701 162485
rect 462635 162420 462636 162484
rect 462700 162420 462701 162484
rect 462635 162419 462701 162420
rect 460979 162348 461045 162349
rect 460979 162284 460980 162348
rect 461044 162284 461045 162348
rect 460979 162283 461045 162284
rect 459234 153718 459266 153954
rect 459502 153718 459586 153954
rect 459822 153718 459854 153954
rect 459234 153634 459854 153718
rect 459234 153398 459266 153634
rect 459502 153398 459586 153634
rect 459822 153398 459854 153634
rect 459234 145308 459854 153398
rect 462954 157674 463574 163000
rect 465950 161805 466010 164870
rect 468526 162621 468586 164870
rect 470992 164661 471052 165106
rect 473440 164930 473500 165106
rect 475888 164930 475948 165106
rect 478472 164930 478532 165106
rect 473440 164870 473554 164930
rect 470989 164660 471055 164661
rect 470989 164596 470990 164660
rect 471054 164596 471055 164660
rect 470989 164595 471055 164596
rect 473494 164253 473554 164870
rect 475886 164870 475948 164930
rect 478462 164870 478532 164930
rect 475886 164253 475946 164870
rect 478462 164253 478522 164870
rect 480920 164661 480980 165106
rect 483368 164930 483428 165106
rect 485952 164930 486012 165106
rect 503224 164930 503284 165106
rect 483368 164870 483490 164930
rect 485952 164870 486066 164930
rect 480917 164660 480983 164661
rect 480917 164596 480918 164660
rect 480982 164596 480983 164660
rect 480917 164595 480983 164596
rect 483430 164253 483490 164870
rect 473491 164252 473557 164253
rect 473491 164188 473492 164252
rect 473556 164188 473557 164252
rect 473491 164187 473557 164188
rect 475883 164252 475949 164253
rect 475883 164188 475884 164252
rect 475948 164188 475949 164252
rect 475883 164187 475949 164188
rect 478459 164252 478525 164253
rect 478459 164188 478460 164252
rect 478524 164188 478525 164252
rect 478459 164187 478525 164188
rect 483427 164252 483493 164253
rect 483427 164188 483428 164252
rect 483492 164188 483493 164252
rect 483427 164187 483493 164188
rect 486006 164117 486066 164870
rect 503118 164870 503284 164930
rect 503360 164930 503420 165106
rect 503360 164870 503546 164930
rect 486003 164116 486069 164117
rect 486003 164052 486004 164116
rect 486068 164052 486069 164116
rect 486003 164051 486069 164052
rect 468523 162620 468589 162621
rect 468523 162556 468524 162620
rect 468588 162556 468589 162620
rect 468523 162555 468589 162556
rect 465947 161804 466013 161805
rect 465947 161740 465948 161804
rect 466012 161740 466013 161804
rect 465947 161739 466013 161740
rect 462954 157438 462986 157674
rect 463222 157438 463306 157674
rect 463542 157438 463574 157674
rect 462954 157354 463574 157438
rect 462954 157118 462986 157354
rect 463222 157118 463306 157354
rect 463542 157118 463574 157354
rect 462954 145308 463574 157118
rect 469794 147454 470414 163000
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 145308 470414 146898
rect 473514 151174 474134 163000
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 145308 474134 150618
rect 477234 154894 477854 163000
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 145308 477854 154338
rect 480954 158614 481574 163000
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 145308 481574 158058
rect 487794 148394 488414 163000
rect 487794 148158 487826 148394
rect 488062 148158 488146 148394
rect 488382 148158 488414 148394
rect 487794 148074 488414 148158
rect 487794 147838 487826 148074
rect 488062 147838 488146 148074
rect 488382 147838 488414 148074
rect 487794 145308 488414 147838
rect 491514 152114 492134 163000
rect 491514 151878 491546 152114
rect 491782 151878 491866 152114
rect 492102 151878 492134 152114
rect 491514 151794 492134 151878
rect 491514 151558 491546 151794
rect 491782 151558 491866 151794
rect 492102 151558 492134 151794
rect 491514 145308 492134 151558
rect 495234 153954 495854 163000
rect 495234 153718 495266 153954
rect 495502 153718 495586 153954
rect 495822 153718 495854 153954
rect 495234 153634 495854 153718
rect 495234 153398 495266 153634
rect 495502 153398 495586 153634
rect 495822 153398 495854 153634
rect 495234 145308 495854 153398
rect 498954 157674 499574 163000
rect 503118 162757 503178 164870
rect 503115 162756 503181 162757
rect 503115 162692 503116 162756
rect 503180 162692 503181 162756
rect 503115 162691 503181 162692
rect 503486 162621 503546 164870
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 503483 162620 503549 162621
rect 503483 162556 503484 162620
rect 503548 162556 503549 162620
rect 503483 162555 503549 162556
rect 498954 157438 498986 157674
rect 499222 157438 499306 157674
rect 499542 157438 499574 157674
rect 498954 157354 499574 157438
rect 498954 157118 498986 157354
rect 499222 157118 499306 157354
rect 499542 157118 499574 157354
rect 498954 145308 499574 157118
rect 505794 147454 506414 163000
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 145308 506414 146898
rect 509514 151174 510134 163000
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 145308 510134 150618
rect 513234 154894 513854 163000
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 510843 145484 510909 145485
rect 510843 145420 510844 145484
rect 510908 145420 510909 145484
rect 510843 145419 510909 145420
rect 498515 144940 498581 144941
rect 498515 144876 498516 144940
rect 498580 144876 498581 144940
rect 498515 144875 498581 144876
rect 499803 144940 499869 144941
rect 499803 144876 499804 144940
rect 499868 144876 499869 144940
rect 499803 144875 499869 144876
rect 498518 143850 498578 144875
rect 499806 143850 499866 144875
rect 510846 143850 510906 145419
rect 513234 145308 513854 154338
rect 516954 158614 517574 163000
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 145308 517574 158058
rect 498464 143790 498578 143850
rect 499688 143790 499866 143850
rect 510840 143790 510906 143850
rect 498464 143202 498524 143790
rect 499688 143202 499748 143790
rect 510840 143202 510900 143790
rect 379470 142110 379714 142170
rect 379283 57220 379349 57221
rect 379283 57156 379284 57220
rect 379348 57156 379349 57220
rect 379283 57155 379349 57156
rect 379099 57084 379165 57085
rect 379099 57020 379100 57084
rect 379164 57020 379165 57084
rect 379099 57019 379165 57020
rect 379654 55230 379714 142110
rect 380272 129454 380620 129486
rect 380272 129218 380328 129454
rect 380564 129218 380620 129454
rect 380272 129134 380620 129218
rect 380272 128898 380328 129134
rect 380564 128898 380620 129134
rect 380272 128866 380620 128898
rect 516000 129454 516348 129486
rect 516000 129218 516056 129454
rect 516292 129218 516348 129454
rect 516000 129134 516348 129218
rect 516000 128898 516056 129134
rect 516292 128898 516348 129134
rect 516000 128866 516348 128898
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 380952 111454 381300 111486
rect 380952 111218 381008 111454
rect 381244 111218 381300 111454
rect 380952 111134 381300 111218
rect 380952 110898 381008 111134
rect 381244 110898 381300 111134
rect 380952 110866 381300 110898
rect 515320 111454 515668 111486
rect 515320 111218 515376 111454
rect 515612 111218 515668 111454
rect 515320 111134 515668 111218
rect 515320 110898 515376 111134
rect 515612 110898 515668 111134
rect 515320 110866 515668 110898
rect 380272 93454 380620 93486
rect 380272 93218 380328 93454
rect 380564 93218 380620 93454
rect 380272 93134 380620 93218
rect 380272 92898 380328 93134
rect 380564 92898 380620 93134
rect 380272 92866 380620 92898
rect 516000 93454 516348 93486
rect 516000 93218 516056 93454
rect 516292 93218 516348 93454
rect 516000 93134 516348 93218
rect 516000 92898 516056 93134
rect 516292 92898 516348 93134
rect 516000 92866 516348 92898
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 380952 75454 381300 75486
rect 380952 75218 381008 75454
rect 381244 75218 381300 75454
rect 380952 75134 381300 75218
rect 380952 74898 381008 75134
rect 381244 74898 381300 75134
rect 380952 74866 381300 74898
rect 515320 75454 515668 75486
rect 515320 75218 515376 75454
rect 515612 75218 515668 75454
rect 515320 75134 515668 75218
rect 515320 74898 515376 75134
rect 515612 74898 515668 75134
rect 515320 74866 515668 74898
rect 396056 59805 396116 60106
rect 397144 59805 397204 60106
rect 396053 59804 396119 59805
rect 396053 59740 396054 59804
rect 396118 59740 396119 59804
rect 396053 59739 396119 59740
rect 397141 59804 397207 59805
rect 397141 59740 397142 59804
rect 397206 59740 397207 59804
rect 397141 59739 397207 59740
rect 398232 59530 398292 60106
rect 399592 59666 399652 60106
rect 400544 59666 400604 60106
rect 399526 59606 399652 59666
rect 400446 59606 400604 59666
rect 398232 59470 398298 59530
rect 398238 58173 398298 59470
rect 398235 58172 398301 58173
rect 398235 58108 398236 58172
rect 398300 58108 398301 58172
rect 398235 58107 398301 58108
rect 377627 55180 377693 55181
rect 377627 55116 377628 55180
rect 377692 55116 377693 55180
rect 377627 55115 377693 55116
rect 379470 55170 379714 55230
rect 379794 57454 380414 58000
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379470 55045 379530 55170
rect 379467 55044 379533 55045
rect 379467 54980 379468 55044
rect 379532 54980 379533 55044
rect 379467 54979 379533 54980
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 374499 3500 374565 3501
rect 374499 3436 374500 3500
rect 374564 3436 374565 3500
rect 374499 3435 374565 3436
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 25174 384134 58000
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 28894 387854 58000
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 32614 391574 58000
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 39454 398414 58000
rect 399526 57901 399586 59606
rect 400446 57901 400506 59606
rect 401768 59530 401828 60106
rect 403128 59669 403188 60106
rect 404216 59669 404276 60106
rect 403125 59668 403191 59669
rect 403125 59604 403126 59668
rect 403190 59604 403191 59668
rect 403125 59603 403191 59604
rect 404213 59668 404279 59669
rect 404213 59604 404214 59668
rect 404278 59604 404279 59668
rect 404213 59603 404279 59604
rect 405440 59530 405500 60106
rect 406528 59530 406588 60106
rect 401734 59470 401828 59530
rect 405414 59470 405500 59530
rect 406518 59470 406588 59530
rect 407616 59530 407676 60106
rect 408296 59530 408356 60106
rect 408704 59530 408764 60106
rect 410064 59530 410124 60106
rect 407616 59470 407682 59530
rect 408296 59470 408418 59530
rect 408704 59470 408786 59530
rect 401734 58173 401794 59470
rect 405414 58173 405474 59470
rect 401731 58172 401797 58173
rect 401731 58108 401732 58172
rect 401796 58108 401797 58172
rect 401731 58107 401797 58108
rect 405411 58172 405477 58173
rect 405411 58108 405412 58172
rect 405476 58108 405477 58172
rect 405411 58107 405477 58108
rect 399523 57900 399589 57901
rect 399523 57836 399524 57900
rect 399588 57836 399589 57900
rect 399523 57835 399589 57836
rect 400443 57900 400509 57901
rect 400443 57836 400444 57900
rect 400508 57836 400509 57900
rect 400443 57835 400509 57836
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 43174 402134 58000
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 46894 405854 58000
rect 406518 57901 406578 59470
rect 407622 57901 407682 59470
rect 408358 57901 408418 59470
rect 408726 57901 408786 59470
rect 410014 59470 410124 59530
rect 410744 59530 410804 60106
rect 411288 59530 411348 60106
rect 412376 59530 412436 60106
rect 413464 59669 413524 60106
rect 413461 59668 413527 59669
rect 413461 59604 413462 59668
rect 413526 59604 413527 59668
rect 413461 59603 413527 59604
rect 413600 59530 413660 60106
rect 410744 59470 410810 59530
rect 411288 59470 411362 59530
rect 412376 59470 412466 59530
rect 406515 57900 406581 57901
rect 406515 57836 406516 57900
rect 406580 57836 406581 57900
rect 406515 57835 406581 57836
rect 407619 57900 407685 57901
rect 407619 57836 407620 57900
rect 407684 57836 407685 57900
rect 407619 57835 407685 57836
rect 408355 57900 408421 57901
rect 408355 57836 408356 57900
rect 408420 57836 408421 57900
rect 408355 57835 408421 57836
rect 408723 57900 408789 57901
rect 408723 57836 408724 57900
rect 408788 57836 408789 57900
rect 408723 57835 408789 57836
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 50614 409574 58000
rect 410014 57901 410074 59470
rect 410011 57900 410077 57901
rect 410011 57836 410012 57900
rect 410076 57836 410077 57900
rect 410011 57835 410077 57836
rect 410750 56541 410810 59470
rect 411302 56949 411362 59470
rect 412406 57901 412466 59470
rect 413510 59470 413660 59530
rect 414552 59530 414612 60106
rect 415912 59530 415972 60106
rect 414552 59470 414674 59530
rect 412403 57900 412469 57901
rect 412403 57836 412404 57900
rect 412468 57836 412469 57900
rect 412403 57835 412469 57836
rect 413510 57085 413570 59470
rect 414614 57901 414674 59470
rect 415534 59470 415972 59530
rect 416048 59530 416108 60106
rect 417000 59805 417060 60106
rect 416997 59804 417063 59805
rect 416997 59740 416998 59804
rect 417062 59740 417063 59804
rect 416997 59739 417063 59740
rect 418088 59533 418148 60106
rect 418496 59805 418556 60106
rect 418493 59804 418559 59805
rect 418493 59740 418494 59804
rect 418558 59740 418559 59804
rect 418493 59739 418559 59740
rect 419448 59669 419508 60106
rect 419445 59668 419511 59669
rect 419445 59604 419446 59668
rect 419510 59604 419511 59668
rect 419445 59603 419511 59604
rect 420672 59533 420732 60106
rect 418088 59532 418173 59533
rect 416048 59470 416146 59530
rect 418088 59470 418108 59532
rect 415534 57901 415594 59470
rect 416086 58173 416146 59470
rect 418107 59468 418108 59470
rect 418172 59468 418173 59532
rect 420672 59532 420749 59533
rect 420672 59470 420684 59532
rect 418107 59467 418173 59468
rect 420683 59468 420684 59470
rect 420748 59468 420749 59532
rect 421080 59530 421140 60106
rect 421760 59669 421820 60106
rect 421757 59668 421823 59669
rect 421757 59604 421758 59668
rect 421822 59604 421823 59668
rect 421757 59603 421823 59604
rect 420683 59467 420749 59468
rect 421054 59470 421140 59530
rect 422848 59530 422908 60106
rect 423528 59669 423588 60106
rect 423936 59805 423996 60106
rect 423933 59804 423999 59805
rect 423933 59740 423934 59804
rect 423998 59740 423999 59804
rect 423933 59739 423999 59740
rect 423525 59668 423591 59669
rect 423525 59604 423526 59668
rect 423590 59604 423591 59668
rect 423525 59603 423591 59604
rect 425296 59530 425356 60106
rect 422848 59470 422954 59530
rect 416083 58172 416149 58173
rect 416083 58108 416084 58172
rect 416148 58108 416149 58172
rect 416083 58107 416149 58108
rect 414611 57900 414677 57901
rect 414611 57836 414612 57900
rect 414676 57836 414677 57900
rect 414611 57835 414677 57836
rect 415531 57900 415597 57901
rect 415531 57836 415532 57900
rect 415596 57836 415597 57900
rect 415531 57835 415597 57836
rect 415794 57454 416414 58000
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 413507 57084 413573 57085
rect 413507 57020 413508 57084
rect 413572 57020 413573 57084
rect 413507 57019 413573 57020
rect 411299 56948 411365 56949
rect 411299 56884 411300 56948
rect 411364 56884 411365 56948
rect 411299 56883 411365 56884
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 410747 56540 410813 56541
rect 410747 56476 410748 56540
rect 410812 56476 410813 56540
rect 410747 56475 410813 56476
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 25174 420134 58000
rect 421054 57221 421114 59470
rect 422894 59397 422954 59470
rect 425286 59470 425356 59530
rect 425976 59530 426036 60106
rect 426384 59530 426444 60106
rect 427608 59530 427668 60106
rect 428288 59530 428348 60106
rect 428696 59530 428756 60106
rect 429784 59530 429844 60106
rect 431008 59530 431068 60106
rect 425976 59470 426082 59530
rect 426384 59470 426450 59530
rect 427608 59470 427738 59530
rect 425286 59397 425346 59470
rect 426022 59397 426082 59470
rect 422891 59396 422957 59397
rect 422891 59332 422892 59396
rect 422956 59332 422957 59396
rect 422891 59331 422957 59332
rect 425283 59396 425349 59397
rect 425283 59332 425284 59396
rect 425348 59332 425349 59396
rect 425283 59331 425349 59332
rect 426019 59396 426085 59397
rect 426019 59332 426020 59396
rect 426084 59332 426085 59396
rect 426019 59331 426085 59332
rect 421051 57220 421117 57221
rect 421051 57156 421052 57220
rect 421116 57156 421117 57220
rect 421051 57155 421117 57156
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 28894 423854 58000
rect 426390 57901 426450 59470
rect 426387 57900 426453 57901
rect 426387 57836 426388 57900
rect 426452 57836 426453 57900
rect 426387 57835 426453 57836
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 32614 427574 58000
rect 427678 57901 427738 59470
rect 428230 59470 428348 59530
rect 428598 59470 428756 59530
rect 429702 59470 429844 59530
rect 430990 59470 431068 59530
rect 431144 59530 431204 60106
rect 432232 59530 432292 60106
rect 433320 59530 433380 60106
rect 433592 59530 433652 60106
rect 431144 59470 431234 59530
rect 432232 59470 432338 59530
rect 433320 59470 433442 59530
rect 428230 59397 428290 59470
rect 428227 59396 428293 59397
rect 428227 59332 428228 59396
rect 428292 59332 428293 59396
rect 428227 59331 428293 59332
rect 428598 57901 428658 59470
rect 429702 57901 429762 59470
rect 427675 57900 427741 57901
rect 427675 57836 427676 57900
rect 427740 57836 427741 57900
rect 427675 57835 427741 57836
rect 428595 57900 428661 57901
rect 428595 57836 428596 57900
rect 428660 57836 428661 57900
rect 428595 57835 428661 57836
rect 429699 57900 429765 57901
rect 429699 57836 429700 57900
rect 429764 57836 429765 57900
rect 429699 57835 429765 57836
rect 430990 57221 431050 59470
rect 431174 57901 431234 59470
rect 432278 57901 432338 59470
rect 431171 57900 431237 57901
rect 431171 57836 431172 57900
rect 431236 57836 431237 57900
rect 431171 57835 431237 57836
rect 432275 57900 432341 57901
rect 432275 57836 432276 57900
rect 432340 57836 432341 57900
rect 432275 57835 432341 57836
rect 433382 57221 433442 59470
rect 433566 59470 433652 59530
rect 434408 59530 434468 60106
rect 435768 59530 435828 60106
rect 436040 59530 436100 60106
rect 436992 59530 437052 60106
rect 434408 59470 434730 59530
rect 435768 59470 435834 59530
rect 433566 57221 433626 59470
rect 430987 57220 431053 57221
rect 430987 57156 430988 57220
rect 431052 57156 431053 57220
rect 430987 57155 431053 57156
rect 433379 57220 433445 57221
rect 433379 57156 433380 57220
rect 433444 57156 433445 57220
rect 433379 57155 433445 57156
rect 433563 57220 433629 57221
rect 433563 57156 433564 57220
rect 433628 57156 433629 57220
rect 433563 57155 433629 57156
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 39454 434414 58000
rect 434670 57901 434730 59470
rect 434667 57900 434733 57901
rect 434667 57836 434668 57900
rect 434732 57836 434733 57900
rect 434667 57835 434733 57836
rect 435774 57221 435834 59470
rect 435958 59470 436100 59530
rect 436878 59470 437052 59530
rect 438080 59530 438140 60106
rect 438488 59530 438548 60106
rect 439168 59530 439228 60106
rect 440936 59530 440996 60106
rect 443520 59530 443580 60106
rect 445968 59530 446028 60106
rect 438080 59470 438410 59530
rect 438488 59470 438594 59530
rect 435958 57901 436018 59470
rect 436878 57901 436938 59470
rect 435955 57900 436021 57901
rect 435955 57836 435956 57900
rect 436020 57836 436021 57900
rect 435955 57835 436021 57836
rect 436875 57900 436941 57901
rect 436875 57836 436876 57900
rect 436940 57836 436941 57900
rect 436875 57835 436941 57836
rect 435771 57220 435837 57221
rect 435771 57156 435772 57220
rect 435836 57156 435837 57220
rect 435771 57155 435837 57156
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 43174 438134 58000
rect 438350 57901 438410 59470
rect 438534 57901 438594 59470
rect 439086 59470 439228 59530
rect 440926 59470 440996 59530
rect 443502 59470 443580 59530
rect 445894 59470 446028 59530
rect 448280 59530 448340 60106
rect 451000 59530 451060 60106
rect 453448 59530 453508 60106
rect 448280 59470 448346 59530
rect 451000 59470 451106 59530
rect 439086 57901 439146 59470
rect 440926 57901 440986 59470
rect 438347 57900 438413 57901
rect 438347 57836 438348 57900
rect 438412 57836 438413 57900
rect 438347 57835 438413 57836
rect 438531 57900 438597 57901
rect 438531 57836 438532 57900
rect 438596 57836 438597 57900
rect 438531 57835 438597 57836
rect 439083 57900 439149 57901
rect 439083 57836 439084 57900
rect 439148 57836 439149 57900
rect 439083 57835 439149 57836
rect 440923 57900 440989 57901
rect 440923 57836 440924 57900
rect 440988 57836 440989 57900
rect 440923 57835 440989 57836
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 46894 441854 58000
rect 443502 57901 443562 59470
rect 443499 57900 443565 57901
rect 443499 57836 443500 57900
rect 443564 57836 443565 57900
rect 443499 57835 443565 57836
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 50614 445574 58000
rect 445894 57901 445954 59470
rect 445891 57900 445957 57901
rect 445891 57836 445892 57900
rect 445956 57836 445957 57900
rect 445891 57835 445957 57836
rect 448286 57357 448346 59470
rect 451046 57901 451106 59470
rect 453438 59470 453508 59530
rect 455896 59530 455956 60106
rect 458480 59530 458540 60106
rect 455896 59470 456442 59530
rect 453438 58445 453498 59470
rect 453435 58444 453501 58445
rect 453435 58380 453436 58444
rect 453500 58380 453501 58444
rect 453435 58379 453501 58380
rect 451043 57900 451109 57901
rect 451043 57836 451044 57900
rect 451108 57836 451109 57900
rect 451043 57835 451109 57836
rect 451794 57454 452414 58000
rect 448283 57356 448349 57357
rect 448283 57292 448284 57356
rect 448348 57292 448349 57356
rect 448283 57291 448349 57292
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 25174 456134 58000
rect 456382 57493 456442 59470
rect 458406 59470 458540 59530
rect 460928 59530 460988 60106
rect 463512 59530 463572 60106
rect 465960 59530 466020 60106
rect 468544 59530 468604 60106
rect 470992 59530 471052 60106
rect 473440 59530 473500 60106
rect 475888 59530 475948 60106
rect 478472 59530 478532 60106
rect 480920 59530 480980 60106
rect 460928 59470 461042 59530
rect 463512 59470 463618 59530
rect 458406 58717 458466 59470
rect 458403 58716 458469 58717
rect 458403 58652 458404 58716
rect 458468 58652 458469 58716
rect 458403 58651 458469 58652
rect 456379 57492 456445 57493
rect 456379 57428 456380 57492
rect 456444 57428 456445 57492
rect 456379 57427 456445 57428
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 28894 459854 58000
rect 460982 57629 461042 59470
rect 463558 58581 463618 59470
rect 465950 59470 466020 59530
rect 468526 59470 468604 59530
rect 470918 59470 471052 59530
rect 473310 59470 473500 59530
rect 475886 59470 475948 59530
rect 478462 59470 478532 59530
rect 480854 59470 480980 59530
rect 483368 59530 483428 60106
rect 485952 59530 486012 60106
rect 503224 59669 503284 60106
rect 503221 59668 503287 59669
rect 503221 59604 503222 59668
rect 503286 59604 503287 59668
rect 503221 59603 503287 59604
rect 503360 59530 503420 60106
rect 483368 59470 483490 59530
rect 485952 59470 486066 59530
rect 465950 59397 466010 59470
rect 465947 59396 466013 59397
rect 465947 59332 465948 59396
rect 466012 59332 466013 59396
rect 465947 59331 466013 59332
rect 463555 58580 463621 58581
rect 463555 58516 463556 58580
rect 463620 58516 463621 58580
rect 463555 58515 463621 58516
rect 460979 57628 461045 57629
rect 460979 57564 460980 57628
rect 461044 57564 461045 57628
rect 460979 57563 461045 57564
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 32614 463574 58000
rect 468526 56677 468586 59470
rect 470918 58853 470978 59470
rect 470915 58852 470981 58853
rect 470915 58788 470916 58852
rect 470980 58788 470981 58852
rect 470915 58787 470981 58788
rect 468523 56676 468589 56677
rect 468523 56612 468524 56676
rect 468588 56612 468589 56676
rect 468523 56611 468589 56612
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 39454 470414 58000
rect 473310 57765 473370 59470
rect 475886 59125 475946 59470
rect 475883 59124 475949 59125
rect 475883 59060 475884 59124
rect 475948 59060 475949 59124
rect 475883 59059 475949 59060
rect 473307 57764 473373 57765
rect 473307 57700 473308 57764
rect 473372 57700 473373 57764
rect 473307 57699 473373 57700
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 43174 474134 58000
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 46894 477854 58000
rect 478462 57901 478522 59470
rect 480854 58989 480914 59470
rect 483430 59261 483490 59470
rect 486006 59261 486066 59470
rect 503302 59470 503420 59530
rect 483427 59260 483493 59261
rect 483427 59196 483428 59260
rect 483492 59196 483493 59260
rect 483427 59195 483493 59196
rect 486003 59260 486069 59261
rect 486003 59196 486004 59260
rect 486068 59196 486069 59260
rect 486003 59195 486069 59196
rect 480851 58988 480917 58989
rect 480851 58924 480852 58988
rect 480916 58924 480917 58988
rect 480851 58923 480917 58924
rect 478459 57900 478525 57901
rect 478459 57836 478460 57900
rect 478524 57836 478525 57900
rect 478459 57835 478525 57836
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 50614 481574 58000
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 57454 488414 58000
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 25174 492134 58000
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 28894 495854 58000
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 32614 499574 58000
rect 503302 57901 503362 59470
rect 503299 57900 503365 57901
rect 503299 57836 503300 57900
rect 503364 57836 503365 57900
rect 503299 57835 503365 57836
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 39454 506414 58000
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 43174 510134 58000
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 46894 513854 58000
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 50614 517574 58000
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 64250 615218 64486 615454
rect 64250 614898 64486 615134
rect 94970 615218 95206 615454
rect 94970 614898 95206 615134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 79610 597218 79846 597454
rect 79610 596898 79846 597134
rect 110330 597218 110566 597454
rect 110330 596898 110566 597134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 64250 579218 64486 579454
rect 64250 578898 64486 579134
rect 94970 579218 95206 579454
rect 94970 578898 95206 579134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 59546 547878 59782 548114
rect 59866 547878 60102 548114
rect 59546 547558 59782 547794
rect 59866 547558 60102 547794
rect 63266 549718 63502 549954
rect 63586 549718 63822 549954
rect 63266 549398 63502 549634
rect 63586 549398 63822 549634
rect 66986 553438 67222 553674
rect 67306 553438 67542 553674
rect 66986 553118 67222 553354
rect 67306 553118 67542 553354
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 91826 544158 92062 544394
rect 92146 544158 92382 544394
rect 91826 543838 92062 544074
rect 92146 543838 92382 544074
rect 95546 547878 95782 548114
rect 95866 547878 96102 548114
rect 95546 547558 95782 547794
rect 95866 547558 96102 547794
rect 99266 549718 99502 549954
rect 99586 549718 99822 549954
rect 99266 549398 99502 549634
rect 99586 549398 99822 549634
rect 102986 553438 103222 553674
rect 103306 553438 103542 553674
rect 102986 553118 103222 553354
rect 103306 553118 103542 553354
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 127826 544158 128062 544394
rect 128146 544158 128382 544394
rect 127826 543838 128062 544074
rect 128146 543838 128382 544074
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 547878 131782 548114
rect 131866 547878 132102 548114
rect 131546 547558 131782 547794
rect 131866 547558 132102 547794
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 144250 615218 144486 615454
rect 144250 614898 144486 615134
rect 174970 615218 175206 615454
rect 174970 614898 175206 615134
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 159610 597218 159846 597454
rect 159610 596898 159846 597134
rect 190330 597218 190566 597454
rect 190330 596898 190566 597134
rect 144250 579218 144486 579454
rect 144250 578898 144486 579134
rect 174970 579218 175206 579454
rect 174970 578898 175206 579134
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 135266 549718 135502 549954
rect 135586 549718 135822 549954
rect 135266 549398 135502 549634
rect 135586 549398 135822 549634
rect 138986 553438 139222 553674
rect 139306 553438 139542 553674
rect 138986 553118 139222 553354
rect 139306 553118 139542 553354
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 163826 544158 164062 544394
rect 164146 544158 164382 544394
rect 163826 543838 164062 544074
rect 164146 543838 164382 544074
rect 167546 547878 167782 548114
rect 167866 547878 168102 548114
rect 167546 547558 167782 547794
rect 167866 547558 168102 547794
rect 171266 549718 171502 549954
rect 171586 549718 171822 549954
rect 171266 549398 171502 549634
rect 171586 549398 171822 549634
rect 174986 553438 175222 553674
rect 175306 553438 175542 553674
rect 174986 553118 175222 553354
rect 175306 553118 175542 553354
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 199826 544158 200062 544394
rect 200146 544158 200382 544394
rect 199826 543838 200062 544074
rect 200146 543838 200382 544074
rect 203546 547878 203782 548114
rect 203866 547878 204102 548114
rect 203546 547558 203782 547794
rect 203866 547558 204102 547794
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 549718 207502 549954
rect 207586 549718 207822 549954
rect 207266 549398 207502 549634
rect 207586 549398 207822 549634
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 224250 615218 224486 615454
rect 224250 614898 224486 615134
rect 254970 615218 255206 615454
rect 254970 614898 255206 615134
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 239610 597218 239846 597454
rect 239610 596898 239846 597134
rect 270330 597218 270566 597454
rect 270330 596898 270566 597134
rect 224250 579218 224486 579454
rect 224250 578898 224486 579134
rect 254970 579218 255206 579454
rect 254970 578898 255206 579134
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 553438 211222 553674
rect 211306 553438 211542 553674
rect 210986 553118 211222 553354
rect 211306 553118 211542 553354
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 235826 544158 236062 544394
rect 236146 544158 236382 544394
rect 235826 543838 236062 544074
rect 236146 543838 236382 544074
rect 239546 547878 239782 548114
rect 239866 547878 240102 548114
rect 239546 547558 239782 547794
rect 239866 547558 240102 547794
rect 243266 549718 243502 549954
rect 243586 549718 243822 549954
rect 243266 549398 243502 549634
rect 243586 549398 243822 549634
rect 246986 553438 247222 553674
rect 247306 553438 247542 553674
rect 246986 553118 247222 553354
rect 247306 553118 247542 553354
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 271826 544158 272062 544394
rect 272146 544158 272382 544394
rect 271826 543838 272062 544074
rect 272146 543838 272382 544074
rect 275546 547878 275782 548114
rect 275866 547878 276102 548114
rect 275546 547558 275782 547794
rect 275866 547558 276102 547794
rect 279266 549718 279502 549954
rect 279586 549718 279822 549954
rect 279266 549398 279502 549634
rect 279586 549398 279822 549634
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 282986 553438 283222 553674
rect 283306 553438 283542 553674
rect 282986 553118 283222 553354
rect 283306 553118 283542 553354
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 79610 525218 79846 525454
rect 79610 524898 79846 525134
rect 110330 525218 110566 525454
rect 110330 524898 110566 525134
rect 141050 525218 141286 525454
rect 141050 524898 141286 525134
rect 171770 525218 172006 525454
rect 171770 524898 172006 525134
rect 202490 525218 202726 525454
rect 202490 524898 202726 525134
rect 233210 525218 233446 525454
rect 233210 524898 233446 525134
rect 263930 525218 264166 525454
rect 263930 524898 264166 525134
rect 294650 525218 294886 525454
rect 294650 524898 294886 525134
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 64250 507218 64486 507454
rect 64250 506898 64486 507134
rect 94970 507218 95206 507454
rect 94970 506898 95206 507134
rect 125690 507218 125926 507454
rect 125690 506898 125926 507134
rect 156410 507218 156646 507454
rect 156410 506898 156646 507134
rect 187130 507218 187366 507454
rect 187130 506898 187366 507134
rect 217850 507218 218086 507454
rect 217850 506898 218086 507134
rect 248570 507218 248806 507454
rect 248570 506898 248806 507134
rect 279290 507218 279526 507454
rect 279290 506898 279526 507134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 79610 489218 79846 489454
rect 79610 488898 79846 489134
rect 110330 489218 110566 489454
rect 110330 488898 110566 489134
rect 141050 489218 141286 489454
rect 141050 488898 141286 489134
rect 171770 489218 172006 489454
rect 171770 488898 172006 489134
rect 202490 489218 202726 489454
rect 202490 488898 202726 489134
rect 233210 489218 233446 489454
rect 233210 488898 233446 489134
rect 263930 489218 264166 489454
rect 263930 488898 264166 489134
rect 294650 489218 294886 489454
rect 294650 488898 294886 489134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 59546 473998 59782 474234
rect 59866 473998 60102 474234
rect 59546 473678 59782 473914
rect 59866 473678 60102 473914
rect 63266 469842 63502 470078
rect 63586 469842 63822 470078
rect 63266 469522 63502 469758
rect 63586 469522 63822 469758
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 81266 468902 81502 469138
rect 81586 468902 81822 469138
rect 81266 468582 81502 468818
rect 81586 468582 81822 468818
rect 84986 465318 85222 465554
rect 85306 465318 85542 465554
rect 84986 464998 85222 465234
rect 85306 464998 85542 465234
rect 91826 470278 92062 470514
rect 92146 470278 92382 470514
rect 91826 469958 92062 470194
rect 92146 469958 92382 470194
rect 95546 473998 95782 474234
rect 95866 473998 96102 474234
rect 95546 473678 95782 473914
rect 95866 473678 96102 473914
rect 99266 469842 99502 470078
rect 99586 469842 99822 470078
rect 99266 469522 99502 469758
rect 99586 469522 99822 469758
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 117266 468902 117502 469138
rect 117586 468902 117822 469138
rect 117266 468582 117502 468818
rect 117586 468582 117822 468818
rect 120986 465318 121222 465554
rect 121306 465318 121542 465554
rect 120986 464998 121222 465234
rect 121306 464998 121542 465234
rect 127826 470278 128062 470514
rect 128146 470278 128382 470514
rect 127826 469958 128062 470194
rect 128146 469958 128382 470194
rect 131546 473998 131782 474234
rect 131866 473998 132102 474234
rect 131546 473678 131782 473914
rect 131866 473678 132102 473914
rect 135266 469842 135502 470078
rect 135586 469842 135822 470078
rect 135266 469522 135502 469758
rect 135586 469522 135822 469758
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 153266 468902 153502 469138
rect 153586 468902 153822 469138
rect 153266 468582 153502 468818
rect 153586 468582 153822 468818
rect 156986 465318 157222 465554
rect 157306 465318 157542 465554
rect 156986 464998 157222 465234
rect 157306 464998 157542 465234
rect 163826 470278 164062 470514
rect 164146 470278 164382 470514
rect 163826 469958 164062 470194
rect 164146 469958 164382 470194
rect 167546 473998 167782 474234
rect 167866 473998 168102 474234
rect 167546 473678 167782 473914
rect 167866 473678 168102 473914
rect 171266 469842 171502 470078
rect 171586 469842 171822 470078
rect 171266 469522 171502 469758
rect 171586 469522 171822 469758
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 189266 468902 189502 469138
rect 189586 468902 189822 469138
rect 189266 468582 189502 468818
rect 189586 468582 189822 468818
rect 192986 465318 193222 465554
rect 193306 465318 193542 465554
rect 192986 464998 193222 465234
rect 193306 464998 193542 465234
rect 60328 453218 60564 453454
rect 60328 452898 60564 453134
rect 196056 453218 196292 453454
rect 196056 452898 196292 453134
rect 61008 435218 61244 435454
rect 61008 434898 61244 435134
rect 195376 435218 195612 435454
rect 195376 434898 195612 435134
rect 60328 417218 60564 417454
rect 60328 416898 60564 417134
rect 196056 417218 196292 417454
rect 196056 416898 196292 417134
rect 61008 399218 61244 399454
rect 61008 398898 61244 399134
rect 195376 399218 195612 399454
rect 195376 398898 195612 399134
rect 60328 381218 60564 381454
rect 60328 380898 60564 381134
rect 196056 381218 196292 381454
rect 196056 380898 196292 381134
rect 59546 365998 59782 366234
rect 59866 365998 60102 366234
rect 59546 365678 59782 365914
rect 59866 365678 60102 365914
rect 63266 369718 63502 369954
rect 63586 369718 63822 369954
rect 63266 369398 63502 369634
rect 63586 369398 63822 369634
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 84986 357318 85222 357554
rect 85306 357318 85542 357554
rect 84986 356998 85222 357234
rect 85306 356998 85542 357234
rect 91826 364158 92062 364394
rect 92146 364158 92382 364394
rect 91826 363838 92062 364074
rect 92146 363838 92382 364074
rect 95546 365998 95782 366234
rect 95866 365998 96102 366234
rect 95546 365678 95782 365914
rect 95866 365678 96102 365914
rect 99266 369718 99502 369954
rect 99586 369718 99822 369954
rect 99266 369398 99502 369634
rect 99586 369398 99822 369634
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 120986 357318 121222 357554
rect 121306 357318 121542 357554
rect 120986 356998 121222 357234
rect 121306 356998 121542 357234
rect 127826 364158 128062 364394
rect 128146 364158 128382 364394
rect 127826 363838 128062 364074
rect 128146 363838 128382 364074
rect 131546 365998 131782 366234
rect 131866 365998 132102 366234
rect 131546 365678 131782 365914
rect 131866 365678 132102 365914
rect 135266 369718 135502 369954
rect 135586 369718 135822 369954
rect 135266 369398 135502 369634
rect 135586 369398 135822 369634
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 156986 357318 157222 357554
rect 157306 357318 157542 357554
rect 156986 356998 157222 357234
rect 157306 356998 157542 357234
rect 163826 364158 164062 364394
rect 164146 364158 164382 364394
rect 163826 363838 164062 364074
rect 164146 363838 164382 364074
rect 167546 365998 167782 366234
rect 167866 365998 168102 366234
rect 167546 365678 167782 365914
rect 167866 365678 168102 365914
rect 171266 369718 171502 369954
rect 171586 369718 171822 369954
rect 171266 369398 171502 369634
rect 171586 369398 171822 369634
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 192986 357318 193222 357554
rect 193306 357318 193542 357554
rect 192986 356998 193222 357234
rect 193306 356998 193542 357234
rect 60328 345218 60564 345454
rect 60328 344898 60564 345134
rect 196056 345218 196292 345454
rect 196056 344898 196292 345134
rect 61008 327218 61244 327454
rect 61008 326898 61244 327134
rect 195376 327218 195612 327454
rect 195376 326898 195612 327134
rect 60328 309218 60564 309454
rect 60328 308898 60564 309134
rect 196056 309218 196292 309454
rect 196056 308898 196292 309134
rect 61008 291218 61244 291454
rect 61008 290898 61244 291134
rect 195376 291218 195612 291454
rect 195376 290898 195612 291134
rect 60328 273218 60564 273454
rect 60328 272898 60564 273134
rect 196056 273218 196292 273454
rect 196056 272898 196292 273134
rect 59546 259878 59782 260114
rect 59866 259878 60102 260114
rect 59546 259558 59782 259794
rect 59866 259558 60102 259794
rect 63266 261718 63502 261954
rect 63586 261718 63822 261954
rect 63266 261398 63502 261634
rect 63586 261398 63822 261634
rect 66986 265438 67222 265674
rect 67306 265438 67542 265674
rect 66986 265118 67222 265354
rect 67306 265118 67542 265354
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 91826 256158 92062 256394
rect 92146 256158 92382 256394
rect 91826 255838 92062 256074
rect 92146 255838 92382 256074
rect 95546 259878 95782 260114
rect 95866 259878 96102 260114
rect 95546 259558 95782 259794
rect 95866 259558 96102 259794
rect 99266 261718 99502 261954
rect 99586 261718 99822 261954
rect 99266 261398 99502 261634
rect 99586 261398 99822 261634
rect 102986 265438 103222 265674
rect 103306 265438 103542 265674
rect 102986 265118 103222 265354
rect 103306 265118 103542 265354
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 127826 256158 128062 256394
rect 128146 256158 128382 256394
rect 127826 255838 128062 256074
rect 128146 255838 128382 256074
rect 131546 259878 131782 260114
rect 131866 259878 132102 260114
rect 131546 259558 131782 259794
rect 131866 259558 132102 259794
rect 135266 261718 135502 261954
rect 135586 261718 135822 261954
rect 135266 261398 135502 261634
rect 135586 261398 135822 261634
rect 138986 265438 139222 265674
rect 139306 265438 139542 265674
rect 138986 265118 139222 265354
rect 139306 265118 139542 265354
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 163826 256158 164062 256394
rect 164146 256158 164382 256394
rect 163826 255838 164062 256074
rect 164146 255838 164382 256074
rect 167546 259878 167782 260114
rect 167866 259878 168102 260114
rect 167546 259558 167782 259794
rect 167866 259558 168102 259794
rect 171266 261718 171502 261954
rect 171586 261718 171822 261954
rect 171266 261398 171502 261634
rect 171586 261398 171822 261634
rect 174986 265438 175222 265674
rect 175306 265438 175542 265674
rect 174986 265118 175222 265354
rect 175306 265118 175542 265354
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 60328 237218 60564 237454
rect 60328 236898 60564 237134
rect 196056 237218 196292 237454
rect 196056 236898 196292 237134
rect 61008 219218 61244 219454
rect 61008 218898 61244 219134
rect 195376 219218 195612 219454
rect 195376 218898 195612 219134
rect 60328 201218 60564 201454
rect 60328 200898 60564 201134
rect 196056 201218 196292 201454
rect 196056 200898 196292 201134
rect 61008 183218 61244 183454
rect 61008 182898 61244 183134
rect 195376 183218 195612 183454
rect 195376 182898 195612 183134
rect 59546 151878 59782 152114
rect 59866 151878 60102 152114
rect 59546 151558 59782 151794
rect 59866 151558 60102 151794
rect 63266 153718 63502 153954
rect 63586 153718 63822 153954
rect 63266 153398 63502 153634
rect 63586 153398 63822 153634
rect 66986 157438 67222 157674
rect 67306 157438 67542 157674
rect 66986 157118 67222 157354
rect 67306 157118 67542 157354
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 91826 148158 92062 148394
rect 92146 148158 92382 148394
rect 91826 147838 92062 148074
rect 92146 147838 92382 148074
rect 95546 151878 95782 152114
rect 95866 151878 96102 152114
rect 95546 151558 95782 151794
rect 95866 151558 96102 151794
rect 99266 153718 99502 153954
rect 99586 153718 99822 153954
rect 99266 153398 99502 153634
rect 99586 153398 99822 153634
rect 102986 157438 103222 157674
rect 103306 157438 103542 157674
rect 102986 157118 103222 157354
rect 103306 157118 103542 157354
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 127826 148158 128062 148394
rect 128146 148158 128382 148394
rect 127826 147838 128062 148074
rect 128146 147838 128382 148074
rect 131546 151878 131782 152114
rect 131866 151878 132102 152114
rect 131546 151558 131782 151794
rect 131866 151558 132102 151794
rect 135266 153718 135502 153954
rect 135586 153718 135822 153954
rect 135266 153398 135502 153634
rect 135586 153398 135822 153634
rect 138986 157438 139222 157674
rect 139306 157438 139542 157674
rect 138986 157118 139222 157354
rect 139306 157118 139542 157354
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 163826 148158 164062 148394
rect 164146 148158 164382 148394
rect 163826 147838 164062 148074
rect 164146 147838 164382 148074
rect 167546 151878 167782 152114
rect 167866 151878 168102 152114
rect 167546 151558 167782 151794
rect 167866 151558 168102 151794
rect 171266 153718 171502 153954
rect 171586 153718 171822 153954
rect 171266 153398 171502 153634
rect 171586 153398 171822 153634
rect 174986 157438 175222 157674
rect 175306 157438 175542 157674
rect 174986 157118 175222 157354
rect 175306 157118 175542 157354
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 60328 129218 60564 129454
rect 60328 128898 60564 129134
rect 196056 129218 196292 129454
rect 196056 128898 196292 129134
rect 61008 111218 61244 111454
rect 61008 110898 61244 111134
rect 195376 111218 195612 111454
rect 195376 110898 195612 111134
rect 60328 93218 60564 93454
rect 60328 92898 60564 93134
rect 196056 93218 196292 93454
rect 196056 92898 196292 93134
rect 61008 75218 61244 75454
rect 61008 74898 61244 75134
rect 195376 75218 195612 75454
rect 195376 74898 195612 75134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 199826 470278 200062 470514
rect 200146 470278 200382 470514
rect 199826 469958 200062 470194
rect 200146 469958 200382 470194
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 364158 200062 364394
rect 200146 364158 200382 364394
rect 199826 363838 200062 364074
rect 200146 363838 200382 364074
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 256158 200062 256394
rect 200146 256158 200382 256394
rect 199826 255838 200062 256074
rect 200146 255838 200382 256074
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 148158 200062 148394
rect 200146 148158 200382 148394
rect 199826 147838 200062 148074
rect 200146 147838 200382 148074
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 203546 473998 203782 474234
rect 203866 473998 204102 474234
rect 203546 473678 203782 473914
rect 203866 473678 204102 473914
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 365998 203782 366234
rect 203866 365998 204102 366234
rect 203546 365678 203782 365914
rect 203866 365678 204102 365914
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 203546 276938 203782 277174
rect 203866 276938 204102 277174
rect 203546 276618 203782 276854
rect 203866 276618 204102 276854
rect 203546 259878 203782 260114
rect 203866 259878 204102 260114
rect 203546 259558 203782 259794
rect 203866 259558 204102 259794
rect 203546 240938 203782 241174
rect 203866 240938 204102 241174
rect 203546 240618 203782 240854
rect 203866 240618 204102 240854
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 151878 203782 152114
rect 203866 151878 204102 152114
rect 203546 151558 203782 151794
rect 203866 151558 204102 151794
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 207266 469842 207502 470078
rect 207586 469842 207822 470078
rect 207266 469522 207502 469758
rect 207586 469522 207822 469758
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 369718 207502 369954
rect 207586 369718 207822 369954
rect 207266 369398 207502 369634
rect 207586 369398 207822 369634
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 207266 280658 207502 280894
rect 207586 280658 207822 280894
rect 207266 280338 207502 280574
rect 207586 280338 207822 280574
rect 207266 261718 207502 261954
rect 207586 261718 207822 261954
rect 207266 261398 207502 261634
rect 207586 261398 207822 261634
rect 207266 244658 207502 244894
rect 207586 244658 207822 244894
rect 207266 244338 207502 244574
rect 207586 244338 207822 244574
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 153718 207502 153954
rect 207586 153718 207822 153954
rect 207266 153398 207502 153634
rect 207586 153398 207822 153634
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 210986 284378 211222 284614
rect 211306 284378 211542 284614
rect 210986 284058 211222 284294
rect 211306 284058 211542 284294
rect 210986 265438 211222 265674
rect 211306 265438 211542 265674
rect 210986 265118 211222 265354
rect 211306 265118 211542 265354
rect 210986 248378 211222 248614
rect 211306 248378 211542 248614
rect 210986 248058 211222 248294
rect 211306 248058 211542 248294
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 210986 157438 211222 157674
rect 211306 157438 211542 157674
rect 210986 157118 211222 157354
rect 211306 157118 211542 157354
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 225266 468902 225502 469138
rect 225586 468902 225822 469138
rect 225266 468582 225502 468818
rect 225586 468582 225822 468818
rect 228986 465318 229222 465554
rect 229306 465318 229542 465554
rect 228986 464998 229222 465234
rect 229306 464998 229542 465234
rect 235826 470278 236062 470514
rect 236146 470278 236382 470514
rect 235826 469958 236062 470194
rect 236146 469958 236382 470194
rect 239546 473998 239782 474234
rect 239866 473998 240102 474234
rect 239546 473678 239782 473914
rect 239866 473678 240102 473914
rect 243266 469842 243502 470078
rect 243586 469842 243822 470078
rect 243266 469522 243502 469758
rect 243586 469522 243822 469758
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 261266 468902 261502 469138
rect 261586 468902 261822 469138
rect 261266 468582 261502 468818
rect 261586 468582 261822 468818
rect 264986 465318 265222 465554
rect 265306 465318 265542 465554
rect 264986 464998 265222 465234
rect 265306 464998 265542 465234
rect 271826 470278 272062 470514
rect 272146 470278 272382 470514
rect 271826 469958 272062 470194
rect 272146 469958 272382 470194
rect 275546 473998 275782 474234
rect 275866 473998 276102 474234
rect 275546 473678 275782 473914
rect 275866 473678 276102 473914
rect 279266 469842 279502 470078
rect 279586 469842 279822 470078
rect 279266 469522 279502 469758
rect 279586 469522 279822 469758
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 297266 468902 297502 469138
rect 297586 468902 297822 469138
rect 297266 468582 297502 468818
rect 297586 468582 297822 468818
rect 300986 465318 301222 465554
rect 301306 465318 301542 465554
rect 300986 464998 301222 465234
rect 301306 464998 301542 465234
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 324250 615218 324486 615454
rect 324250 614898 324486 615134
rect 354970 615218 355206 615454
rect 354970 614898 355206 615134
rect 385690 615218 385926 615454
rect 385690 614898 385926 615134
rect 416410 615218 416646 615454
rect 416410 614898 416646 615134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 339610 597218 339846 597454
rect 339610 596898 339846 597134
rect 370330 597218 370566 597454
rect 370330 596898 370566 597134
rect 401050 597218 401286 597454
rect 401050 596898 401286 597134
rect 324250 579218 324486 579454
rect 324250 578898 324486 579134
rect 354970 579218 355206 579454
rect 354970 578898 355206 579134
rect 385690 579218 385926 579454
rect 385690 578898 385926 579134
rect 416410 579218 416646 579454
rect 416410 578898 416646 579134
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 339610 561218 339846 561454
rect 339610 560898 339846 561134
rect 370330 561218 370566 561454
rect 370330 560898 370566 561134
rect 401050 561218 401286 561454
rect 401050 560898 401286 561134
rect 324250 543218 324486 543454
rect 324250 542898 324486 543134
rect 354970 543218 355206 543454
rect 354970 542898 355206 543134
rect 385690 543218 385926 543454
rect 385690 542898 385926 543134
rect 416410 543218 416646 543454
rect 416410 542898 416646 543134
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 339610 525218 339846 525454
rect 339610 524898 339846 525134
rect 370330 525218 370566 525454
rect 370330 524898 370566 525134
rect 401050 525218 401286 525454
rect 401050 524898 401286 525134
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 220328 453218 220564 453454
rect 220328 452898 220564 453134
rect 356056 453218 356292 453454
rect 356056 452898 356292 453134
rect 221008 435218 221244 435454
rect 221008 434898 221244 435134
rect 355376 435218 355612 435454
rect 355376 434898 355612 435134
rect 220328 417218 220564 417454
rect 220328 416898 220564 417134
rect 356056 417218 356292 417454
rect 356056 416898 356292 417134
rect 221008 399218 221244 399454
rect 221008 398898 221244 399134
rect 355376 399218 355612 399454
rect 355376 398898 355612 399134
rect 220328 381218 220564 381454
rect 220328 380898 220564 381134
rect 356056 381218 356292 381454
rect 356056 380898 356292 381134
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 228986 357318 229222 357554
rect 229306 357318 229542 357554
rect 228986 356998 229222 357234
rect 229306 356998 229542 357234
rect 235826 364158 236062 364394
rect 236146 364158 236382 364394
rect 235826 363838 236062 364074
rect 236146 363838 236382 364074
rect 239546 365998 239782 366234
rect 239866 365998 240102 366234
rect 239546 365678 239782 365914
rect 239866 365678 240102 365914
rect 243266 369718 243502 369954
rect 243586 369718 243822 369954
rect 243266 369398 243502 369634
rect 243586 369398 243822 369634
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 264986 357318 265222 357554
rect 265306 357318 265542 357554
rect 264986 356998 265222 357234
rect 265306 356998 265542 357234
rect 271826 364158 272062 364394
rect 272146 364158 272382 364394
rect 271826 363838 272062 364074
rect 272146 363838 272382 364074
rect 275546 365998 275782 366234
rect 275866 365998 276102 366234
rect 275546 365678 275782 365914
rect 275866 365678 276102 365914
rect 279266 369718 279502 369954
rect 279586 369718 279822 369954
rect 279266 369398 279502 369634
rect 279586 369398 279822 369634
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 300986 357318 301222 357554
rect 301306 357318 301542 357554
rect 300986 356998 301222 357234
rect 301306 356998 301542 357234
rect 307826 364158 308062 364394
rect 308146 364158 308382 364394
rect 307826 363838 308062 364074
rect 308146 363838 308382 364074
rect 311546 365998 311782 366234
rect 311866 365998 312102 366234
rect 311546 365678 311782 365914
rect 311866 365678 312102 365914
rect 315266 369718 315502 369954
rect 315586 369718 315822 369954
rect 315266 369398 315502 369634
rect 315586 369398 315822 369634
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 336986 357318 337222 357554
rect 337306 357318 337542 357554
rect 336986 356998 337222 357234
rect 337306 356998 337542 357234
rect 343826 364158 344062 364394
rect 344146 364158 344382 364394
rect 343826 363838 344062 364074
rect 344146 363838 344382 364074
rect 347546 365998 347782 366234
rect 347866 365998 348102 366234
rect 347546 365678 347782 365914
rect 347866 365678 348102 365914
rect 351266 369718 351502 369954
rect 351586 369718 351822 369954
rect 351266 369398 351502 369634
rect 351586 369398 351822 369634
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 220328 345218 220564 345454
rect 220328 344898 220564 345134
rect 356056 345218 356292 345454
rect 356056 344898 356292 345134
rect 221008 327218 221244 327454
rect 221008 326898 221244 327134
rect 355376 327218 355612 327454
rect 355376 326898 355612 327134
rect 220328 309218 220564 309454
rect 220328 308898 220564 309134
rect 356056 309218 356292 309454
rect 356056 308898 356292 309134
rect 221008 291218 221244 291454
rect 221008 290898 221244 291134
rect 355376 291218 355612 291454
rect 355376 290898 355612 291134
rect 220328 273218 220564 273454
rect 220328 272898 220564 273134
rect 356056 273218 356292 273454
rect 356056 272898 356292 273134
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 235826 256158 236062 256394
rect 236146 256158 236382 256394
rect 235826 255838 236062 256074
rect 236146 255838 236382 256074
rect 239546 259878 239782 260114
rect 239866 259878 240102 260114
rect 239546 259558 239782 259794
rect 239866 259558 240102 259794
rect 243266 261718 243502 261954
rect 243586 261718 243822 261954
rect 243266 261398 243502 261634
rect 243586 261398 243822 261634
rect 246986 265438 247222 265674
rect 247306 265438 247542 265674
rect 246986 265118 247222 265354
rect 247306 265118 247542 265354
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 271826 256158 272062 256394
rect 272146 256158 272382 256394
rect 271826 255838 272062 256074
rect 272146 255838 272382 256074
rect 275546 259878 275782 260114
rect 275866 259878 276102 260114
rect 275546 259558 275782 259794
rect 275866 259558 276102 259794
rect 279266 261718 279502 261954
rect 279586 261718 279822 261954
rect 279266 261398 279502 261634
rect 279586 261398 279822 261634
rect 282986 265438 283222 265674
rect 283306 265438 283542 265674
rect 282986 265118 283222 265354
rect 283306 265118 283542 265354
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 307826 256158 308062 256394
rect 308146 256158 308382 256394
rect 307826 255838 308062 256074
rect 308146 255838 308382 256074
rect 311546 259878 311782 260114
rect 311866 259878 312102 260114
rect 311546 259558 311782 259794
rect 311866 259558 312102 259794
rect 315266 261718 315502 261954
rect 315586 261718 315822 261954
rect 315266 261398 315502 261634
rect 315586 261398 315822 261634
rect 318986 265438 319222 265674
rect 319306 265438 319542 265674
rect 318986 265118 319222 265354
rect 319306 265118 319542 265354
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 343826 256158 344062 256394
rect 344146 256158 344382 256394
rect 343826 255838 344062 256074
rect 344146 255838 344382 256074
rect 347546 259878 347782 260114
rect 347866 259878 348102 260114
rect 347546 259558 347782 259794
rect 347866 259558 348102 259794
rect 351266 261718 351502 261954
rect 351586 261718 351822 261954
rect 351266 261398 351502 261634
rect 351586 261398 351822 261634
rect 354986 265438 355222 265674
rect 355306 265438 355542 265674
rect 354986 265118 355222 265354
rect 355306 265118 355542 265354
rect 220328 237218 220564 237454
rect 220328 236898 220564 237134
rect 356056 237218 356292 237454
rect 356056 236898 356292 237134
rect 221008 219218 221244 219454
rect 221008 218898 221244 219134
rect 355376 219218 355612 219454
rect 355376 218898 355612 219134
rect 220328 201218 220564 201454
rect 220328 200898 220564 201134
rect 356056 201218 356292 201454
rect 356056 200898 356292 201134
rect 221008 183218 221244 183454
rect 221008 182898 221244 183134
rect 355376 183218 355612 183454
rect 355376 182898 355612 183134
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 235826 148158 236062 148394
rect 236146 148158 236382 148394
rect 235826 147838 236062 148074
rect 236146 147838 236382 148074
rect 239546 151878 239782 152114
rect 239866 151878 240102 152114
rect 239546 151558 239782 151794
rect 239866 151558 240102 151794
rect 243266 153718 243502 153954
rect 243586 153718 243822 153954
rect 243266 153398 243502 153634
rect 243586 153398 243822 153634
rect 246986 157438 247222 157674
rect 247306 157438 247542 157674
rect 246986 157118 247222 157354
rect 247306 157118 247542 157354
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 271826 148158 272062 148394
rect 272146 148158 272382 148394
rect 271826 147838 272062 148074
rect 272146 147838 272382 148074
rect 275546 151878 275782 152114
rect 275866 151878 276102 152114
rect 275546 151558 275782 151794
rect 275866 151558 276102 151794
rect 279266 153718 279502 153954
rect 279586 153718 279822 153954
rect 279266 153398 279502 153634
rect 279586 153398 279822 153634
rect 282986 157438 283222 157674
rect 283306 157438 283542 157674
rect 282986 157118 283222 157354
rect 283306 157118 283542 157354
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 307826 148158 308062 148394
rect 308146 148158 308382 148394
rect 307826 147838 308062 148074
rect 308146 147838 308382 148074
rect 311546 151878 311782 152114
rect 311866 151878 312102 152114
rect 311546 151558 311782 151794
rect 311866 151558 312102 151794
rect 315266 153718 315502 153954
rect 315586 153718 315822 153954
rect 315266 153398 315502 153634
rect 315586 153398 315822 153634
rect 318986 157438 319222 157674
rect 319306 157438 319542 157674
rect 318986 157118 319222 157354
rect 319306 157118 319542 157354
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 343826 148158 344062 148394
rect 344146 148158 344382 148394
rect 343826 147838 344062 148074
rect 344146 147838 344382 148074
rect 347546 151878 347782 152114
rect 347866 151878 348102 152114
rect 347546 151558 347782 151794
rect 347866 151558 348102 151794
rect 351266 153718 351502 153954
rect 351586 153718 351822 153954
rect 351266 153398 351502 153634
rect 351586 153398 351822 153634
rect 354986 157438 355222 157674
rect 355306 157438 355542 157674
rect 354986 157118 355222 157354
rect 355306 157118 355542 157354
rect 220328 129218 220564 129454
rect 220328 128898 220564 129134
rect 356056 129218 356292 129454
rect 356056 128898 356292 129134
rect 221008 111218 221244 111454
rect 221008 110898 221244 111134
rect 355376 111218 355612 111454
rect 355376 110898 355612 111134
rect 220328 93218 220564 93454
rect 220328 92898 220564 93134
rect 356056 93218 356292 93454
rect 356056 92898 356292 93134
rect 221008 75218 221244 75454
rect 221008 74898 221244 75134
rect 355376 75218 355612 75454
rect 355376 74898 355612 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 357318 373222 357554
rect 373306 357318 373542 357554
rect 372986 356998 373222 357234
rect 373306 356998 373542 357234
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 464250 615218 464486 615454
rect 464250 614898 464486 615134
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 464250 579218 464486 579454
rect 464250 578898 464486 579134
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 479610 597218 479846 597454
rect 479610 596898 479846 597134
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 494970 615218 495206 615454
rect 494970 614898 495206 615134
rect 494970 579218 495206 579454
rect 494970 578898 495206 579134
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 380328 453218 380564 453454
rect 380328 452898 380564 453134
rect 516056 453218 516292 453454
rect 516056 452898 516292 453134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 381008 435218 381244 435454
rect 381008 434898 381244 435134
rect 515376 435218 515612 435454
rect 515376 434898 515612 435134
rect 380328 417218 380564 417454
rect 380328 416898 380564 417134
rect 516056 417218 516292 417454
rect 516056 416898 516292 417134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 381008 399218 381244 399454
rect 381008 398898 381244 399134
rect 515376 399218 515612 399454
rect 515376 398898 515612 399134
rect 380328 381218 380564 381454
rect 380328 380898 380564 381134
rect 516056 381218 516292 381454
rect 516056 380898 516292 381134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 379826 364158 380062 364394
rect 380146 364158 380382 364394
rect 379826 363838 380062 364074
rect 380146 363838 380382 364074
rect 383546 365998 383782 366234
rect 383866 365998 384102 366234
rect 383546 365678 383782 365914
rect 383866 365678 384102 365914
rect 387266 369718 387502 369954
rect 387586 369718 387822 369954
rect 387266 369398 387502 369634
rect 387586 369398 387822 369634
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 408986 357318 409222 357554
rect 409306 357318 409542 357554
rect 408986 356998 409222 357234
rect 409306 356998 409542 357234
rect 415826 364158 416062 364394
rect 416146 364158 416382 364394
rect 415826 363838 416062 364074
rect 416146 363838 416382 364074
rect 419546 365998 419782 366234
rect 419866 365998 420102 366234
rect 419546 365678 419782 365914
rect 419866 365678 420102 365914
rect 423266 369718 423502 369954
rect 423586 369718 423822 369954
rect 423266 369398 423502 369634
rect 423586 369398 423822 369634
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 444986 357318 445222 357554
rect 445306 357318 445542 357554
rect 444986 356998 445222 357234
rect 445306 356998 445542 357234
rect 451826 364158 452062 364394
rect 452146 364158 452382 364394
rect 451826 363838 452062 364074
rect 452146 363838 452382 364074
rect 455546 365998 455782 366234
rect 455866 365998 456102 366234
rect 455546 365678 455782 365914
rect 455866 365678 456102 365914
rect 459266 369718 459502 369954
rect 459586 369718 459822 369954
rect 459266 369398 459502 369634
rect 459586 369398 459822 369634
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 480986 357318 481222 357554
rect 481306 357318 481542 357554
rect 480986 356998 481222 357234
rect 481306 356998 481542 357234
rect 487826 364158 488062 364394
rect 488146 364158 488382 364394
rect 487826 363838 488062 364074
rect 488146 363838 488382 364074
rect 491546 365998 491782 366234
rect 491866 365998 492102 366234
rect 491546 365678 491782 365914
rect 491866 365678 492102 365914
rect 495266 369718 495502 369954
rect 495586 369718 495822 369954
rect 495266 369398 495502 369634
rect 495586 369398 495822 369634
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 516986 357318 517222 357554
rect 517306 357318 517542 357554
rect 516986 356998 517222 357234
rect 517306 356998 517542 357234
rect 380328 345218 380564 345454
rect 380328 344898 380564 345134
rect 516056 345218 516292 345454
rect 516056 344898 516292 345134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 381008 327218 381244 327454
rect 381008 326898 381244 327134
rect 515376 327218 515612 327454
rect 515376 326898 515612 327134
rect 380328 309218 380564 309454
rect 380328 308898 380564 309134
rect 516056 309218 516292 309454
rect 516056 308898 516292 309134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 381008 291218 381244 291454
rect 381008 290898 381244 291134
rect 515376 291218 515612 291454
rect 515376 290898 515612 291134
rect 380328 273218 380564 273454
rect 380328 272898 380564 273134
rect 516056 273218 516292 273454
rect 516056 272898 516292 273134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 379826 256158 380062 256394
rect 380146 256158 380382 256394
rect 379826 255838 380062 256074
rect 380146 255838 380382 256074
rect 383546 259878 383782 260114
rect 383866 259878 384102 260114
rect 383546 259558 383782 259794
rect 383866 259558 384102 259794
rect 387266 261718 387502 261954
rect 387586 261718 387822 261954
rect 387266 261398 387502 261634
rect 387586 261398 387822 261634
rect 390986 265438 391222 265674
rect 391306 265438 391542 265674
rect 390986 265118 391222 265354
rect 391306 265118 391542 265354
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 415826 256158 416062 256394
rect 416146 256158 416382 256394
rect 415826 255838 416062 256074
rect 416146 255838 416382 256074
rect 419546 259878 419782 260114
rect 419866 259878 420102 260114
rect 419546 259558 419782 259794
rect 419866 259558 420102 259794
rect 423266 261718 423502 261954
rect 423586 261718 423822 261954
rect 423266 261398 423502 261634
rect 423586 261398 423822 261634
rect 426986 265438 427222 265674
rect 427306 265438 427542 265674
rect 426986 265118 427222 265354
rect 427306 265118 427542 265354
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 451826 256158 452062 256394
rect 452146 256158 452382 256394
rect 451826 255838 452062 256074
rect 452146 255838 452382 256074
rect 455546 259878 455782 260114
rect 455866 259878 456102 260114
rect 455546 259558 455782 259794
rect 455866 259558 456102 259794
rect 459266 261718 459502 261954
rect 459586 261718 459822 261954
rect 459266 261398 459502 261634
rect 459586 261398 459822 261634
rect 462986 265438 463222 265674
rect 463306 265438 463542 265674
rect 462986 265118 463222 265354
rect 463306 265118 463542 265354
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 487826 256158 488062 256394
rect 488146 256158 488382 256394
rect 487826 255838 488062 256074
rect 488146 255838 488382 256074
rect 491546 259878 491782 260114
rect 491866 259878 492102 260114
rect 491546 259558 491782 259794
rect 491866 259558 492102 259794
rect 495266 261718 495502 261954
rect 495586 261718 495822 261954
rect 495266 261398 495502 261634
rect 495586 261398 495822 261634
rect 498986 265438 499222 265674
rect 499306 265438 499542 265674
rect 498986 265118 499222 265354
rect 499306 265118 499542 265354
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 380328 237218 380564 237454
rect 380328 236898 380564 237134
rect 516056 237218 516292 237454
rect 516056 236898 516292 237134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 381008 219218 381244 219454
rect 381008 218898 381244 219134
rect 515376 219218 515612 219454
rect 515376 218898 515612 219134
rect 380328 201218 380564 201454
rect 380328 200898 380564 201134
rect 516056 201218 516292 201454
rect 516056 200898 516292 201134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 381008 183218 381244 183454
rect 381008 182898 381244 183134
rect 515376 183218 515612 183454
rect 515376 182898 515612 183134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 379826 148158 380062 148394
rect 380146 148158 380382 148394
rect 379826 147838 380062 148074
rect 380146 147838 380382 148074
rect 383546 151878 383782 152114
rect 383866 151878 384102 152114
rect 383546 151558 383782 151794
rect 383866 151558 384102 151794
rect 387266 153718 387502 153954
rect 387586 153718 387822 153954
rect 387266 153398 387502 153634
rect 387586 153398 387822 153634
rect 390986 157438 391222 157674
rect 391306 157438 391542 157674
rect 390986 157118 391222 157354
rect 391306 157118 391542 157354
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 415826 148158 416062 148394
rect 416146 148158 416382 148394
rect 415826 147838 416062 148074
rect 416146 147838 416382 148074
rect 419546 151878 419782 152114
rect 419866 151878 420102 152114
rect 419546 151558 419782 151794
rect 419866 151558 420102 151794
rect 423266 153718 423502 153954
rect 423586 153718 423822 153954
rect 423266 153398 423502 153634
rect 423586 153398 423822 153634
rect 426986 157438 427222 157674
rect 427306 157438 427542 157674
rect 426986 157118 427222 157354
rect 427306 157118 427542 157354
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 451826 148158 452062 148394
rect 452146 148158 452382 148394
rect 451826 147838 452062 148074
rect 452146 147838 452382 148074
rect 455546 151878 455782 152114
rect 455866 151878 456102 152114
rect 455546 151558 455782 151794
rect 455866 151558 456102 151794
rect 459266 153718 459502 153954
rect 459586 153718 459822 153954
rect 459266 153398 459502 153634
rect 459586 153398 459822 153634
rect 462986 157438 463222 157674
rect 463306 157438 463542 157674
rect 462986 157118 463222 157354
rect 463306 157118 463542 157354
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 487826 148158 488062 148394
rect 488146 148158 488382 148394
rect 487826 147838 488062 148074
rect 488146 147838 488382 148074
rect 491546 151878 491782 152114
rect 491866 151878 492102 152114
rect 491546 151558 491782 151794
rect 491866 151558 492102 151794
rect 495266 153718 495502 153954
rect 495586 153718 495822 153954
rect 495266 153398 495502 153634
rect 495586 153398 495822 153634
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 498986 157438 499222 157674
rect 499306 157438 499542 157674
rect 498986 157118 499222 157354
rect 499306 157118 499542 157354
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 380328 129218 380564 129454
rect 380328 128898 380564 129134
rect 516056 129218 516292 129454
rect 516056 128898 516292 129134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 381008 111218 381244 111454
rect 381008 110898 381244 111134
rect 515376 111218 515612 111454
rect 515376 110898 515612 111134
rect 380328 93218 380564 93454
rect 380328 92898 380564 93134
rect 516056 93218 516292 93454
rect 516056 92898 516292 93134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 381008 75218 381244 75454
rect 381008 74898 381244 75134
rect 515376 75218 515612 75454
rect 515376 74898 515612 75134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 64250 615454
rect 64486 615218 94970 615454
rect 95206 615218 144250 615454
rect 144486 615218 174970 615454
rect 175206 615218 224250 615454
rect 224486 615218 254970 615454
rect 255206 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 324250 615454
rect 324486 615218 354970 615454
rect 355206 615218 385690 615454
rect 385926 615218 416410 615454
rect 416646 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 464250 615454
rect 464486 615218 494970 615454
rect 495206 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 64250 615134
rect 64486 614898 94970 615134
rect 95206 614898 144250 615134
rect 144486 614898 174970 615134
rect 175206 614898 224250 615134
rect 224486 614898 254970 615134
rect 255206 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 324250 615134
rect 324486 614898 354970 615134
rect 355206 614898 385690 615134
rect 385926 614898 416410 615134
rect 416646 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 464250 615134
rect 464486 614898 494970 615134
rect 495206 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 79610 597454
rect 79846 597218 110330 597454
rect 110566 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 159610 597454
rect 159846 597218 190330 597454
rect 190566 597218 239610 597454
rect 239846 597218 270330 597454
rect 270566 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 339610 597454
rect 339846 597218 370330 597454
rect 370566 597218 401050 597454
rect 401286 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 479610 597454
rect 479846 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 79610 597134
rect 79846 596898 110330 597134
rect 110566 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 159610 597134
rect 159846 596898 190330 597134
rect 190566 596898 239610 597134
rect 239846 596898 270330 597134
rect 270566 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 339610 597134
rect 339846 596898 370330 597134
rect 370566 596898 401050 597134
rect 401286 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 479610 597134
rect 479846 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 64250 579454
rect 64486 579218 94970 579454
rect 95206 579218 144250 579454
rect 144486 579218 174970 579454
rect 175206 579218 224250 579454
rect 224486 579218 254970 579454
rect 255206 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 324250 579454
rect 324486 579218 354970 579454
rect 355206 579218 385690 579454
rect 385926 579218 416410 579454
rect 416646 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 464250 579454
rect 464486 579218 494970 579454
rect 495206 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 64250 579134
rect 64486 578898 94970 579134
rect 95206 578898 144250 579134
rect 144486 578898 174970 579134
rect 175206 578898 224250 579134
rect 224486 578898 254970 579134
rect 255206 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 324250 579134
rect 324486 578898 354970 579134
rect 355206 578898 385690 579134
rect 385926 578898 416410 579134
rect 416646 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 464250 579134
rect 464486 578898 494970 579134
rect 495206 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 339610 561454
rect 339846 561218 370330 561454
rect 370566 561218 401050 561454
rect 401286 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 339610 561134
rect 339846 560898 370330 561134
rect 370566 560898 401050 561134
rect 401286 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect 66954 553674 283574 553706
rect 66954 553438 66986 553674
rect 67222 553438 67306 553674
rect 67542 553438 102986 553674
rect 103222 553438 103306 553674
rect 103542 553438 138986 553674
rect 139222 553438 139306 553674
rect 139542 553438 174986 553674
rect 175222 553438 175306 553674
rect 175542 553438 210986 553674
rect 211222 553438 211306 553674
rect 211542 553438 246986 553674
rect 247222 553438 247306 553674
rect 247542 553438 282986 553674
rect 283222 553438 283306 553674
rect 283542 553438 283574 553674
rect 66954 553354 283574 553438
rect 66954 553118 66986 553354
rect 67222 553118 67306 553354
rect 67542 553118 102986 553354
rect 103222 553118 103306 553354
rect 103542 553118 138986 553354
rect 139222 553118 139306 553354
rect 139542 553118 174986 553354
rect 175222 553118 175306 553354
rect 175542 553118 210986 553354
rect 211222 553118 211306 553354
rect 211542 553118 246986 553354
rect 247222 553118 247306 553354
rect 247542 553118 282986 553354
rect 283222 553118 283306 553354
rect 283542 553118 283574 553354
rect 66954 553086 283574 553118
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect 63234 549954 279854 549986
rect 63234 549718 63266 549954
rect 63502 549718 63586 549954
rect 63822 549718 99266 549954
rect 99502 549718 99586 549954
rect 99822 549718 135266 549954
rect 135502 549718 135586 549954
rect 135822 549718 171266 549954
rect 171502 549718 171586 549954
rect 171822 549718 207266 549954
rect 207502 549718 207586 549954
rect 207822 549718 243266 549954
rect 243502 549718 243586 549954
rect 243822 549718 279266 549954
rect 279502 549718 279586 549954
rect 279822 549718 279854 549954
rect 63234 549634 279854 549718
rect 63234 549398 63266 549634
rect 63502 549398 63586 549634
rect 63822 549398 99266 549634
rect 99502 549398 99586 549634
rect 99822 549398 135266 549634
rect 135502 549398 135586 549634
rect 135822 549398 171266 549634
rect 171502 549398 171586 549634
rect 171822 549398 207266 549634
rect 207502 549398 207586 549634
rect 207822 549398 243266 549634
rect 243502 549398 243586 549634
rect 243822 549398 279266 549634
rect 279502 549398 279586 549634
rect 279822 549398 279854 549634
rect 63234 549366 279854 549398
rect 59514 548114 276134 548146
rect 59514 547878 59546 548114
rect 59782 547878 59866 548114
rect 60102 547878 95546 548114
rect 95782 547878 95866 548114
rect 96102 547878 131546 548114
rect 131782 547878 131866 548114
rect 132102 547878 167546 548114
rect 167782 547878 167866 548114
rect 168102 547878 203546 548114
rect 203782 547878 203866 548114
rect 204102 547878 239546 548114
rect 239782 547878 239866 548114
rect 240102 547878 275546 548114
rect 275782 547878 275866 548114
rect 276102 547878 276134 548114
rect 59514 547794 276134 547878
rect 59514 547558 59546 547794
rect 59782 547558 59866 547794
rect 60102 547558 95546 547794
rect 95782 547558 95866 547794
rect 96102 547558 131546 547794
rect 131782 547558 131866 547794
rect 132102 547558 167546 547794
rect 167782 547558 167866 547794
rect 168102 547558 203546 547794
rect 203782 547558 203866 547794
rect 204102 547558 239546 547794
rect 239782 547558 239866 547794
rect 240102 547558 275546 547794
rect 275782 547558 275866 547794
rect 276102 547558 276134 547794
rect 59514 547526 276134 547558
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect 91794 544394 272414 544426
rect 91794 544158 91826 544394
rect 92062 544158 92146 544394
rect 92382 544158 127826 544394
rect 128062 544158 128146 544394
rect 128382 544158 163826 544394
rect 164062 544158 164146 544394
rect 164382 544158 199826 544394
rect 200062 544158 200146 544394
rect 200382 544158 235826 544394
rect 236062 544158 236146 544394
rect 236382 544158 271826 544394
rect 272062 544158 272146 544394
rect 272382 544158 272414 544394
rect 91794 544074 272414 544158
rect 91794 543838 91826 544074
rect 92062 543838 92146 544074
rect 92382 543838 127826 544074
rect 128062 543838 128146 544074
rect 128382 543838 163826 544074
rect 164062 543838 164146 544074
rect 164382 543838 199826 544074
rect 200062 543838 200146 544074
rect 200382 543838 235826 544074
rect 236062 543838 236146 544074
rect 236382 543838 271826 544074
rect 272062 543838 272146 544074
rect 272382 543838 272414 544074
rect 91794 543806 272414 543838
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 324250 543454
rect 324486 543218 354970 543454
rect 355206 543218 385690 543454
rect 385926 543218 416410 543454
rect 416646 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 324250 543134
rect 324486 542898 354970 543134
rect 355206 542898 385690 543134
rect 385926 542898 416410 543134
rect 416646 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 79610 525454
rect 79846 525218 110330 525454
rect 110566 525218 141050 525454
rect 141286 525218 171770 525454
rect 172006 525218 202490 525454
rect 202726 525218 233210 525454
rect 233446 525218 263930 525454
rect 264166 525218 294650 525454
rect 294886 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 339610 525454
rect 339846 525218 370330 525454
rect 370566 525218 401050 525454
rect 401286 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 79610 525134
rect 79846 524898 110330 525134
rect 110566 524898 141050 525134
rect 141286 524898 171770 525134
rect 172006 524898 202490 525134
rect 202726 524898 233210 525134
rect 233446 524898 263930 525134
rect 264166 524898 294650 525134
rect 294886 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 339610 525134
rect 339846 524898 370330 525134
rect 370566 524898 401050 525134
rect 401286 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 64250 507454
rect 64486 507218 94970 507454
rect 95206 507218 125690 507454
rect 125926 507218 156410 507454
rect 156646 507218 187130 507454
rect 187366 507218 217850 507454
rect 218086 507218 248570 507454
rect 248806 507218 279290 507454
rect 279526 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 64250 507134
rect 64486 506898 94970 507134
rect 95206 506898 125690 507134
rect 125926 506898 156410 507134
rect 156646 506898 187130 507134
rect 187366 506898 217850 507134
rect 218086 506898 248570 507134
rect 248806 506898 279290 507134
rect 279526 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 79610 489454
rect 79846 489218 110330 489454
rect 110566 489218 141050 489454
rect 141286 489218 171770 489454
rect 172006 489218 202490 489454
rect 202726 489218 233210 489454
rect 233446 489218 263930 489454
rect 264166 489218 294650 489454
rect 294886 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 79610 489134
rect 79846 488898 110330 489134
rect 110566 488898 141050 489134
rect 141286 488898 171770 489134
rect 172006 488898 202490 489134
rect 202726 488898 233210 489134
rect 233446 488898 263930 489134
rect 264166 488898 294650 489134
rect 294886 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect 59514 474234 276134 474266
rect 59514 473998 59546 474234
rect 59782 473998 59866 474234
rect 60102 473998 95546 474234
rect 95782 473998 95866 474234
rect 96102 473998 131546 474234
rect 131782 473998 131866 474234
rect 132102 473998 167546 474234
rect 167782 473998 167866 474234
rect 168102 473998 203546 474234
rect 203782 473998 203866 474234
rect 204102 473998 239546 474234
rect 239782 473998 239866 474234
rect 240102 473998 275546 474234
rect 275782 473998 275866 474234
rect 276102 473998 276134 474234
rect 59514 473914 276134 473998
rect 59514 473678 59546 473914
rect 59782 473678 59866 473914
rect 60102 473678 95546 473914
rect 95782 473678 95866 473914
rect 96102 473678 131546 473914
rect 131782 473678 131866 473914
rect 132102 473678 167546 473914
rect 167782 473678 167866 473914
rect 168102 473678 203546 473914
rect 203782 473678 203866 473914
rect 204102 473678 239546 473914
rect 239782 473678 239866 473914
rect 240102 473678 275546 473914
rect 275782 473678 275866 473914
rect 276102 473678 276134 473914
rect 59514 473646 276134 473678
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect 91794 470514 272414 470546
rect 91794 470278 91826 470514
rect 92062 470278 92146 470514
rect 92382 470278 127826 470514
rect 128062 470278 128146 470514
rect 128382 470278 163826 470514
rect 164062 470278 164146 470514
rect 164382 470278 199826 470514
rect 200062 470278 200146 470514
rect 200382 470278 235826 470514
rect 236062 470278 236146 470514
rect 236382 470278 271826 470514
rect 272062 470278 272146 470514
rect 272382 470278 272414 470514
rect 91794 470194 272414 470278
rect 91794 470110 91826 470194
rect 63234 470078 91826 470110
rect 63234 469842 63266 470078
rect 63502 469842 63586 470078
rect 63822 469958 91826 470078
rect 92062 469958 92146 470194
rect 92382 470078 127826 470194
rect 92382 469958 99266 470078
rect 63822 469842 99266 469958
rect 99502 469842 99586 470078
rect 99822 469958 127826 470078
rect 128062 469958 128146 470194
rect 128382 470078 163826 470194
rect 128382 469958 135266 470078
rect 99822 469842 135266 469958
rect 135502 469842 135586 470078
rect 135822 469958 163826 470078
rect 164062 469958 164146 470194
rect 164382 470078 199826 470194
rect 164382 469958 171266 470078
rect 135822 469842 171266 469958
rect 171502 469842 171586 470078
rect 171822 469958 199826 470078
rect 200062 469958 200146 470194
rect 200382 470078 235826 470194
rect 200382 469958 207266 470078
rect 171822 469842 207266 469958
rect 207502 469842 207586 470078
rect 207822 469958 235826 470078
rect 236062 469958 236146 470194
rect 236382 470078 271826 470194
rect 236382 469958 243266 470078
rect 207822 469842 243266 469958
rect 243502 469842 243586 470078
rect 243822 469958 271826 470078
rect 272062 469958 272146 470194
rect 272382 470110 272414 470194
rect 272382 470078 279854 470110
rect 272382 469958 279266 470078
rect 243822 469842 279266 469958
rect 279502 469842 279586 470078
rect 279822 469842 279854 470078
rect 63234 469758 279854 469842
rect 63234 469522 63266 469758
rect 63502 469522 63586 469758
rect 63822 469522 99266 469758
rect 99502 469522 99586 469758
rect 99822 469522 135266 469758
rect 135502 469522 135586 469758
rect 135822 469522 171266 469758
rect 171502 469522 171586 469758
rect 171822 469522 207266 469758
rect 207502 469522 207586 469758
rect 207822 469522 243266 469758
rect 243502 469522 243586 469758
rect 243822 469522 279266 469758
rect 279502 469522 279586 469758
rect 279822 469522 279854 469758
rect 63234 469490 279854 469522
rect 81234 469138 297854 469170
rect 81234 468902 81266 469138
rect 81502 468902 81586 469138
rect 81822 468902 117266 469138
rect 117502 468902 117586 469138
rect 117822 468902 153266 469138
rect 153502 468902 153586 469138
rect 153822 468902 189266 469138
rect 189502 468902 189586 469138
rect 189822 468902 225266 469138
rect 225502 468902 225586 469138
rect 225822 468902 261266 469138
rect 261502 468902 261586 469138
rect 261822 468902 297266 469138
rect 297502 468902 297586 469138
rect 297822 468902 297854 469138
rect 81234 468818 297854 468902
rect 81234 468582 81266 468818
rect 81502 468582 81586 468818
rect 81822 468582 117266 468818
rect 117502 468582 117586 468818
rect 117822 468582 153266 468818
rect 153502 468582 153586 468818
rect 153822 468582 189266 468818
rect 189502 468582 189586 468818
rect 189822 468582 225266 468818
rect 225502 468582 225586 468818
rect 225822 468582 261266 468818
rect 261502 468582 261586 468818
rect 261822 468582 297266 468818
rect 297502 468582 297586 468818
rect 297822 468582 297854 468818
rect 81234 468550 297854 468582
rect 84954 465554 301574 465586
rect 84954 465318 84986 465554
rect 85222 465318 85306 465554
rect 85542 465318 120986 465554
rect 121222 465318 121306 465554
rect 121542 465318 156986 465554
rect 157222 465318 157306 465554
rect 157542 465318 192986 465554
rect 193222 465318 193306 465554
rect 193542 465318 228986 465554
rect 229222 465318 229306 465554
rect 229542 465318 264986 465554
rect 265222 465318 265306 465554
rect 265542 465318 300986 465554
rect 301222 465318 301306 465554
rect 301542 465318 301574 465554
rect 84954 465234 301574 465318
rect 84954 464998 84986 465234
rect 85222 464998 85306 465234
rect 85542 464998 120986 465234
rect 121222 464998 121306 465234
rect 121542 464998 156986 465234
rect 157222 464998 157306 465234
rect 157542 464998 192986 465234
rect 193222 464998 193306 465234
rect 193542 464998 228986 465234
rect 229222 464998 229306 465234
rect 229542 464998 264986 465234
rect 265222 464998 265306 465234
rect 265542 464998 300986 465234
rect 301222 464998 301306 465234
rect 301542 464998 301574 465234
rect 84954 464966 301574 464998
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 60328 453454
rect 60564 453218 196056 453454
rect 196292 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 220328 453454
rect 220564 453218 356056 453454
rect 356292 453218 380328 453454
rect 380564 453218 516056 453454
rect 516292 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 60328 453134
rect 60564 452898 196056 453134
rect 196292 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 220328 453134
rect 220564 452898 356056 453134
rect 356292 452898 380328 453134
rect 380564 452898 516056 453134
rect 516292 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 61008 435454
rect 61244 435218 195376 435454
rect 195612 435218 221008 435454
rect 221244 435218 355376 435454
rect 355612 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 381008 435454
rect 381244 435218 515376 435454
rect 515612 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 61008 435134
rect 61244 434898 195376 435134
rect 195612 434898 221008 435134
rect 221244 434898 355376 435134
rect 355612 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 381008 435134
rect 381244 434898 515376 435134
rect 515612 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 60328 417454
rect 60564 417218 196056 417454
rect 196292 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 220328 417454
rect 220564 417218 356056 417454
rect 356292 417218 380328 417454
rect 380564 417218 516056 417454
rect 516292 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 60328 417134
rect 60564 416898 196056 417134
rect 196292 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 220328 417134
rect 220564 416898 356056 417134
rect 356292 416898 380328 417134
rect 380564 416898 516056 417134
rect 516292 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 61008 399454
rect 61244 399218 195376 399454
rect 195612 399218 221008 399454
rect 221244 399218 355376 399454
rect 355612 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 381008 399454
rect 381244 399218 515376 399454
rect 515612 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 61008 399134
rect 61244 398898 195376 399134
rect 195612 398898 221008 399134
rect 221244 398898 355376 399134
rect 355612 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 381008 399134
rect 381244 398898 515376 399134
rect 515612 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 60328 381454
rect 60564 381218 196056 381454
rect 196292 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 220328 381454
rect 220564 381218 356056 381454
rect 356292 381218 380328 381454
rect 380564 381218 516056 381454
rect 516292 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 60328 381134
rect 60564 380898 196056 381134
rect 196292 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 220328 381134
rect 220564 380898 356056 381134
rect 356292 380898 380328 381134
rect 380564 380898 516056 381134
rect 516292 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect 63234 369954 495854 369986
rect 63234 369718 63266 369954
rect 63502 369718 63586 369954
rect 63822 369718 99266 369954
rect 99502 369718 99586 369954
rect 99822 369718 135266 369954
rect 135502 369718 135586 369954
rect 135822 369718 171266 369954
rect 171502 369718 171586 369954
rect 171822 369718 207266 369954
rect 207502 369718 207586 369954
rect 207822 369718 243266 369954
rect 243502 369718 243586 369954
rect 243822 369718 279266 369954
rect 279502 369718 279586 369954
rect 279822 369718 315266 369954
rect 315502 369718 315586 369954
rect 315822 369718 351266 369954
rect 351502 369718 351586 369954
rect 351822 369718 387266 369954
rect 387502 369718 387586 369954
rect 387822 369718 423266 369954
rect 423502 369718 423586 369954
rect 423822 369718 459266 369954
rect 459502 369718 459586 369954
rect 459822 369718 495266 369954
rect 495502 369718 495586 369954
rect 495822 369718 495854 369954
rect 63234 369634 495854 369718
rect 63234 369398 63266 369634
rect 63502 369398 63586 369634
rect 63822 369398 99266 369634
rect 99502 369398 99586 369634
rect 99822 369398 135266 369634
rect 135502 369398 135586 369634
rect 135822 369398 171266 369634
rect 171502 369398 171586 369634
rect 171822 369398 207266 369634
rect 207502 369398 207586 369634
rect 207822 369398 243266 369634
rect 243502 369398 243586 369634
rect 243822 369398 279266 369634
rect 279502 369398 279586 369634
rect 279822 369398 315266 369634
rect 315502 369398 315586 369634
rect 315822 369398 351266 369634
rect 351502 369398 351586 369634
rect 351822 369398 387266 369634
rect 387502 369398 387586 369634
rect 387822 369398 423266 369634
rect 423502 369398 423586 369634
rect 423822 369398 459266 369634
rect 459502 369398 459586 369634
rect 459822 369398 495266 369634
rect 495502 369398 495586 369634
rect 495822 369398 495854 369634
rect 63234 369366 495854 369398
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect 59514 366234 492134 366266
rect 59514 365998 59546 366234
rect 59782 365998 59866 366234
rect 60102 365998 95546 366234
rect 95782 365998 95866 366234
rect 96102 365998 131546 366234
rect 131782 365998 131866 366234
rect 132102 365998 167546 366234
rect 167782 365998 167866 366234
rect 168102 365998 203546 366234
rect 203782 365998 203866 366234
rect 204102 365998 239546 366234
rect 239782 365998 239866 366234
rect 240102 365998 275546 366234
rect 275782 365998 275866 366234
rect 276102 365998 311546 366234
rect 311782 365998 311866 366234
rect 312102 365998 347546 366234
rect 347782 365998 347866 366234
rect 348102 365998 383546 366234
rect 383782 365998 383866 366234
rect 384102 365998 419546 366234
rect 419782 365998 419866 366234
rect 420102 365998 455546 366234
rect 455782 365998 455866 366234
rect 456102 365998 491546 366234
rect 491782 365998 491866 366234
rect 492102 365998 492134 366234
rect 59514 365914 492134 365998
rect 59514 365678 59546 365914
rect 59782 365678 59866 365914
rect 60102 365678 95546 365914
rect 95782 365678 95866 365914
rect 96102 365678 131546 365914
rect 131782 365678 131866 365914
rect 132102 365678 167546 365914
rect 167782 365678 167866 365914
rect 168102 365678 203546 365914
rect 203782 365678 203866 365914
rect 204102 365678 239546 365914
rect 239782 365678 239866 365914
rect 240102 365678 275546 365914
rect 275782 365678 275866 365914
rect 276102 365678 311546 365914
rect 311782 365678 311866 365914
rect 312102 365678 347546 365914
rect 347782 365678 347866 365914
rect 348102 365678 383546 365914
rect 383782 365678 383866 365914
rect 384102 365678 419546 365914
rect 419782 365678 419866 365914
rect 420102 365678 455546 365914
rect 455782 365678 455866 365914
rect 456102 365678 491546 365914
rect 491782 365678 491866 365914
rect 492102 365678 492134 365914
rect 59514 365646 492134 365678
rect 91794 364394 488414 364426
rect 91794 364158 91826 364394
rect 92062 364158 92146 364394
rect 92382 364158 127826 364394
rect 128062 364158 128146 364394
rect 128382 364158 163826 364394
rect 164062 364158 164146 364394
rect 164382 364158 199826 364394
rect 200062 364158 200146 364394
rect 200382 364158 235826 364394
rect 236062 364158 236146 364394
rect 236382 364158 271826 364394
rect 272062 364158 272146 364394
rect 272382 364158 307826 364394
rect 308062 364158 308146 364394
rect 308382 364158 343826 364394
rect 344062 364158 344146 364394
rect 344382 364158 379826 364394
rect 380062 364158 380146 364394
rect 380382 364158 415826 364394
rect 416062 364158 416146 364394
rect 416382 364158 451826 364394
rect 452062 364158 452146 364394
rect 452382 364158 487826 364394
rect 488062 364158 488146 364394
rect 488382 364158 488414 364394
rect 91794 364074 488414 364158
rect 91794 363838 91826 364074
rect 92062 363838 92146 364074
rect 92382 363838 127826 364074
rect 128062 363838 128146 364074
rect 128382 363838 163826 364074
rect 164062 363838 164146 364074
rect 164382 363838 199826 364074
rect 200062 363838 200146 364074
rect 200382 363838 235826 364074
rect 236062 363838 236146 364074
rect 236382 363838 271826 364074
rect 272062 363838 272146 364074
rect 272382 363838 307826 364074
rect 308062 363838 308146 364074
rect 308382 363838 343826 364074
rect 344062 363838 344146 364074
rect 344382 363838 379826 364074
rect 380062 363838 380146 364074
rect 380382 363838 415826 364074
rect 416062 363838 416146 364074
rect 416382 363838 451826 364074
rect 452062 363838 452146 364074
rect 452382 363838 487826 364074
rect 488062 363838 488146 364074
rect 488382 363838 488414 364074
rect 91794 363806 488414 363838
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect 84954 357554 517574 357586
rect 84954 357318 84986 357554
rect 85222 357318 85306 357554
rect 85542 357318 120986 357554
rect 121222 357318 121306 357554
rect 121542 357318 156986 357554
rect 157222 357318 157306 357554
rect 157542 357318 192986 357554
rect 193222 357318 193306 357554
rect 193542 357318 228986 357554
rect 229222 357318 229306 357554
rect 229542 357318 264986 357554
rect 265222 357318 265306 357554
rect 265542 357318 300986 357554
rect 301222 357318 301306 357554
rect 301542 357318 336986 357554
rect 337222 357318 337306 357554
rect 337542 357318 372986 357554
rect 373222 357318 373306 357554
rect 373542 357318 408986 357554
rect 409222 357318 409306 357554
rect 409542 357318 444986 357554
rect 445222 357318 445306 357554
rect 445542 357318 480986 357554
rect 481222 357318 481306 357554
rect 481542 357318 516986 357554
rect 517222 357318 517306 357554
rect 517542 357318 517574 357554
rect 84954 357234 517574 357318
rect 84954 356998 84986 357234
rect 85222 356998 85306 357234
rect 85542 356998 120986 357234
rect 121222 356998 121306 357234
rect 121542 356998 156986 357234
rect 157222 356998 157306 357234
rect 157542 356998 192986 357234
rect 193222 356998 193306 357234
rect 193542 356998 228986 357234
rect 229222 356998 229306 357234
rect 229542 356998 264986 357234
rect 265222 356998 265306 357234
rect 265542 356998 300986 357234
rect 301222 356998 301306 357234
rect 301542 356998 336986 357234
rect 337222 356998 337306 357234
rect 337542 356998 372986 357234
rect 373222 356998 373306 357234
rect 373542 356998 408986 357234
rect 409222 356998 409306 357234
rect 409542 356998 444986 357234
rect 445222 356998 445306 357234
rect 445542 356998 480986 357234
rect 481222 356998 481306 357234
rect 481542 356998 516986 357234
rect 517222 356998 517306 357234
rect 517542 356998 517574 357234
rect 84954 356966 517574 356998
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 60328 345454
rect 60564 345218 196056 345454
rect 196292 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 220328 345454
rect 220564 345218 356056 345454
rect 356292 345218 380328 345454
rect 380564 345218 516056 345454
rect 516292 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 60328 345134
rect 60564 344898 196056 345134
rect 196292 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 220328 345134
rect 220564 344898 356056 345134
rect 356292 344898 380328 345134
rect 380564 344898 516056 345134
rect 516292 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 61008 327454
rect 61244 327218 195376 327454
rect 195612 327218 221008 327454
rect 221244 327218 355376 327454
rect 355612 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 381008 327454
rect 381244 327218 515376 327454
rect 515612 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 61008 327134
rect 61244 326898 195376 327134
rect 195612 326898 221008 327134
rect 221244 326898 355376 327134
rect 355612 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 381008 327134
rect 381244 326898 515376 327134
rect 515612 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 60328 309454
rect 60564 309218 196056 309454
rect 196292 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 220328 309454
rect 220564 309218 356056 309454
rect 356292 309218 380328 309454
rect 380564 309218 516056 309454
rect 516292 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 60328 309134
rect 60564 308898 196056 309134
rect 196292 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 220328 309134
rect 220564 308898 356056 309134
rect 356292 308898 380328 309134
rect 380564 308898 516056 309134
rect 516292 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 61008 291454
rect 61244 291218 195376 291454
rect 195612 291218 221008 291454
rect 221244 291218 355376 291454
rect 355612 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 381008 291454
rect 381244 291218 515376 291454
rect 515612 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 61008 291134
rect 61244 290898 195376 291134
rect 195612 290898 221008 291134
rect 221244 290898 355376 291134
rect 355612 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 381008 291134
rect 381244 290898 515376 291134
rect 515612 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 60328 273454
rect 60564 273218 196056 273454
rect 196292 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 220328 273454
rect 220564 273218 356056 273454
rect 356292 273218 380328 273454
rect 380564 273218 516056 273454
rect 516292 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 60328 273134
rect 60564 272898 196056 273134
rect 196292 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 220328 273134
rect 220564 272898 356056 273134
rect 356292 272898 380328 273134
rect 380564 272898 516056 273134
rect 516292 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect 66954 265674 499574 265706
rect 66954 265438 66986 265674
rect 67222 265438 67306 265674
rect 67542 265438 102986 265674
rect 103222 265438 103306 265674
rect 103542 265438 138986 265674
rect 139222 265438 139306 265674
rect 139542 265438 174986 265674
rect 175222 265438 175306 265674
rect 175542 265438 210986 265674
rect 211222 265438 211306 265674
rect 211542 265438 246986 265674
rect 247222 265438 247306 265674
rect 247542 265438 282986 265674
rect 283222 265438 283306 265674
rect 283542 265438 318986 265674
rect 319222 265438 319306 265674
rect 319542 265438 354986 265674
rect 355222 265438 355306 265674
rect 355542 265438 390986 265674
rect 391222 265438 391306 265674
rect 391542 265438 426986 265674
rect 427222 265438 427306 265674
rect 427542 265438 462986 265674
rect 463222 265438 463306 265674
rect 463542 265438 498986 265674
rect 499222 265438 499306 265674
rect 499542 265438 499574 265674
rect 66954 265354 499574 265438
rect 66954 265118 66986 265354
rect 67222 265118 67306 265354
rect 67542 265118 102986 265354
rect 103222 265118 103306 265354
rect 103542 265118 138986 265354
rect 139222 265118 139306 265354
rect 139542 265118 174986 265354
rect 175222 265118 175306 265354
rect 175542 265118 210986 265354
rect 211222 265118 211306 265354
rect 211542 265118 246986 265354
rect 247222 265118 247306 265354
rect 247542 265118 282986 265354
rect 283222 265118 283306 265354
rect 283542 265118 318986 265354
rect 319222 265118 319306 265354
rect 319542 265118 354986 265354
rect 355222 265118 355306 265354
rect 355542 265118 390986 265354
rect 391222 265118 391306 265354
rect 391542 265118 426986 265354
rect 427222 265118 427306 265354
rect 427542 265118 462986 265354
rect 463222 265118 463306 265354
rect 463542 265118 498986 265354
rect 499222 265118 499306 265354
rect 499542 265118 499574 265354
rect 66954 265086 499574 265118
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect 63234 261954 495854 261986
rect 63234 261718 63266 261954
rect 63502 261718 63586 261954
rect 63822 261718 99266 261954
rect 99502 261718 99586 261954
rect 99822 261718 135266 261954
rect 135502 261718 135586 261954
rect 135822 261718 171266 261954
rect 171502 261718 171586 261954
rect 171822 261718 207266 261954
rect 207502 261718 207586 261954
rect 207822 261718 243266 261954
rect 243502 261718 243586 261954
rect 243822 261718 279266 261954
rect 279502 261718 279586 261954
rect 279822 261718 315266 261954
rect 315502 261718 315586 261954
rect 315822 261718 351266 261954
rect 351502 261718 351586 261954
rect 351822 261718 387266 261954
rect 387502 261718 387586 261954
rect 387822 261718 423266 261954
rect 423502 261718 423586 261954
rect 423822 261718 459266 261954
rect 459502 261718 459586 261954
rect 459822 261718 495266 261954
rect 495502 261718 495586 261954
rect 495822 261718 495854 261954
rect 63234 261634 495854 261718
rect 63234 261398 63266 261634
rect 63502 261398 63586 261634
rect 63822 261398 99266 261634
rect 99502 261398 99586 261634
rect 99822 261398 135266 261634
rect 135502 261398 135586 261634
rect 135822 261398 171266 261634
rect 171502 261398 171586 261634
rect 171822 261398 207266 261634
rect 207502 261398 207586 261634
rect 207822 261398 243266 261634
rect 243502 261398 243586 261634
rect 243822 261398 279266 261634
rect 279502 261398 279586 261634
rect 279822 261398 315266 261634
rect 315502 261398 315586 261634
rect 315822 261398 351266 261634
rect 351502 261398 351586 261634
rect 351822 261398 387266 261634
rect 387502 261398 387586 261634
rect 387822 261398 423266 261634
rect 423502 261398 423586 261634
rect 423822 261398 459266 261634
rect 459502 261398 459586 261634
rect 459822 261398 495266 261634
rect 495502 261398 495586 261634
rect 495822 261398 495854 261634
rect 63234 261366 495854 261398
rect 59514 260114 492134 260146
rect 59514 259878 59546 260114
rect 59782 259878 59866 260114
rect 60102 259878 95546 260114
rect 95782 259878 95866 260114
rect 96102 259878 131546 260114
rect 131782 259878 131866 260114
rect 132102 259878 167546 260114
rect 167782 259878 167866 260114
rect 168102 259878 203546 260114
rect 203782 259878 203866 260114
rect 204102 259878 239546 260114
rect 239782 259878 239866 260114
rect 240102 259878 275546 260114
rect 275782 259878 275866 260114
rect 276102 259878 311546 260114
rect 311782 259878 311866 260114
rect 312102 259878 347546 260114
rect 347782 259878 347866 260114
rect 348102 259878 383546 260114
rect 383782 259878 383866 260114
rect 384102 259878 419546 260114
rect 419782 259878 419866 260114
rect 420102 259878 455546 260114
rect 455782 259878 455866 260114
rect 456102 259878 491546 260114
rect 491782 259878 491866 260114
rect 492102 259878 492134 260114
rect 59514 259794 492134 259878
rect 59514 259558 59546 259794
rect 59782 259558 59866 259794
rect 60102 259558 95546 259794
rect 95782 259558 95866 259794
rect 96102 259558 131546 259794
rect 131782 259558 131866 259794
rect 132102 259558 167546 259794
rect 167782 259558 167866 259794
rect 168102 259558 203546 259794
rect 203782 259558 203866 259794
rect 204102 259558 239546 259794
rect 239782 259558 239866 259794
rect 240102 259558 275546 259794
rect 275782 259558 275866 259794
rect 276102 259558 311546 259794
rect 311782 259558 311866 259794
rect 312102 259558 347546 259794
rect 347782 259558 347866 259794
rect 348102 259558 383546 259794
rect 383782 259558 383866 259794
rect 384102 259558 419546 259794
rect 419782 259558 419866 259794
rect 420102 259558 455546 259794
rect 455782 259558 455866 259794
rect 456102 259558 491546 259794
rect 491782 259558 491866 259794
rect 492102 259558 492134 259794
rect 59514 259526 492134 259558
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect 91794 256394 488414 256426
rect 91794 256158 91826 256394
rect 92062 256158 92146 256394
rect 92382 256158 127826 256394
rect 128062 256158 128146 256394
rect 128382 256158 163826 256394
rect 164062 256158 164146 256394
rect 164382 256158 199826 256394
rect 200062 256158 200146 256394
rect 200382 256158 235826 256394
rect 236062 256158 236146 256394
rect 236382 256158 271826 256394
rect 272062 256158 272146 256394
rect 272382 256158 307826 256394
rect 308062 256158 308146 256394
rect 308382 256158 343826 256394
rect 344062 256158 344146 256394
rect 344382 256158 379826 256394
rect 380062 256158 380146 256394
rect 380382 256158 415826 256394
rect 416062 256158 416146 256394
rect 416382 256158 451826 256394
rect 452062 256158 452146 256394
rect 452382 256158 487826 256394
rect 488062 256158 488146 256394
rect 488382 256158 488414 256394
rect 91794 256074 488414 256158
rect 91794 255838 91826 256074
rect 92062 255838 92146 256074
rect 92382 255838 127826 256074
rect 128062 255838 128146 256074
rect 128382 255838 163826 256074
rect 164062 255838 164146 256074
rect 164382 255838 199826 256074
rect 200062 255838 200146 256074
rect 200382 255838 235826 256074
rect 236062 255838 236146 256074
rect 236382 255838 271826 256074
rect 272062 255838 272146 256074
rect 272382 255838 307826 256074
rect 308062 255838 308146 256074
rect 308382 255838 343826 256074
rect 344062 255838 344146 256074
rect 344382 255838 379826 256074
rect 380062 255838 380146 256074
rect 380382 255838 415826 256074
rect 416062 255838 416146 256074
rect 416382 255838 451826 256074
rect 452062 255838 452146 256074
rect 452382 255838 487826 256074
rect 488062 255838 488146 256074
rect 488382 255838 488414 256074
rect 91794 255806 488414 255838
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 60328 237454
rect 60564 237218 196056 237454
rect 196292 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 220328 237454
rect 220564 237218 356056 237454
rect 356292 237218 380328 237454
rect 380564 237218 516056 237454
rect 516292 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 60328 237134
rect 60564 236898 196056 237134
rect 196292 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 220328 237134
rect 220564 236898 356056 237134
rect 356292 236898 380328 237134
rect 380564 236898 516056 237134
rect 516292 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 61008 219454
rect 61244 219218 195376 219454
rect 195612 219218 221008 219454
rect 221244 219218 355376 219454
rect 355612 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 381008 219454
rect 381244 219218 515376 219454
rect 515612 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 61008 219134
rect 61244 218898 195376 219134
rect 195612 218898 221008 219134
rect 221244 218898 355376 219134
rect 355612 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 381008 219134
rect 381244 218898 515376 219134
rect 515612 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 60328 201454
rect 60564 201218 196056 201454
rect 196292 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 220328 201454
rect 220564 201218 356056 201454
rect 356292 201218 380328 201454
rect 380564 201218 516056 201454
rect 516292 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 60328 201134
rect 60564 200898 196056 201134
rect 196292 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 220328 201134
rect 220564 200898 356056 201134
rect 356292 200898 380328 201134
rect 380564 200898 516056 201134
rect 516292 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 61008 183454
rect 61244 183218 195376 183454
rect 195612 183218 221008 183454
rect 221244 183218 355376 183454
rect 355612 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 381008 183454
rect 381244 183218 515376 183454
rect 515612 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 61008 183134
rect 61244 182898 195376 183134
rect 195612 182898 221008 183134
rect 221244 182898 355376 183134
rect 355612 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 381008 183134
rect 381244 182898 515376 183134
rect 515612 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect 66954 157674 499574 157706
rect 66954 157438 66986 157674
rect 67222 157438 67306 157674
rect 67542 157438 102986 157674
rect 103222 157438 103306 157674
rect 103542 157438 138986 157674
rect 139222 157438 139306 157674
rect 139542 157438 174986 157674
rect 175222 157438 175306 157674
rect 175542 157438 210986 157674
rect 211222 157438 211306 157674
rect 211542 157438 246986 157674
rect 247222 157438 247306 157674
rect 247542 157438 282986 157674
rect 283222 157438 283306 157674
rect 283542 157438 318986 157674
rect 319222 157438 319306 157674
rect 319542 157438 354986 157674
rect 355222 157438 355306 157674
rect 355542 157438 390986 157674
rect 391222 157438 391306 157674
rect 391542 157438 426986 157674
rect 427222 157438 427306 157674
rect 427542 157438 462986 157674
rect 463222 157438 463306 157674
rect 463542 157438 498986 157674
rect 499222 157438 499306 157674
rect 499542 157438 499574 157674
rect 66954 157354 499574 157438
rect 66954 157118 66986 157354
rect 67222 157118 67306 157354
rect 67542 157118 102986 157354
rect 103222 157118 103306 157354
rect 103542 157118 138986 157354
rect 139222 157118 139306 157354
rect 139542 157118 174986 157354
rect 175222 157118 175306 157354
rect 175542 157118 210986 157354
rect 211222 157118 211306 157354
rect 211542 157118 246986 157354
rect 247222 157118 247306 157354
rect 247542 157118 282986 157354
rect 283222 157118 283306 157354
rect 283542 157118 318986 157354
rect 319222 157118 319306 157354
rect 319542 157118 354986 157354
rect 355222 157118 355306 157354
rect 355542 157118 390986 157354
rect 391222 157118 391306 157354
rect 391542 157118 426986 157354
rect 427222 157118 427306 157354
rect 427542 157118 462986 157354
rect 463222 157118 463306 157354
rect 463542 157118 498986 157354
rect 499222 157118 499306 157354
rect 499542 157118 499574 157354
rect 66954 157086 499574 157118
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect 63234 153954 495854 153986
rect 63234 153718 63266 153954
rect 63502 153718 63586 153954
rect 63822 153718 99266 153954
rect 99502 153718 99586 153954
rect 99822 153718 135266 153954
rect 135502 153718 135586 153954
rect 135822 153718 171266 153954
rect 171502 153718 171586 153954
rect 171822 153718 207266 153954
rect 207502 153718 207586 153954
rect 207822 153718 243266 153954
rect 243502 153718 243586 153954
rect 243822 153718 279266 153954
rect 279502 153718 279586 153954
rect 279822 153718 315266 153954
rect 315502 153718 315586 153954
rect 315822 153718 351266 153954
rect 351502 153718 351586 153954
rect 351822 153718 387266 153954
rect 387502 153718 387586 153954
rect 387822 153718 423266 153954
rect 423502 153718 423586 153954
rect 423822 153718 459266 153954
rect 459502 153718 459586 153954
rect 459822 153718 495266 153954
rect 495502 153718 495586 153954
rect 495822 153718 495854 153954
rect 63234 153634 495854 153718
rect 63234 153398 63266 153634
rect 63502 153398 63586 153634
rect 63822 153398 99266 153634
rect 99502 153398 99586 153634
rect 99822 153398 135266 153634
rect 135502 153398 135586 153634
rect 135822 153398 171266 153634
rect 171502 153398 171586 153634
rect 171822 153398 207266 153634
rect 207502 153398 207586 153634
rect 207822 153398 243266 153634
rect 243502 153398 243586 153634
rect 243822 153398 279266 153634
rect 279502 153398 279586 153634
rect 279822 153398 315266 153634
rect 315502 153398 315586 153634
rect 315822 153398 351266 153634
rect 351502 153398 351586 153634
rect 351822 153398 387266 153634
rect 387502 153398 387586 153634
rect 387822 153398 423266 153634
rect 423502 153398 423586 153634
rect 423822 153398 459266 153634
rect 459502 153398 459586 153634
rect 459822 153398 495266 153634
rect 495502 153398 495586 153634
rect 495822 153398 495854 153634
rect 63234 153366 495854 153398
rect 59514 152114 492134 152146
rect 59514 151878 59546 152114
rect 59782 151878 59866 152114
rect 60102 151878 95546 152114
rect 95782 151878 95866 152114
rect 96102 151878 131546 152114
rect 131782 151878 131866 152114
rect 132102 151878 167546 152114
rect 167782 151878 167866 152114
rect 168102 151878 203546 152114
rect 203782 151878 203866 152114
rect 204102 151878 239546 152114
rect 239782 151878 239866 152114
rect 240102 151878 275546 152114
rect 275782 151878 275866 152114
rect 276102 151878 311546 152114
rect 311782 151878 311866 152114
rect 312102 151878 347546 152114
rect 347782 151878 347866 152114
rect 348102 151878 383546 152114
rect 383782 151878 383866 152114
rect 384102 151878 419546 152114
rect 419782 151878 419866 152114
rect 420102 151878 455546 152114
rect 455782 151878 455866 152114
rect 456102 151878 491546 152114
rect 491782 151878 491866 152114
rect 492102 151878 492134 152114
rect 59514 151794 492134 151878
rect 59514 151558 59546 151794
rect 59782 151558 59866 151794
rect 60102 151558 95546 151794
rect 95782 151558 95866 151794
rect 96102 151558 131546 151794
rect 131782 151558 131866 151794
rect 132102 151558 167546 151794
rect 167782 151558 167866 151794
rect 168102 151558 203546 151794
rect 203782 151558 203866 151794
rect 204102 151558 239546 151794
rect 239782 151558 239866 151794
rect 240102 151558 275546 151794
rect 275782 151558 275866 151794
rect 276102 151558 311546 151794
rect 311782 151558 311866 151794
rect 312102 151558 347546 151794
rect 347782 151558 347866 151794
rect 348102 151558 383546 151794
rect 383782 151558 383866 151794
rect 384102 151558 419546 151794
rect 419782 151558 419866 151794
rect 420102 151558 455546 151794
rect 455782 151558 455866 151794
rect 456102 151558 491546 151794
rect 491782 151558 491866 151794
rect 492102 151558 492134 151794
rect 59514 151526 492134 151558
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect 91794 148394 488414 148426
rect 91794 148158 91826 148394
rect 92062 148158 92146 148394
rect 92382 148158 127826 148394
rect 128062 148158 128146 148394
rect 128382 148158 163826 148394
rect 164062 148158 164146 148394
rect 164382 148158 199826 148394
rect 200062 148158 200146 148394
rect 200382 148158 235826 148394
rect 236062 148158 236146 148394
rect 236382 148158 271826 148394
rect 272062 148158 272146 148394
rect 272382 148158 307826 148394
rect 308062 148158 308146 148394
rect 308382 148158 343826 148394
rect 344062 148158 344146 148394
rect 344382 148158 379826 148394
rect 380062 148158 380146 148394
rect 380382 148158 415826 148394
rect 416062 148158 416146 148394
rect 416382 148158 451826 148394
rect 452062 148158 452146 148394
rect 452382 148158 487826 148394
rect 488062 148158 488146 148394
rect 488382 148158 488414 148394
rect 91794 148074 488414 148158
rect 91794 147838 91826 148074
rect 92062 147838 92146 148074
rect 92382 147838 127826 148074
rect 128062 147838 128146 148074
rect 128382 147838 163826 148074
rect 164062 147838 164146 148074
rect 164382 147838 199826 148074
rect 200062 147838 200146 148074
rect 200382 147838 235826 148074
rect 236062 147838 236146 148074
rect 236382 147838 271826 148074
rect 272062 147838 272146 148074
rect 272382 147838 307826 148074
rect 308062 147838 308146 148074
rect 308382 147838 343826 148074
rect 344062 147838 344146 148074
rect 344382 147838 379826 148074
rect 380062 147838 380146 148074
rect 380382 147838 415826 148074
rect 416062 147838 416146 148074
rect 416382 147838 451826 148074
rect 452062 147838 452146 148074
rect 452382 147838 487826 148074
rect 488062 147838 488146 148074
rect 488382 147838 488414 148074
rect 91794 147806 488414 147838
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 60328 129454
rect 60564 129218 196056 129454
rect 196292 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 220328 129454
rect 220564 129218 356056 129454
rect 356292 129218 380328 129454
rect 380564 129218 516056 129454
rect 516292 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 60328 129134
rect 60564 128898 196056 129134
rect 196292 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 220328 129134
rect 220564 128898 356056 129134
rect 356292 128898 380328 129134
rect 380564 128898 516056 129134
rect 516292 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 61008 111454
rect 61244 111218 195376 111454
rect 195612 111218 221008 111454
rect 221244 111218 355376 111454
rect 355612 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 381008 111454
rect 381244 111218 515376 111454
rect 515612 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 61008 111134
rect 61244 110898 195376 111134
rect 195612 110898 221008 111134
rect 221244 110898 355376 111134
rect 355612 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 381008 111134
rect 381244 110898 515376 111134
rect 515612 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 60328 93454
rect 60564 93218 196056 93454
rect 196292 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 220328 93454
rect 220564 93218 356056 93454
rect 356292 93218 380328 93454
rect 380564 93218 516056 93454
rect 516292 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 60328 93134
rect 60564 92898 196056 93134
rect 196292 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 220328 93134
rect 220564 92898 356056 93134
rect 356292 92898 380328 93134
rect 380564 92898 516056 93134
rect 516292 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 61008 75454
rect 61244 75218 195376 75454
rect 195612 75218 221008 75454
rect 221244 75218 355376 75454
rect 355612 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 381008 75454
rect 381244 75218 515376 75454
rect 515612 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 61008 75134
rect 61244 74898 195376 75134
rect 195612 74898 221008 75134
rect 221244 74898 355376 75134
rect 355612 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 381008 75134
rect 381244 74898 515376 75134
rect 515612 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_2kbyte_1rw1r_32x512_8  agent_1_sram2k_inst0
timestamp 0
transform 1 0 60000 0 1 60000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  agent_1_sram2k_inst1
timestamp 0
transform 1 0 60000 0 1 165000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  agent_1_sram2k_inst2
timestamp 0
transform 1 0 60000 0 1 270000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  codemaker_sram2k_inst0
timestamp 0
transform 1 0 380000 0 1 60000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  codemaker_sram2k_inst1
timestamp 0
transform 1 0 380000 0 1 165000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  codemaker_sram2k_inst2
timestamp 0
transform 1 0 380000 0 1 270000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  codemaker_sram2k_inst3
timestamp 0
transform 1 0 380000 0 1 375000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst0
timestamp 0
transform 1 0 60000 0 1 375000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst1
timestamp 0
transform 1 0 220000 0 1 60000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst2
timestamp 0
transform 1 0 220000 0 1 165000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst3
timestamp 0
transform 1 0 220000 0 1 270000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst4
timestamp 0
transform 1 0 220000 0 1 375000
box 0 0 136620 83308
use VerySimpleCPU_core  inst_agent_1
timestamp 0
transform 1 0 60000 0 1 560000
box 0 0 60955 63099
use VerySimpleCPU_core  inst_codemaker
timestamp 0
transform 1 0 220000 0 1 560000
box 0 0 60955 63099
use VerySimpleCPU_core  inst_control_tower
timestamp 0
transform 1 0 140000 0 1 560000
box 0 0 60955 63099
use main_controller  inst_main_controller
timestamp 0
transform 1 0 60000 0 1 480000
box 0 0 240000 60000
use main_memory  inst_main_memory
timestamp 0
transform 1 0 320000 0 1 520000
box 0 0 108889 111033
use uart  inst_uart
timestamp 0
transform 1 0 460000 0 1 570000
box 0 0 50000 50000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 145308 74414 163000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 145308 110414 163000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 145308 146414 163000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 145308 182414 163000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 145308 218414 163000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 145308 254414 163000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 145308 290414 163000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 145308 326414 163000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 145308 398414 163000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 145308 434414 163000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 145308 470414 163000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 145308 506414 163000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 250308 74414 268000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 250308 110414 268000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 250308 146414 268000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 250308 182414 268000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 250308 218414 268000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 250308 254414 268000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 250308 290414 268000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 250308 326414 268000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 250308 398414 268000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 250308 434414 268000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 250308 470414 268000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 250308 506414 268000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 355308 74414 373000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 355308 110414 373000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 355308 146414 373000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 355308 182414 373000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 355308 218414 373000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 355308 254414 373000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 355308 290414 373000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 355308 326414 373000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 355308 398414 373000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 355308 434414 373000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 355308 470414 373000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 355308 506414 373000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 460308 74414 478000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 460308 110414 478000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 460308 146414 478000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 460308 182414 478000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 460308 218414 478000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 460308 254414 478000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 460308 290414 478000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 460308 326414 518000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 518000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 460308 398414 518000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 542000 74414 558000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 542000 110414 558000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 542000 146414 558000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 542000 182414 558000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 542000 218414 558000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 542000 254414 558000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 460308 470414 568000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 460308 506414 568000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 625099 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 625099 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 625099 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 625099 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 625099 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 625099 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 542000 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 633033 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 633033 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 633033 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 460308 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 622000 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 622000 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 145308 78134 163000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 145308 114134 163000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 145308 150134 163000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 145308 186134 163000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 145308 222134 163000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 145308 258134 163000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 145308 294134 163000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 145308 330134 163000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 145308 402134 163000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 145308 438134 163000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 145308 474134 163000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 145308 510134 163000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 250308 78134 268000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 250308 114134 268000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 250308 150134 268000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 250308 186134 268000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 250308 222134 268000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 250308 258134 268000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 250308 294134 268000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 250308 330134 268000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 250308 402134 268000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 250308 438134 268000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 250308 474134 268000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 250308 510134 268000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 355308 78134 373000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 355308 114134 373000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 355308 150134 373000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 355308 186134 373000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 355308 222134 373000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 355308 258134 373000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 355308 294134 373000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 355308 330134 373000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 355308 402134 373000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 355308 438134 373000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 355308 474134 373000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 355308 510134 373000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 460308 78134 478000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 460308 114134 478000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 460308 150134 478000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 460308 186134 478000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 460308 222134 478000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 460308 258134 478000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 460308 294134 478000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 460308 330134 518000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 518000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 460308 402134 518000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 542000 78134 558000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 542000 114134 558000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 542000 150134 558000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 542000 186134 558000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 542000 222134 558000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 542000 258134 558000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 460308 474134 568000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 460308 510134 568000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 625099 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 625099 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 625099 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 625099 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 625099 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 625099 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 542000 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 633033 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 633033 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 633033 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 460308 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 622000 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 622000 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s 81234 468550 297854 469170 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 145308 81854 163000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 145308 117854 163000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 145308 153854 163000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 145308 189854 163000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 145308 225854 163000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 145308 261854 163000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 145308 297854 163000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 145308 333854 163000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 145308 405854 163000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 145308 441854 163000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 145308 477854 163000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 145308 513854 163000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 250308 81854 268000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 250308 117854 268000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 250308 153854 268000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 250308 189854 268000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 250308 225854 268000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 250308 261854 268000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 250308 297854 268000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 250308 333854 268000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 250308 405854 268000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 250308 441854 268000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 250308 477854 268000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 250308 513854 268000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 355308 81854 373000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 355308 117854 373000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 355308 153854 373000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 355308 189854 373000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 355308 225854 373000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 355308 261854 373000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 355308 297854 373000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 355308 333854 373000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 355308 405854 373000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 355308 441854 373000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 355308 477854 373000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 355308 513854 373000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 460308 81854 478000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 460308 117854 478000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 460308 153854 478000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 460308 189854 478000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 460308 225854 478000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 460308 261854 478000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 460308 297854 478000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 460308 333854 518000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 518000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 460308 405854 518000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 542000 81854 558000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 542000 117854 558000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 542000 153854 558000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 542000 189854 558000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 542000 225854 558000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 542000 261854 558000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 460308 477854 568000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 625099 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 625099 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 625099 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 625099 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 625099 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 625099 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 542000 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 633033 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 633033 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 633033 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 460308 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 622000 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 460308 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s 84954 356966 517574 357586 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s 84954 464966 301574 465586 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 145308 85574 163000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 145308 121574 163000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 145308 157574 163000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 145308 193574 163000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 145308 229574 163000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 145308 265574 163000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 145308 301574 163000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 145308 337574 163000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 145308 409574 163000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 145308 445574 163000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 145308 481574 163000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 145308 517574 163000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 250308 85574 268000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 250308 121574 268000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 250308 157574 268000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 250308 193574 268000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 250308 229574 268000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 250308 265574 268000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 250308 301574 268000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 250308 337574 268000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 250308 409574 268000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 250308 445574 268000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 250308 481574 268000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 250308 517574 268000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 355308 85574 373000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 355308 121574 373000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 355308 157574 373000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 355308 193574 373000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 355308 229574 373000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 355308 265574 373000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 355308 301574 373000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 355308 337574 373000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 355308 409574 373000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 355308 445574 373000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 355308 481574 373000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 355308 517574 373000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 460308 85574 478000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 460308 121574 478000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 460308 157574 478000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 460308 193574 478000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 460308 229574 478000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 460308 265574 478000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 460308 301574 478000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 460308 337574 518000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 518000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 460308 409574 518000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 542000 85574 558000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 542000 121574 558000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 542000 157574 558000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 542000 193574 558000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 542000 229574 558000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 542000 265574 558000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 460308 481574 568000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 625099 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 625099 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 625099 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 625099 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 625099 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 625099 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 542000 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 633033 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 633033 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 633033 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 460308 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 622000 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 460308 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 63234 153366 495854 153986 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 63234 261366 495854 261986 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 63234 369366 495854 369986 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 63234 469490 279854 470110 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 63234 549366 279854 549986 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 145308 63854 163000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 145308 99854 163000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 145308 135854 163000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 145308 171854 163000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 145308 243854 163000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 145308 279854 163000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 145308 315854 163000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 145308 351854 163000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 145308 387854 163000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 145308 423854 163000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 145308 459854 163000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 145308 495854 163000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 250308 63854 268000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 250308 99854 268000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 250308 135854 268000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 250308 171854 268000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 250308 243854 268000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 250308 279854 268000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 250308 315854 268000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 250308 351854 268000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 250308 387854 268000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 250308 423854 268000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 250308 459854 268000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 250308 495854 268000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 355308 63854 373000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 355308 99854 373000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 355308 135854 373000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 355308 171854 373000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 355308 243854 373000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 355308 279854 373000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 355308 315854 373000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 355308 351854 373000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 355308 387854 373000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 355308 423854 373000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 355308 459854 373000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 355308 495854 373000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 460308 63854 478000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 460308 99854 478000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 460308 135854 478000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 460308 171854 478000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 478000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 460308 243854 478000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 460308 279854 478000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 460308 351854 518000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 460308 387854 518000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 460308 423854 518000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 542000 63854 558000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 542000 99854 558000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 542000 171854 558000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 542000 243854 558000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 542000 279854 558000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 460308 459854 568000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 460308 495854 568000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 625099 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 625099 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 542000 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 625099 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 542000 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 625099 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 625099 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 460308 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 633033 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 633033 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 633033 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 622000 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 622000 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 66954 157086 499574 157706 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 66954 265086 499574 265706 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 66954 553086 283574 553706 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 145308 67574 163000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 145308 103574 163000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 145308 139574 163000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 145308 175574 163000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 145308 247574 163000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 145308 283574 163000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 145308 319574 163000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 145308 355574 163000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 145308 391574 163000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 145308 427574 163000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 145308 463574 163000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 145308 499574 163000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 250308 67574 268000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 250308 103574 268000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 250308 139574 268000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 250308 175574 268000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 250308 247574 268000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 250308 283574 268000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 250308 319574 268000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 250308 355574 268000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 250308 391574 268000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 250308 427574 268000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 250308 463574 268000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 250308 499574 268000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 355308 67574 373000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 355308 103574 373000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 355308 139574 373000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 355308 175574 373000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 355308 247574 373000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 355308 283574 373000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 355308 319574 373000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 355308 355574 373000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 355308 391574 373000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 355308 427574 373000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 355308 463574 373000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 355308 499574 373000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 460308 67574 478000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 460308 103574 478000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 460308 139574 478000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 460308 175574 478000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 478000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 460308 247574 478000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 460308 283574 478000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 460308 319574 518000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 460308 355574 518000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 460308 391574 518000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 460308 427574 518000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 542000 67574 558000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 542000 103574 558000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 542000 139574 558000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 542000 175574 558000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 542000 247574 558000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 542000 283574 558000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 460308 463574 568000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 460308 499574 568000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 625099 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 625099 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 625099 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 625099 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 542000 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 625099 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 625099 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 633033 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 633033 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 633033 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 633033 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 622000 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 622000 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 91794 147806 488414 148426 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 91794 255806 488414 256426 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 91794 363806 488414 364426 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 91794 469926 272414 470546 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 91794 543806 272414 544426 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 145308 92414 163000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 145308 128414 163000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 145308 164414 163000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 145308 236414 163000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 145308 272414 163000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 145308 308414 163000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 145308 344414 163000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 145308 380414 163000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 145308 416414 163000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 145308 452414 163000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 145308 488414 163000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 250308 92414 268000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 250308 128414 268000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 250308 164414 268000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 250308 236414 268000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 250308 272414 268000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 250308 308414 268000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 250308 344414 268000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 250308 380414 268000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 250308 416414 268000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 250308 452414 268000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 250308 488414 268000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 355308 92414 373000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 355308 128414 373000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 355308 164414 373000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 355308 236414 373000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 355308 272414 373000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 355308 308414 373000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 355308 344414 373000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 355308 380414 373000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 355308 416414 373000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 355308 452414 373000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 355308 488414 373000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 460308 92414 478000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 460308 128414 478000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 460308 164414 478000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 478000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 460308 236414 478000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 460308 272414 478000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 460308 344414 518000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 460308 380414 518000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 460308 416414 518000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 542000 92414 558000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 542000 164414 558000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 542000 200414 558000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 542000 236414 558000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 542000 272414 558000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 460308 488414 568000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 625099 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 542000 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 625099 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 625099 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 625099 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 625099 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 460308 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 633033 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 633033 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 633033 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 460308 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 622000 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 59514 151526 492134 152146 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 59514 259526 492134 260146 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 59514 365646 492134 366266 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 59514 473646 276134 474266 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 59514 547526 276134 548146 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 145308 60134 163000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 145308 96134 163000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 145308 132134 163000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 145308 168134 163000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 145308 240134 163000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 145308 276134 163000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 145308 312134 163000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 145308 348134 163000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 145308 384134 163000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 145308 420134 163000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 145308 456134 163000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 145308 492134 163000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 250308 60134 268000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 250308 96134 268000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 250308 132134 268000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 250308 168134 268000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 250308 240134 268000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 250308 276134 268000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 250308 312134 268000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 250308 348134 268000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 250308 384134 268000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 250308 420134 268000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 250308 456134 268000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 250308 492134 268000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 355308 60134 373000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 355308 96134 373000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 355308 132134 373000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 355308 168134 373000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 355308 240134 373000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 355308 276134 373000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 355308 312134 373000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 355308 348134 373000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 355308 384134 373000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 355308 420134 373000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 355308 456134 373000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 355308 492134 373000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 460308 60134 478000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 460308 96134 478000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 460308 132134 478000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 460308 168134 478000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 478000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 460308 240134 478000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 460308 276134 478000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 460308 348134 518000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 460308 384134 518000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 460308 420134 518000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 542000 60134 558000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 542000 96134 558000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 542000 168134 558000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 542000 240134 558000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 542000 276134 558000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 460308 492134 568000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 625099 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 625099 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 542000 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 625099 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 542000 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 625099 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 625099 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 460308 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 633033 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 633033 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 633033 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 460308 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 622000 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
