magic
tech sky130A
magscale 1 2
timestamp 1655467073
<< metal1 >>
rect 235166 700340 235172 700392
rect 235224 700380 235230 700392
rect 307018 700380 307024 700392
rect 235224 700352 307024 700380
rect 235224 700340 235230 700352
rect 307018 700340 307024 700352
rect 307076 700340 307082 700392
rect 429838 700340 429844 700392
rect 429896 700380 429902 700392
rect 434714 700380 434720 700392
rect 429896 700352 434720 700380
rect 429896 700340 429902 700352
rect 434714 700340 434720 700352
rect 434772 700340 434778 700392
rect 170306 700272 170312 700324
rect 170364 700312 170370 700324
rect 434806 700312 434812 700324
rect 170364 700284 434812 700312
rect 170364 700272 170370 700284
rect 434806 700272 434812 700284
rect 434864 700272 434870 700324
rect 364334 692044 364340 692096
rect 364392 692084 364398 692096
rect 427814 692084 427820 692096
rect 364392 692056 427820 692084
rect 364392 692044 364398 692056
rect 427814 692044 427820 692056
rect 427872 692044 427878 692096
rect 147306 683136 147312 683188
rect 147364 683176 147370 683188
rect 580166 683176 580172 683188
rect 147364 683148 580172 683176
rect 147364 683136 147370 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 59170 654780 59176 654832
rect 59228 654820 59234 654832
rect 542354 654820 542360 654832
rect 59228 654792 542360 654820
rect 59228 654780 59234 654792
rect 542354 654780 542360 654792
rect 542412 654780 542418 654832
rect 104894 653352 104900 653404
rect 104952 653392 104958 653404
rect 434898 653392 434904 653404
rect 104952 653364 434904 653392
rect 104952 653352 104958 653364
rect 434898 653352 434904 653364
rect 434956 653352 434962 653404
rect 299474 651992 299480 652044
rect 299532 652032 299538 652044
rect 405826 652032 405832 652044
rect 299532 652004 405832 652032
rect 299532 651992 299538 652004
rect 405826 651992 405832 652004
rect 405884 651992 405890 652044
rect 324222 649272 324228 649324
rect 324280 649312 324286 649324
rect 494054 649312 494060 649324
rect 324280 649284 494060 649312
rect 324280 649272 324286 649284
rect 494054 649272 494060 649284
rect 494112 649272 494118 649324
rect 311158 648116 311164 648168
rect 311216 648156 311222 648168
rect 337562 648156 337568 648168
rect 311216 648128 337568 648156
rect 311216 648116 311222 648128
rect 337562 648116 337568 648128
rect 337620 648116 337626 648168
rect 316770 648048 316776 648100
rect 316828 648088 316834 648100
rect 342254 648088 342260 648100
rect 316828 648060 342260 648088
rect 316828 648048 316834 648060
rect 342254 648048 342260 648060
rect 342312 648048 342318 648100
rect 323762 647980 323768 648032
rect 323820 648020 323826 648032
rect 401686 648020 401692 648032
rect 323820 647992 401692 648020
rect 323820 647980 323826 647992
rect 401686 647980 401692 647992
rect 401744 647980 401750 648032
rect 322382 647912 322388 647964
rect 322440 647952 322446 647964
rect 346578 647952 346584 647964
rect 322440 647924 346584 647952
rect 322440 647912 322446 647924
rect 346578 647912 346584 647924
rect 346636 647912 346642 647964
rect 322290 647844 322296 647896
rect 322348 647884 322354 647896
rect 355594 647884 355600 647896
rect 322348 647856 355600 647884
rect 322348 647844 322354 647856
rect 355594 647844 355600 647856
rect 355652 647844 355658 647896
rect 323578 647776 323584 647828
rect 323636 647816 323642 647828
rect 369118 647816 369124 647828
rect 323636 647788 369124 647816
rect 323636 647776 323642 647788
rect 369118 647776 369124 647788
rect 369176 647776 369182 647828
rect 318150 647708 318156 647760
rect 318208 647748 318214 647760
rect 364610 647748 364616 647760
rect 318208 647720 364616 647748
rect 318208 647708 318214 647720
rect 364610 647708 364616 647720
rect 364668 647708 364674 647760
rect 320910 647640 320916 647692
rect 320968 647680 320974 647692
rect 373994 647680 374000 647692
rect 320968 647652 374000 647680
rect 320968 647640 320974 647652
rect 373994 647640 374000 647652
rect 374052 647640 374058 647692
rect 324866 647572 324872 647624
rect 324924 647612 324930 647624
rect 378134 647612 378140 647624
rect 324924 647584 378140 647612
rect 324924 647572 324930 647584
rect 378134 647572 378140 647584
rect 378192 647572 378198 647624
rect 324774 647504 324780 647556
rect 324832 647544 324838 647556
rect 387794 647544 387800 647556
rect 324832 647516 387800 647544
rect 324832 647504 324838 647516
rect 387794 647504 387800 647516
rect 387852 647504 387858 647556
rect 313918 647436 313924 647488
rect 313976 647476 313982 647488
rect 383654 647476 383660 647488
rect 313976 647448 383660 647476
rect 313976 647436 313982 647448
rect 383654 647436 383660 647448
rect 383712 647436 383718 647488
rect 320818 647368 320824 647420
rect 320876 647408 320882 647420
rect 392302 647408 392308 647420
rect 320876 647380 392308 647408
rect 320876 647368 320882 647380
rect 392302 647368 392308 647380
rect 392360 647368 392366 647420
rect 322198 647300 322204 647352
rect 322256 647340 322262 647352
rect 432874 647340 432880 647352
rect 322256 647312 432880 647340
rect 322256 647300 322262 647312
rect 432874 647300 432880 647312
rect 432932 647300 432938 647352
rect 323670 647232 323676 647284
rect 323728 647272 323734 647284
rect 328546 647272 328552 647284
rect 323728 647244 328552 647272
rect 323728 647232 323734 647244
rect 328546 647232 328552 647244
rect 328604 647232 328610 647284
rect 391934 647232 391940 647284
rect 391992 647272 391998 647284
rect 396810 647272 396816 647284
rect 391992 647244 396816 647272
rect 391992 647232 391998 647244
rect 396810 647232 396816 647244
rect 396868 647232 396874 647284
rect 419534 647232 419540 647284
rect 419592 647272 419598 647284
rect 457438 647272 457444 647284
rect 419592 647244 457444 647272
rect 419592 647232 419598 647244
rect 457438 647232 457444 647244
rect 457496 647232 457502 647284
rect 235074 646484 235080 646536
rect 235132 646524 235138 646536
rect 391934 646524 391940 646536
rect 235132 646496 391940 646524
rect 235132 646484 235138 646496
rect 391934 646484 391940 646496
rect 391992 646484 391998 646536
rect 322566 646416 322572 646468
rect 322624 646456 322630 646468
rect 436186 646456 436192 646468
rect 322624 646428 436192 646456
rect 322624 646416 322630 646428
rect 436186 646416 436192 646428
rect 436244 646416 436250 646468
rect 322474 646348 322480 646400
rect 322532 646388 322538 646400
rect 436094 646388 436100 646400
rect 322532 646360 436100 646388
rect 322532 646348 322538 646360
rect 436094 646348 436100 646360
rect 436152 646348 436158 646400
rect 319438 646280 319444 646332
rect 319496 646320 319502 646332
rect 436278 646320 436284 646332
rect 319496 646292 436284 646320
rect 319496 646280 319502 646292
rect 436278 646280 436284 646292
rect 436336 646280 436342 646332
rect 234338 646212 234344 646264
rect 234396 646252 234402 646264
rect 360194 646252 360200 646264
rect 234396 646224 360200 646252
rect 234396 646212 234402 646224
rect 360194 646212 360200 646224
rect 360252 646212 360258 646264
rect 316862 646144 316868 646196
rect 316920 646184 316926 646196
rect 457530 646184 457536 646196
rect 316920 646156 457536 646184
rect 316920 646144 316926 646156
rect 457530 646144 457536 646156
rect 457588 646144 457594 646196
rect 319530 646076 319536 646128
rect 319588 646116 319594 646128
rect 494790 646116 494796 646128
rect 319588 646088 494796 646116
rect 319588 646076 319594 646088
rect 494790 646076 494796 646088
rect 494848 646076 494854 646128
rect 239398 646008 239404 646060
rect 239456 646048 239462 646060
rect 433334 646048 433340 646060
rect 239456 646020 433340 646048
rect 239456 646008 239462 646020
rect 433334 646008 433340 646020
rect 433392 646008 433398 646060
rect 18598 645940 18604 645992
rect 18656 645980 18662 645992
rect 414842 645980 414848 645992
rect 18656 645952 414848 645980
rect 18656 645940 18662 645952
rect 414842 645940 414848 645952
rect 414900 645940 414906 645992
rect 238018 645872 238024 645924
rect 238076 645912 238082 645924
rect 419534 645912 419540 645924
rect 238076 645884 419540 645912
rect 238076 645872 238082 645884
rect 419534 645872 419540 645884
rect 419592 645872 419598 645924
rect 147490 645328 147496 645380
rect 147548 645368 147554 645380
rect 164510 645368 164516 645380
rect 147548 645340 164516 645368
rect 147548 645328 147554 645340
rect 164510 645328 164516 645340
rect 164568 645328 164574 645380
rect 145466 645260 145472 645312
rect 145524 645300 145530 645312
rect 145524 645272 156828 645300
rect 145524 645260 145530 645272
rect 144914 645124 144920 645176
rect 144972 645164 144978 645176
rect 156598 645164 156604 645176
rect 144972 645136 156604 645164
rect 144972 645124 144978 645136
rect 156598 645124 156604 645136
rect 156656 645124 156662 645176
rect 156800 645164 156828 645272
rect 196066 645164 196072 645176
rect 156800 645136 196072 645164
rect 196066 645124 196072 645136
rect 196124 645124 196130 645176
rect 238846 645124 238852 645176
rect 238904 645164 238910 645176
rect 580350 645164 580356 645176
rect 238904 645136 580356 645164
rect 238904 645124 238910 645136
rect 580350 645124 580356 645136
rect 580408 645124 580414 645176
rect 142798 645056 142804 645108
rect 142856 645096 142862 645108
rect 161474 645096 161480 645108
rect 142856 645068 161480 645096
rect 142856 645056 142862 645068
rect 161474 645056 161480 645068
rect 161532 645056 161538 645108
rect 215018 645056 215024 645108
rect 215076 645096 215082 645108
rect 245654 645096 245660 645108
rect 215076 645068 245660 645096
rect 215076 645056 215082 645068
rect 245654 645056 245660 645068
rect 245712 645056 245718 645108
rect 322658 645056 322664 645108
rect 322716 645096 322722 645108
rect 457714 645096 457720 645108
rect 322716 645068 457720 645096
rect 322716 645056 322722 645068
rect 457714 645056 457720 645068
rect 457772 645056 457778 645108
rect 115382 644988 115388 645040
rect 115440 645028 115446 645040
rect 124582 645028 124588 645040
rect 115440 645000 124588 645028
rect 115440 644988 115446 645000
rect 124582 644988 124588 645000
rect 124640 644988 124646 645040
rect 148778 644988 148784 645040
rect 148836 645028 148842 645040
rect 148836 645000 156552 645028
rect 148836 644988 148842 645000
rect 86402 644920 86408 644972
rect 86460 644960 86466 644972
rect 124214 644960 124220 644972
rect 86460 644932 124220 644960
rect 86460 644920 86466 644932
rect 124214 644920 124220 644932
rect 124272 644920 124278 644972
rect 148962 644920 148968 644972
rect 149020 644960 149026 644972
rect 156414 644960 156420 644972
rect 149020 644932 156420 644960
rect 149020 644920 149026 644932
rect 156414 644920 156420 644932
rect 156472 644920 156478 644972
rect 94774 644852 94780 644904
rect 94832 644892 94838 644904
rect 120902 644892 120908 644904
rect 94832 644864 120908 644892
rect 94832 644852 94838 644864
rect 120902 644852 120908 644864
rect 120960 644852 120966 644904
rect 147582 644852 147588 644904
rect 147640 644892 147646 644904
rect 155218 644892 155224 644904
rect 147640 644864 155224 644892
rect 147640 644852 147646 644864
rect 155218 644852 155224 644864
rect 155276 644852 155282 644904
rect 156524 644892 156552 645000
rect 156690 644988 156696 645040
rect 156748 645028 156754 645040
rect 207658 645028 207664 645040
rect 156748 645000 207664 645028
rect 156748 644988 156754 645000
rect 207658 644988 207664 645000
rect 207716 644988 207722 645040
rect 226426 644988 226432 645040
rect 226484 645028 226490 645040
rect 300302 645028 300308 645040
rect 226484 645000 300308 645028
rect 226484 644988 226490 645000
rect 300302 644988 300308 645000
rect 300360 644988 300366 645040
rect 314102 644988 314108 645040
rect 314160 645028 314166 645040
rect 456978 645028 456984 645040
rect 314160 645000 456984 645028
rect 314160 644988 314166 645000
rect 456978 644988 456984 645000
rect 457036 644988 457042 645040
rect 156598 644920 156604 644972
rect 156656 644960 156662 644972
rect 172882 644960 172888 644972
rect 156656 644932 172888 644960
rect 156656 644920 156662 644932
rect 172882 644920 172888 644932
rect 172940 644920 172946 644972
rect 214282 644920 214288 644972
rect 214340 644960 214346 644972
rect 289262 644960 289268 644972
rect 214340 644932 289268 644960
rect 214340 644920 214346 644932
rect 289262 644920 289268 644932
rect 289320 644920 289326 644972
rect 318058 644920 318064 644972
rect 318116 644960 318122 644972
rect 471606 644960 471612 644972
rect 318116 644932 471612 644960
rect 318116 644920 318122 644932
rect 471606 644920 471612 644932
rect 471664 644920 471670 644972
rect 176102 644892 176108 644904
rect 156524 644864 176108 644892
rect 176102 644852 176108 644864
rect 176160 644852 176166 644904
rect 232498 644852 232504 644904
rect 232556 644892 232562 644904
rect 271966 644892 271972 644904
rect 232556 644864 271972 644892
rect 232556 644852 232562 644864
rect 271966 644852 271972 644864
rect 272024 644852 272030 644904
rect 304258 644852 304264 644904
rect 304316 644892 304322 644904
rect 457622 644892 457628 644904
rect 304316 644864 457628 644892
rect 304316 644852 304322 644864
rect 457622 644852 457628 644864
rect 457680 644852 457686 644904
rect 106366 644784 106372 644836
rect 106424 644824 106430 644836
rect 121638 644824 121644 644836
rect 106424 644796 121644 644824
rect 106424 644784 106430 644796
rect 121638 644784 121644 644796
rect 121696 644784 121702 644836
rect 143350 644784 143356 644836
rect 143408 644824 143414 644836
rect 184474 644824 184480 644836
rect 143408 644796 184480 644824
rect 143408 644784 143414 644796
rect 184474 644784 184480 644796
rect 184532 644784 184538 644836
rect 231118 644784 231124 644836
rect 231176 644824 231182 644836
rect 248782 644824 248788 644836
rect 231176 644796 248788 644824
rect 231176 644784 231182 644796
rect 248782 644784 248788 644796
rect 248840 644784 248846 644836
rect 249150 644784 249156 644836
rect 249208 644824 249214 644836
rect 295518 644824 295524 644836
rect 249208 644796 295524 644824
rect 249208 644784 249214 644796
rect 295518 644784 295524 644796
rect 295576 644784 295582 644836
rect 314010 644784 314016 644836
rect 314068 644824 314074 644836
rect 483198 644824 483204 644836
rect 314068 644796 483204 644824
rect 314068 644784 314074 644796
rect 483198 644784 483204 644796
rect 483256 644784 483262 644836
rect 109586 644716 109592 644768
rect 109644 644756 109650 644768
rect 126974 644756 126980 644768
rect 109644 644728 126980 644756
rect 109644 644716 109650 644728
rect 126974 644716 126980 644728
rect 127032 644716 127038 644768
rect 149698 644716 149704 644768
rect 149756 644756 149762 644768
rect 190454 644756 190460 644768
rect 149756 644728 190460 644756
rect 149756 644716 149762 644728
rect 190454 644716 190460 644728
rect 190512 644716 190518 644768
rect 222930 644716 222936 644768
rect 222988 644756 222994 644768
rect 277670 644756 277676 644768
rect 222988 644728 277676 644756
rect 222988 644716 222994 644728
rect 277670 644716 277676 644728
rect 277728 644716 277734 644768
rect 319622 644716 319628 644768
rect 319680 644756 319686 644768
rect 511994 644756 512000 644768
rect 319680 644728 512000 644756
rect 319680 644716 319686 644728
rect 511994 644716 512000 644728
rect 512052 644716 512058 644768
rect 55122 644648 55128 644700
rect 55180 644688 55186 644700
rect 80606 644688 80612 644700
rect 55180 644660 80612 644688
rect 55180 644648 55186 644660
rect 80606 644648 80612 644660
rect 80664 644648 80670 644700
rect 103790 644648 103796 644700
rect 103848 644688 103854 644700
rect 121454 644688 121460 644700
rect 103848 644660 121460 644688
rect 103848 644648 103854 644660
rect 121454 644648 121460 644660
rect 121512 644648 121518 644700
rect 149790 644648 149796 644700
rect 149848 644688 149854 644700
rect 199286 644688 199292 644700
rect 149848 644660 199292 644688
rect 149848 644648 149854 644660
rect 199286 644648 199292 644660
rect 199344 644648 199350 644700
rect 239674 644648 239680 644700
rect 239732 644688 239738 644700
rect 297726 644688 297732 644700
rect 239732 644660 297732 644688
rect 239732 644648 239738 644660
rect 297726 644648 297732 644660
rect 297784 644648 297790 644700
rect 316954 644648 316960 644700
rect 317012 644688 317018 644700
rect 512086 644688 512092 644700
rect 317012 644660 512092 644688
rect 317012 644648 317018 644660
rect 512086 644648 512092 644660
rect 512144 644648 512150 644700
rect 54938 644580 54944 644632
rect 54996 644620 55002 644632
rect 92198 644620 92204 644632
rect 54996 644592 92204 644620
rect 54996 644580 55002 644592
rect 92198 644580 92204 644592
rect 92256 644580 92262 644632
rect 100570 644580 100576 644632
rect 100628 644620 100634 644632
rect 124398 644620 124404 644632
rect 100628 644592 124404 644620
rect 100628 644580 100634 644592
rect 124398 644580 124404 644592
rect 124456 644580 124462 644632
rect 148870 644580 148876 644632
rect 148928 644620 148934 644632
rect 148928 644592 161474 644620
rect 148928 644580 148934 644592
rect 55030 644512 55036 644564
rect 55088 644552 55094 644564
rect 88978 644552 88984 644564
rect 55088 644524 88984 644552
rect 55088 644512 55094 644524
rect 88978 644512 88984 644524
rect 89036 644512 89042 644564
rect 112162 644512 112168 644564
rect 112220 644552 112226 644564
rect 120994 644552 121000 644564
rect 112220 644524 121000 644552
rect 112220 644512 112226 644524
rect 120994 644512 121000 644524
rect 121052 644512 121058 644564
rect 148410 644512 148416 644564
rect 148468 644552 148474 644564
rect 153194 644552 153200 644564
rect 148468 644524 153200 644552
rect 148468 644512 148474 644524
rect 153194 644512 153200 644524
rect 153252 644512 153258 644564
rect 155218 644512 155224 644564
rect 155276 644552 155282 644564
rect 158714 644552 158720 644564
rect 155276 644524 158720 644552
rect 155276 644512 155282 644524
rect 158714 644512 158720 644524
rect 158772 644512 158778 644564
rect 161446 644552 161474 644592
rect 239582 644580 239588 644632
rect 239640 644620 239646 644632
rect 251358 644620 251364 644632
rect 239640 644592 251364 644620
rect 239640 644580 239646 644592
rect 251358 644580 251364 644592
rect 251416 644580 251422 644632
rect 317046 644580 317052 644632
rect 317104 644620 317110 644632
rect 512178 644620 512184 644632
rect 317104 644592 512184 644620
rect 317104 644580 317110 644592
rect 512178 644580 512184 644592
rect 512236 644580 512242 644632
rect 201862 644552 201868 644564
rect 161446 644524 201868 644552
rect 201862 644512 201868 644524
rect 201920 644512 201926 644564
rect 237466 644512 237472 644564
rect 237524 644552 237530 644564
rect 254486 644552 254492 644564
rect 237524 644524 254492 644552
rect 237524 644512 237530 644524
rect 254486 644512 254492 644524
rect 254544 644512 254550 644564
rect 305638 644512 305644 644564
rect 305696 644552 305702 644564
rect 501230 644552 501236 644564
rect 305696 644524 501236 644552
rect 305696 644512 305702 644524
rect 501230 644512 501236 644524
rect 501288 644512 501294 644564
rect 59354 644444 59360 644496
rect 59412 644484 59418 644496
rect 97994 644484 98000 644496
rect 59412 644456 98000 644484
rect 59412 644444 59418 644456
rect 97994 644444 98000 644456
rect 98052 644444 98058 644496
rect 117958 644444 117964 644496
rect 118016 644484 118022 644496
rect 124490 644484 124496 644496
rect 118016 644456 124496 644484
rect 118016 644444 118022 644456
rect 124490 644444 124496 644456
rect 124548 644444 124554 644496
rect 134058 644444 134064 644496
rect 134116 644484 134122 644496
rect 149974 644484 149980 644496
rect 134116 644456 149980 644484
rect 134116 644444 134122 644456
rect 149974 644444 149980 644456
rect 150032 644444 150038 644496
rect 205542 644444 205548 644496
rect 205600 644484 205606 644496
rect 211154 644484 211160 644496
rect 205600 644456 211160 644484
rect 205600 644444 205606 644456
rect 211154 644444 211160 644456
rect 211212 644444 211218 644496
rect 239490 644444 239496 644496
rect 239548 644484 239554 644496
rect 242894 644484 242900 644496
rect 239548 644456 242900 644484
rect 239548 644444 239554 644456
rect 242894 644444 242900 644456
rect 242952 644444 242958 644496
rect 3418 643696 3424 643748
rect 3476 643736 3482 643748
rect 321002 643736 321008 643748
rect 3476 643708 321008 643736
rect 3476 643696 3482 643708
rect 321002 643696 321008 643708
rect 321060 643696 321066 643748
rect 238110 643560 238116 643612
rect 238168 643600 238174 643612
rect 268654 643600 268660 643612
rect 238168 643572 268660 643600
rect 238168 643560 238174 643572
rect 268654 643560 268660 643572
rect 268712 643560 268718 643612
rect 126238 643492 126244 643544
rect 126296 643532 126302 643544
rect 187694 643532 187700 643544
rect 126296 643504 187700 643532
rect 126296 643492 126302 643504
rect 187694 643492 187700 643504
rect 187752 643492 187758 643544
rect 220078 643492 220084 643544
rect 220136 643532 220142 643544
rect 257062 643532 257068 643544
rect 220136 643504 257068 643532
rect 220136 643492 220142 643504
rect 257062 643492 257068 643504
rect 257120 643492 257126 643544
rect 149882 643424 149888 643476
rect 149940 643464 149946 643476
rect 170306 643464 170312 643476
rect 149940 643436 170312 643464
rect 149940 643424 149946 643436
rect 170306 643424 170312 643436
rect 170364 643424 170370 643476
rect 228358 643424 228364 643476
rect 228416 643464 228422 643476
rect 266538 643464 266544 643476
rect 228416 643436 266544 643464
rect 228416 643424 228422 643436
rect 266538 643424 266544 643436
rect 266596 643424 266602 643476
rect 56318 643356 56324 643408
rect 56376 643396 56382 643408
rect 71590 643396 71596 643408
rect 56376 643368 71596 643396
rect 56376 643356 56382 643368
rect 71590 643356 71596 643368
rect 71648 643356 71654 643408
rect 141878 643356 141884 643408
rect 141936 643396 141942 643408
rect 167086 643396 167092 643408
rect 141936 643368 167092 643396
rect 141936 643356 141942 643368
rect 167086 643356 167092 643368
rect 167144 643356 167150 643408
rect 220170 643356 220176 643408
rect 220228 643396 220234 643408
rect 260374 643396 260380 643408
rect 220228 643368 260380 643396
rect 220228 643356 220234 643368
rect 260374 643356 260380 643368
rect 260432 643356 260438 643408
rect 56502 643288 56508 643340
rect 56560 643328 56566 643340
rect 65794 643328 65800 643340
rect 56560 643300 65800 643328
rect 56560 643288 56566 643300
rect 65794 643288 65800 643300
rect 65852 643288 65858 643340
rect 137646 643288 137652 643340
rect 137704 643328 137710 643340
rect 179000 643328 179006 643340
rect 137704 643300 179006 643328
rect 137704 643288 137710 643300
rect 179000 643288 179006 643300
rect 179058 643288 179064 643340
rect 231210 643288 231216 643340
rect 231268 643328 231274 643340
rect 280246 643328 280252 643340
rect 231268 643300 280252 643328
rect 231268 643288 231274 643300
rect 280246 643288 280252 643300
rect 280304 643288 280310 643340
rect 59262 643220 59268 643272
rect 59320 643260 59326 643272
rect 74810 643260 74816 643272
rect 59320 643232 74816 643260
rect 59320 643220 59326 643232
rect 74810 643220 74816 643232
rect 74868 643220 74874 643272
rect 144178 643220 144184 643272
rect 144236 643260 144242 643272
rect 193812 643260 193818 643272
rect 144236 643232 193818 643260
rect 144236 643220 144242 643232
rect 193812 643220 193818 643232
rect 193870 643220 193876 643272
rect 236638 643220 236644 643272
rect 236696 643260 236702 643272
rect 291838 643260 291844 643272
rect 236696 643232 291844 643260
rect 236696 643220 236702 643232
rect 291838 643220 291844 643232
rect 291896 643220 291902 643272
rect 56410 643152 56416 643204
rect 56468 643192 56474 643204
rect 77386 643192 77392 643204
rect 56468 643164 77392 643192
rect 56468 643152 56474 643164
rect 77386 643152 77392 643164
rect 77444 643152 77450 643204
rect 83182 643152 83188 643204
rect 83240 643192 83246 643204
rect 124306 643192 124312 643204
rect 83240 643164 124312 643192
rect 83240 643152 83246 643164
rect 124306 643152 124312 643164
rect 124364 643152 124370 643204
rect 125410 643152 125416 643204
rect 125468 643192 125474 643204
rect 182220 643192 182226 643204
rect 125468 643164 182226 643192
rect 125468 643152 125474 643164
rect 182220 643152 182226 643164
rect 182278 643152 182284 643204
rect 215938 643152 215944 643204
rect 215996 643192 216002 643204
rect 274634 643192 274640 643204
rect 215996 643164 274640 643192
rect 215996 643152 216002 643164
rect 274634 643152 274640 643164
rect 274692 643152 274698 643204
rect 69290 643084 69296 643136
rect 69348 643124 69354 643136
rect 122834 643124 122840 643136
rect 69348 643096 122840 643124
rect 69348 643084 69354 643096
rect 122834 643084 122840 643096
rect 122892 643084 122898 643136
rect 146110 643084 146116 643136
rect 146168 643124 146174 643136
rect 155494 643124 155500 643136
rect 146168 643096 155500 643124
rect 146168 643084 146174 643096
rect 155494 643084 155500 643096
rect 155552 643084 155558 643136
rect 217318 643084 217324 643136
rect 217376 643124 217382 643136
rect 286134 643124 286140 643136
rect 217376 643096 286140 643124
rect 217376 643084 217382 643096
rect 286134 643084 286140 643096
rect 286192 643084 286198 643136
rect 312538 643084 312544 643136
rect 312596 643124 312602 643136
rect 321554 643124 321560 643136
rect 312596 643096 321560 643124
rect 312596 643084 312602 643096
rect 321554 643084 321560 643096
rect 321612 643084 321618 643136
rect 54846 642336 54852 642388
rect 54904 642376 54910 642388
rect 62942 642376 62948 642388
rect 54904 642348 62948 642376
rect 54904 642336 54910 642348
rect 62942 642336 62948 642348
rect 63000 642336 63006 642388
rect 223574 642336 223580 642388
rect 223632 642376 223638 642388
rect 249150 642376 249156 642388
rect 223632 642348 249156 642376
rect 223632 642336 223638 642348
rect 249150 642336 249156 642348
rect 249208 642336 249214 642388
rect 262950 642376 262956 642388
rect 258046 642348 262956 642376
rect 222838 641860 222844 641912
rect 222896 641900 222902 641912
rect 258046 641900 258074 642348
rect 262950 642336 262956 642348
rect 263008 642336 263014 642388
rect 283558 642376 283564 642388
rect 277366 642348 283564 642376
rect 222896 641872 258074 641900
rect 222896 641860 222902 641872
rect 214558 641792 214564 641844
rect 214616 641832 214622 641844
rect 277366 641832 277394 642348
rect 283558 642336 283564 642348
rect 283616 642336 283622 642388
rect 214616 641804 277394 641832
rect 214616 641792 214622 641804
rect 57882 641724 57888 641776
rect 57940 641764 57946 641776
rect 146202 641764 146208 641776
rect 57940 641736 146208 641764
rect 57940 641724 57946 641736
rect 146202 641724 146208 641736
rect 146260 641764 146266 641776
rect 238018 641764 238024 641776
rect 146260 641736 238024 641764
rect 146260 641724 146266 641736
rect 238018 641724 238024 641736
rect 238076 641724 238082 641776
rect 140038 640296 140044 640348
rect 140096 640336 140102 640348
rect 146294 640336 146300 640348
rect 140096 640308 146300 640336
rect 140096 640296 140102 640308
rect 146294 640296 146300 640308
rect 146352 640296 146358 640348
rect 235258 640296 235264 640348
rect 235316 640336 235322 640348
rect 237374 640336 237380 640348
rect 235316 640308 237380 640336
rect 235316 640296 235322 640308
rect 237374 640296 237380 640308
rect 237432 640296 237438 640348
rect 465166 640296 465172 640348
rect 465224 640336 465230 640348
rect 580258 640336 580264 640348
rect 465224 640308 580264 640336
rect 465224 640296 465230 640308
rect 580258 640296 580264 640308
rect 580316 640296 580322 640348
rect 309870 638936 309876 638988
rect 309928 638976 309934 638988
rect 321554 638976 321560 638988
rect 309928 638948 321560 638976
rect 309928 638936 309934 638948
rect 321554 638936 321560 638948
rect 321612 638936 321618 638988
rect 238938 638596 238944 638648
rect 238996 638636 239002 638648
rect 239766 638636 239772 638648
rect 238996 638608 239772 638636
rect 238996 638596 239002 638608
rect 239766 638596 239772 638608
rect 239824 638596 239830 638648
rect 215754 638188 215760 638240
rect 215812 638228 215818 638240
rect 237466 638228 237472 638240
rect 215812 638200 237472 638228
rect 215812 638188 215818 638200
rect 237466 638188 237472 638200
rect 237524 638188 237530 638240
rect 233602 633428 233608 633480
rect 233660 633468 233666 633480
rect 237374 633468 237380 633480
rect 233660 633440 237380 633468
rect 233660 633428 233666 633440
rect 237374 633428 237380 633440
rect 237432 633428 237438 633480
rect 307110 633428 307116 633480
rect 307168 633468 307174 633480
rect 321554 633468 321560 633480
rect 307168 633440 321560 633468
rect 307168 633428 307174 633440
rect 321554 633428 321560 633440
rect 321612 633428 321618 633480
rect 141234 630640 141240 630692
rect 141292 630680 141298 630692
rect 146294 630680 146300 630692
rect 141292 630652 146300 630680
rect 141292 630640 141298 630652
rect 146294 630640 146300 630652
rect 146352 630640 146358 630692
rect 232590 630640 232596 630692
rect 232648 630680 232654 630692
rect 237374 630680 237380 630692
rect 232648 630652 237380 630680
rect 232648 630640 232654 630652
rect 237374 630640 237380 630652
rect 237432 630640 237438 630692
rect 309778 629280 309784 629332
rect 309836 629320 309842 629332
rect 321554 629320 321560 629332
rect 309836 629292 321560 629320
rect 309836 629280 309842 629292
rect 321554 629280 321560 629292
rect 321612 629280 321618 629332
rect 132586 627920 132592 627972
rect 132644 627960 132650 627972
rect 146294 627960 146300 627972
rect 132644 627932 146300 627960
rect 132644 627920 132650 627932
rect 146294 627920 146300 627932
rect 146352 627920 146358 627972
rect 224310 625132 224316 625184
rect 224368 625172 224374 625184
rect 237374 625172 237380 625184
rect 224368 625144 237380 625172
rect 224368 625132 224374 625144
rect 237374 625132 237380 625144
rect 237432 625132 237438 625184
rect 305730 625132 305736 625184
rect 305788 625172 305794 625184
rect 321554 625172 321560 625184
rect 305788 625144 321560 625172
rect 305788 625132 305794 625144
rect 321554 625132 321560 625144
rect 321612 625132 321618 625184
rect 218606 620984 218612 621036
rect 218664 621024 218670 621036
rect 237374 621024 237380 621036
rect 218664 620996 237380 621024
rect 218664 620984 218670 620996
rect 237374 620984 237380 620996
rect 237432 620984 237438 621036
rect 312630 619624 312636 619676
rect 312688 619664 312694 619676
rect 321554 619664 321560 619676
rect 312688 619636 321560 619664
rect 312688 619624 312694 619636
rect 321554 619624 321560 619636
rect 321612 619624 321618 619676
rect 314194 615476 314200 615528
rect 314252 615516 314258 615528
rect 321554 615516 321560 615528
rect 314252 615488 321560 615516
rect 314252 615476 314258 615488
rect 321554 615476 321560 615488
rect 321612 615476 321618 615528
rect 233878 612756 233884 612808
rect 233936 612796 233942 612808
rect 237374 612796 237380 612808
rect 233936 612768 237380 612796
rect 233936 612756 233942 612768
rect 237374 612756 237380 612768
rect 237432 612756 237438 612808
rect 129090 609968 129096 610020
rect 129148 610008 129154 610020
rect 146294 610008 146300 610020
rect 129148 609980 146300 610008
rect 129148 609968 129154 609980
rect 146294 609968 146300 609980
rect 146352 609968 146358 610020
rect 217410 609968 217416 610020
rect 217468 610008 217474 610020
rect 237374 610008 237380 610020
rect 217468 609980 237380 610008
rect 217468 609968 217474 609980
rect 237374 609968 237380 609980
rect 237432 609968 237438 610020
rect 311250 609968 311256 610020
rect 311308 610008 311314 610020
rect 321554 610008 321560 610020
rect 311308 609980 321560 610008
rect 311308 609968 311314 609980
rect 321554 609968 321560 609980
rect 321612 609968 321618 610020
rect 302786 609220 302792 609272
rect 302844 609260 302850 609272
rect 303154 609260 303160 609272
rect 302844 609232 303160 609260
rect 302844 609220 302850 609232
rect 303154 609220 303160 609232
rect 303212 609260 303218 609272
rect 322658 609260 322664 609272
rect 303212 609232 322664 609260
rect 303212 609220 303218 609232
rect 322658 609220 322664 609232
rect 322716 609220 322722 609272
rect 124030 608608 124036 608660
rect 124088 608648 124094 608660
rect 145558 608648 145564 608660
rect 124088 608620 145564 608648
rect 124088 608608 124094 608620
rect 145558 608608 145564 608620
rect 145616 608608 145622 608660
rect 220262 607180 220268 607232
rect 220320 607220 220326 607232
rect 237374 607220 237380 607232
rect 220320 607192 237380 607220
rect 220320 607180 220326 607192
rect 237374 607180 237380 607192
rect 237432 607180 237438 607232
rect 229738 603100 229744 603152
rect 229796 603140 229802 603152
rect 237374 603140 237380 603152
rect 229796 603112 237380 603140
rect 229796 603100 229802 603112
rect 237374 603100 237380 603112
rect 237432 603100 237438 603152
rect 232866 600312 232872 600364
rect 232924 600352 232930 600364
rect 237374 600352 237380 600364
rect 232924 600324 237380 600352
rect 232924 600312 232930 600324
rect 237374 600312 237380 600324
rect 237432 600312 237438 600364
rect 308398 600312 308404 600364
rect 308456 600352 308462 600364
rect 321554 600352 321560 600364
rect 308456 600324 321560 600352
rect 308456 600312 308462 600324
rect 321554 600312 321560 600324
rect 321612 600312 321618 600364
rect 126882 597524 126888 597576
rect 126940 597564 126946 597576
rect 146294 597564 146300 597576
rect 126940 597536 146300 597564
rect 126940 597524 126946 597536
rect 146294 597524 146300 597536
rect 146352 597524 146358 597576
rect 235350 597524 235356 597576
rect 235408 597564 235414 597576
rect 237374 597564 237380 597576
rect 235408 597536 237380 597564
rect 235408 597524 235414 597536
rect 237374 597524 237380 597536
rect 237432 597524 237438 597576
rect 305822 596164 305828 596216
rect 305880 596204 305886 596216
rect 321554 596204 321560 596216
rect 305880 596176 321560 596204
rect 305880 596164 305886 596176
rect 321554 596164 321560 596176
rect 321612 596164 321618 596216
rect 144270 594804 144276 594856
rect 144328 594844 144334 594856
rect 146938 594844 146944 594856
rect 144328 594816 146944 594844
rect 144328 594804 144334 594816
rect 146938 594804 146944 594816
rect 146996 594804 147002 594856
rect 216030 594804 216036 594856
rect 216088 594844 216094 594856
rect 237374 594844 237380 594856
rect 216088 594816 237380 594844
rect 216088 594804 216094 594816
rect 237374 594804 237380 594816
rect 237432 594804 237438 594856
rect 513282 592016 513288 592068
rect 513340 592056 513346 592068
rect 578878 592056 578884 592068
rect 513340 592028 578884 592056
rect 513340 592016 513346 592028
rect 578878 592016 578884 592028
rect 578936 592016 578942 592068
rect 139762 590656 139768 590708
rect 139820 590696 139826 590708
rect 146294 590696 146300 590708
rect 139820 590668 146300 590696
rect 139820 590656 139826 590668
rect 146294 590656 146300 590668
rect 146352 590656 146358 590708
rect 217502 590656 217508 590708
rect 217560 590696 217566 590708
rect 237374 590696 237380 590708
rect 217560 590668 237380 590696
rect 217560 590656 217566 590668
rect 237374 590656 237380 590668
rect 237432 590656 237438 590708
rect 317138 590656 317144 590708
rect 317196 590696 317202 590708
rect 321554 590696 321560 590708
rect 317196 590668 321560 590696
rect 317196 590656 317202 590668
rect 321554 590656 321560 590668
rect 321612 590656 321618 590708
rect 227162 587868 227168 587920
rect 227220 587908 227226 587920
rect 237374 587908 237380 587920
rect 227220 587880 237380 587908
rect 227220 587868 227226 587880
rect 237374 587868 237380 587880
rect 237432 587868 237438 587920
rect 219250 585148 219256 585200
rect 219308 585188 219314 585200
rect 237374 585188 237380 585200
rect 219308 585160 237380 585188
rect 219308 585148 219314 585160
rect 237374 585148 237380 585160
rect 237432 585148 237438 585200
rect 123110 584944 123116 584996
rect 123168 584984 123174 584996
rect 123570 584984 123576 584996
rect 123168 584956 123576 584984
rect 123168 584944 123174 584956
rect 123570 584944 123576 584956
rect 123628 584944 123634 584996
rect 148318 583040 148324 583092
rect 148376 583080 148382 583092
rect 148778 583080 148784 583092
rect 148376 583052 148784 583080
rect 148376 583040 148382 583052
rect 148778 583040 148784 583052
rect 148836 583040 148842 583092
rect 148778 582904 148784 582956
rect 148836 582944 148842 582956
rect 148962 582944 148968 582956
rect 148836 582916 148968 582944
rect 148836 582904 148842 582916
rect 148962 582904 148968 582916
rect 149020 582904 149026 582956
rect 223482 582360 223488 582412
rect 223540 582400 223546 582412
rect 237374 582400 237380 582412
rect 223540 582372 237380 582400
rect 223540 582360 223546 582372
rect 237374 582360 237380 582372
rect 237432 582360 237438 582412
rect 120718 581748 120724 581800
rect 120776 581788 120782 581800
rect 121178 581788 121184 581800
rect 120776 581760 121184 581788
rect 120776 581748 120782 581760
rect 121178 581748 121184 581760
rect 121236 581748 121242 581800
rect 57422 581204 57428 581256
rect 57480 581244 57486 581256
rect 59906 581244 59912 581256
rect 57480 581216 59912 581244
rect 57480 581204 57486 581216
rect 59906 581204 59912 581216
rect 59964 581204 59970 581256
rect 3142 580932 3148 580984
rect 3200 580972 3206 580984
rect 305822 580972 305828 580984
rect 3200 580944 305828 580972
rect 3200 580932 3206 580944
rect 305822 580932 305828 580944
rect 305880 580932 305886 580984
rect 145558 580864 145564 580916
rect 145616 580904 145622 580916
rect 213914 580904 213920 580916
rect 145616 580876 213920 580904
rect 145616 580864 145622 580876
rect 213914 580864 213920 580876
rect 213972 580904 213978 580916
rect 302786 580904 302792 580916
rect 213972 580876 302792 580904
rect 213972 580864 213978 580876
rect 302786 580864 302792 580876
rect 302844 580864 302850 580916
rect 58802 580660 58808 580712
rect 58860 580700 58866 580712
rect 60918 580700 60924 580712
rect 58860 580672 60924 580700
rect 58860 580660 58866 580672
rect 60918 580660 60924 580672
rect 60976 580660 60982 580712
rect 119338 580660 119344 580712
rect 119396 580700 119402 580712
rect 123110 580700 123116 580712
rect 119396 580672 123116 580700
rect 119396 580660 119402 580672
rect 123110 580660 123116 580672
rect 123168 580660 123174 580712
rect 147122 580660 147128 580712
rect 147180 580700 147186 580712
rect 151078 580700 151084 580712
rect 147180 580672 151084 580700
rect 147180 580660 147186 580672
rect 151078 580660 151084 580672
rect 151136 580660 151142 580712
rect 57330 580592 57336 580644
rect 57388 580632 57394 580644
rect 61378 580632 61384 580644
rect 57388 580604 61384 580632
rect 57388 580592 57394 580604
rect 61378 580592 61384 580604
rect 61436 580592 61442 580644
rect 112530 580252 112536 580304
rect 112588 580292 112594 580304
rect 123570 580292 123576 580304
rect 112588 580264 123576 580292
rect 112588 580252 112594 580264
rect 123570 580252 123576 580264
rect 123628 580252 123634 580304
rect 199378 580252 199384 580304
rect 199436 580292 199442 580304
rect 212626 580292 212632 580304
rect 199436 580264 212632 580292
rect 199436 580252 199442 580264
rect 212626 580252 212632 580264
rect 212684 580252 212690 580304
rect 59170 579572 59176 579624
rect 59228 579612 59234 579624
rect 62390 579612 62396 579624
rect 59228 579584 62396 579612
rect 59228 579572 59234 579584
rect 62390 579572 62396 579584
rect 62448 579572 62454 579624
rect 148594 579572 148600 579624
rect 148652 579612 148658 579624
rect 150526 579612 150532 579624
rect 148652 579584 150532 579612
rect 148652 579572 148658 579584
rect 150526 579572 150532 579584
rect 150584 579572 150590 579624
rect 295242 579572 295248 579624
rect 295300 579612 295306 579624
rect 319622 579612 319628 579624
rect 295300 579584 319628 579612
rect 295300 579572 295306 579584
rect 319622 579572 319628 579584
rect 319680 579572 319686 579624
rect 289538 579504 289544 579556
rect 289596 579544 289602 579556
rect 316862 579544 316868 579556
rect 289596 579516 316868 579544
rect 289596 579504 289602 579516
rect 316862 579504 316868 579516
rect 316920 579504 316926 579556
rect 107562 579436 107568 579488
rect 107620 579476 107626 579488
rect 124582 579476 124588 579488
rect 107620 579448 124588 579476
rect 107620 579436 107626 579448
rect 124582 579436 124588 579448
rect 124640 579436 124646 579488
rect 288802 579436 288808 579488
rect 288860 579476 288866 579488
rect 317046 579476 317052 579488
rect 288860 579448 317052 579476
rect 288860 579436 288866 579448
rect 317046 579436 317052 579448
rect 317104 579436 317110 579488
rect 97442 579368 97448 579420
rect 97500 579408 97506 579420
rect 120994 579408 121000 579420
rect 97500 579380 121000 579408
rect 97500 579368 97506 579380
rect 120994 579368 121000 579380
rect 121052 579368 121058 579420
rect 288066 579368 288072 579420
rect 288124 579408 288130 579420
rect 316954 579408 316960 579420
rect 288124 579380 316960 579408
rect 288124 579368 288130 579380
rect 316954 579368 316960 579380
rect 317012 579368 317018 579420
rect 98178 579300 98184 579352
rect 98236 579340 98242 579352
rect 126974 579340 126980 579352
rect 98236 579312 126980 579340
rect 98236 579300 98242 579312
rect 126974 579300 126980 579312
rect 127032 579300 127038 579352
rect 148870 579300 148876 579352
rect 148928 579340 148934 579352
rect 155494 579340 155500 579352
rect 148928 579312 155500 579340
rect 148928 579300 148934 579312
rect 155494 579300 155500 579312
rect 155552 579300 155558 579352
rect 286318 579300 286324 579352
rect 286376 579340 286382 579352
rect 319438 579340 319444 579352
rect 286376 579312 319444 579340
rect 286376 579300 286382 579312
rect 319438 579300 319444 579312
rect 319496 579300 319502 579352
rect 93946 579232 93952 579284
rect 94004 579272 94010 579284
rect 124398 579272 124404 579284
rect 94004 579244 124404 579272
rect 94004 579232 94010 579244
rect 124398 579232 124404 579244
rect 124456 579232 124462 579284
rect 149790 579232 149796 579284
rect 149848 579272 149854 579284
rect 156230 579272 156236 579284
rect 149848 579244 156236 579272
rect 149848 579232 149854 579244
rect 156230 579232 156236 579244
rect 156288 579232 156294 579284
rect 165522 579232 165528 579284
rect 165580 579272 165586 579284
rect 211154 579272 211160 579284
rect 165580 579244 211160 579272
rect 165580 579232 165586 579244
rect 211154 579232 211160 579244
rect 211212 579232 211218 579284
rect 258718 579232 258724 579284
rect 258776 579272 258782 579284
rect 322474 579272 322480 579284
rect 258776 579244 322480 579272
rect 258776 579232 258782 579244
rect 322474 579232 322480 579244
rect 322532 579232 322538 579284
rect 58434 579164 58440 579216
rect 58492 579204 58498 579216
rect 68830 579204 68836 579216
rect 58492 579176 68836 579204
rect 58492 579164 58498 579176
rect 68830 579164 68836 579176
rect 68888 579164 68894 579216
rect 87414 579164 87420 579216
rect 87472 579204 87478 579216
rect 121638 579204 121644 579216
rect 87472 579176 121644 579204
rect 87472 579164 87478 579176
rect 121638 579164 121644 579176
rect 121696 579164 121702 579216
rect 123110 579164 123116 579216
rect 123168 579204 123174 579216
rect 211706 579204 211712 579216
rect 123168 579176 211712 579204
rect 123168 579164 123174 579176
rect 211706 579164 211712 579176
rect 211764 579164 211770 579216
rect 245838 579164 245844 579216
rect 245896 579204 245902 579216
rect 322566 579204 322572 579216
rect 245896 579176 322572 579204
rect 245896 579164 245902 579176
rect 322566 579164 322572 579176
rect 322624 579164 322630 579216
rect 57698 579096 57704 579148
rect 57756 579136 57762 579148
rect 71038 579136 71044 579148
rect 57756 579108 71044 579136
rect 57756 579096 57762 579108
rect 71038 579096 71044 579108
rect 71096 579096 71102 579148
rect 88150 579096 88156 579148
rect 88208 579136 88214 579148
rect 124490 579136 124496 579148
rect 88208 579108 124496 579136
rect 88208 579096 88214 579108
rect 124490 579096 124496 579108
rect 124548 579096 124554 579148
rect 148962 579096 148968 579148
rect 149020 579136 149026 579148
rect 159082 579136 159088 579148
rect 149020 579108 159088 579136
rect 149020 579096 149026 579108
rect 159082 579096 159088 579108
rect 159140 579096 159146 579148
rect 200666 579096 200672 579148
rect 200724 579136 200730 579148
rect 301406 579136 301412 579148
rect 200724 579108 301412 579136
rect 200724 579096 200730 579108
rect 301406 579096 301412 579108
rect 301464 579096 301470 579148
rect 57606 579028 57612 579080
rect 57664 579068 57670 579080
rect 83182 579068 83188 579080
rect 57664 579040 83188 579068
rect 57664 579028 57670 579040
rect 83182 579028 83188 579040
rect 83240 579028 83246 579080
rect 84562 579028 84568 579080
rect 84620 579068 84626 579080
rect 122098 579068 122104 579080
rect 84620 579040 122104 579068
rect 84620 579028 84626 579040
rect 122098 579028 122104 579040
rect 122156 579028 122162 579080
rect 148318 579028 148324 579080
rect 148376 579068 148382 579080
rect 161934 579068 161940 579080
rect 148376 579040 161940 579068
rect 148376 579028 148382 579040
rect 161934 579028 161940 579040
rect 161992 579028 161998 579080
rect 196342 579028 196348 579080
rect 196400 579068 196406 579080
rect 302602 579068 302608 579080
rect 196400 579040 302608 579068
rect 196400 579028 196406 579040
rect 302602 579028 302608 579040
rect 302660 579028 302666 579080
rect 66714 578960 66720 579012
rect 66772 579000 66778 579012
rect 120718 579000 120724 579012
rect 66772 578972 120724 579000
rect 66772 578960 66778 578972
rect 120718 578960 120724 578972
rect 120776 578960 120782 579012
rect 148778 578960 148784 579012
rect 148836 579000 148842 579012
rect 164878 579000 164884 579012
rect 148836 578972 164884 579000
rect 148836 578960 148842 578972
rect 164878 578960 164884 578972
rect 164936 578960 164942 579012
rect 184198 578960 184204 579012
rect 184256 579000 184262 579012
rect 301038 579000 301044 579012
rect 184256 578972 301044 579000
rect 184256 578960 184262 578972
rect 301038 578960 301044 578972
rect 301096 578960 301102 579012
rect 63770 578892 63776 578944
rect 63828 578932 63834 578944
rect 122282 578932 122288 578944
rect 63828 578904 122288 578932
rect 63828 578892 63834 578904
rect 122282 578892 122288 578904
rect 122340 578892 122346 578944
rect 149698 578892 149704 578944
rect 149756 578932 149762 578944
rect 151814 578932 151820 578944
rect 149756 578904 151820 578932
rect 149756 578892 149762 578904
rect 151814 578892 151820 578904
rect 151872 578892 151878 578944
rect 179874 578892 179880 578944
rect 179932 578932 179938 578944
rect 301590 578932 301596 578944
rect 179932 578904 301596 578932
rect 179932 578892 179938 578904
rect 301590 578892 301596 578904
rect 301648 578892 301654 578944
rect 147214 578824 147220 578876
rect 147272 578864 147278 578876
rect 166258 578864 166264 578876
rect 147272 578836 166264 578864
rect 147272 578824 147278 578836
rect 166258 578824 166264 578836
rect 166316 578824 166322 578876
rect 290182 578824 290188 578876
rect 290240 578864 290246 578876
rect 314010 578864 314016 578876
rect 290240 578836 314016 578864
rect 290240 578824 290246 578836
rect 314010 578824 314016 578836
rect 314068 578824 314074 578876
rect 297358 578756 297364 578808
rect 297416 578796 297422 578808
rect 319530 578796 319536 578808
rect 297416 578768 319536 578796
rect 297416 578756 297422 578768
rect 319530 578756 319536 578768
rect 319588 578756 319594 578808
rect 292390 578688 292396 578740
rect 292448 578728 292454 578740
rect 314102 578728 314108 578740
rect 292448 578700 314108 578728
rect 292448 578688 292454 578700
rect 314102 578688 314108 578700
rect 314160 578688 314166 578740
rect 106918 578144 106924 578196
rect 106976 578184 106982 578196
rect 108574 578184 108580 578196
rect 106976 578156 108580 578184
rect 106976 578144 106982 578156
rect 108574 578144 108580 578156
rect 108632 578144 108638 578196
rect 116578 578144 116584 578196
rect 116636 578184 116642 578196
rect 117406 578184 117412 578196
rect 116636 578156 117412 578184
rect 116636 578144 116642 578156
rect 117406 578144 117412 578156
rect 117464 578144 117470 578196
rect 191098 578144 191104 578196
rect 191156 578184 191162 578196
rect 195422 578184 195428 578196
rect 191156 578156 195428 578184
rect 191156 578144 191162 578156
rect 195422 578144 195428 578156
rect 195480 578144 195486 578196
rect 192478 578076 192484 578128
rect 192536 578116 192542 578128
rect 198734 578116 198740 578128
rect 192536 578088 198740 578116
rect 192536 578076 192542 578088
rect 198734 578076 198740 578088
rect 198792 578076 198798 578128
rect 174170 577940 174176 577992
rect 174228 577980 174234 577992
rect 189626 577980 189632 577992
rect 174228 577952 189632 577980
rect 174228 577940 174234 577952
rect 189626 577940 189632 577952
rect 189684 577940 189690 577992
rect 162670 577872 162676 577924
rect 162728 577912 162734 577924
rect 178034 577912 178040 577924
rect 162728 577884 178040 577912
rect 162728 577872 162734 577884
rect 178034 577872 178040 577884
rect 178092 577872 178098 577924
rect 164142 577804 164148 577856
rect 164200 577844 164206 577856
rect 183830 577844 183836 577856
rect 164200 577816 183836 577844
rect 164200 577804 164206 577816
rect 183830 577804 183836 577816
rect 183888 577804 183894 577856
rect 227898 577804 227904 577856
rect 227956 577844 227962 577856
rect 265526 577844 265532 577856
rect 227956 577816 265532 577844
rect 227956 577804 227962 577816
rect 265526 577804 265532 577816
rect 265584 577804 265590 577856
rect 77018 577736 77024 577788
rect 77076 577776 77082 577788
rect 86770 577776 86776 577788
rect 77076 577748 86776 577776
rect 77076 577736 77082 577748
rect 86770 577736 86776 577748
rect 86828 577736 86834 577788
rect 94498 577736 94504 577788
rect 94556 577776 94562 577788
rect 104158 577776 104164 577788
rect 94556 577748 104164 577776
rect 94556 577736 94562 577748
rect 104158 577736 104164 577748
rect 104216 577736 104222 577788
rect 150342 577736 150348 577788
rect 150400 577776 150406 577788
rect 151170 577776 151176 577788
rect 150400 577748 151176 577776
rect 150400 577736 150406 577748
rect 151170 577736 151176 577748
rect 151228 577736 151234 577788
rect 154850 577736 154856 577788
rect 154908 577776 154914 577788
rect 181254 577776 181260 577788
rect 154908 577748 181260 577776
rect 154908 577736 154914 577748
rect 181254 577736 181260 577748
rect 181312 577736 181318 577788
rect 232222 577736 232228 577788
rect 232280 577776 232286 577788
rect 279694 577776 279700 577788
rect 232280 577748 279700 577776
rect 232280 577736 232286 577748
rect 279694 577736 279700 577748
rect 279752 577736 279758 577788
rect 60274 577668 60280 577720
rect 60332 577708 60338 577720
rect 71130 577708 71136 577720
rect 60332 577680 71136 577708
rect 60332 577668 60338 577680
rect 71130 577668 71136 577680
rect 71188 577668 71194 577720
rect 75270 577668 75276 577720
rect 75328 577708 75334 577720
rect 96982 577708 96988 577720
rect 75328 577680 96988 577708
rect 75328 577668 75334 577680
rect 96982 577668 96988 577680
rect 97040 577668 97046 577720
rect 100202 577668 100208 577720
rect 100260 577708 100266 577720
rect 115198 577708 115204 577720
rect 100260 577680 115204 577708
rect 100260 577668 100266 577680
rect 115198 577668 115204 577680
rect 115256 577668 115262 577720
rect 159818 577668 159824 577720
rect 159876 577708 159882 577720
rect 192846 577708 192852 577720
rect 159876 577680 192852 577708
rect 159876 577668 159882 577680
rect 192846 577668 192852 577680
rect 192904 577668 192910 577720
rect 197998 577668 198004 577720
rect 198056 577708 198062 577720
rect 210234 577708 210240 577720
rect 198056 577680 210240 577708
rect 198056 577668 198062 577680
rect 210234 577668 210240 577680
rect 210292 577668 210298 577720
rect 220722 577668 220728 577720
rect 220780 577708 220786 577720
rect 268102 577708 268108 577720
rect 220780 577680 268108 577708
rect 220780 577668 220786 577680
rect 268102 577668 268108 577680
rect 268160 577668 268166 577720
rect 273898 577668 273904 577720
rect 273956 577708 273962 577720
rect 282914 577708 282920 577720
rect 273956 577680 282920 577708
rect 273956 577668 273962 577680
rect 282914 577668 282920 577680
rect 282972 577668 282978 577720
rect 289078 577668 289084 577720
rect 289136 577708 289142 577720
rect 300302 577708 300308 577720
rect 289136 577680 300308 577708
rect 289136 577668 289142 577680
rect 300302 577668 300308 577680
rect 300360 577668 300366 577720
rect 58894 577600 58900 577652
rect 58952 577640 58958 577652
rect 74534 577640 74540 577652
rect 58952 577612 74540 577640
rect 58952 577600 58958 577612
rect 74534 577600 74540 577612
rect 74592 577600 74598 577652
rect 86034 577600 86040 577652
rect 86092 577640 86098 577652
rect 108298 577640 108304 577652
rect 86092 577612 108304 577640
rect 86092 577600 86098 577612
rect 108298 577600 108304 577612
rect 108356 577600 108362 577652
rect 116670 577600 116676 577652
rect 116728 577640 116734 577652
rect 120166 577640 120172 577652
rect 116728 577612 120172 577640
rect 116728 577600 116734 577612
rect 120166 577600 120172 577612
rect 120224 577600 120230 577652
rect 130470 577600 130476 577652
rect 130528 577640 130534 577652
rect 163866 577640 163872 577652
rect 130528 577612 163872 577640
rect 130528 577600 130534 577612
rect 163866 577600 163872 577612
rect 163924 577600 163930 577652
rect 169846 577600 169852 577652
rect 169904 577640 169910 577652
rect 175458 577640 175464 577652
rect 169904 577612 175464 577640
rect 169904 577600 169910 577612
rect 175458 577600 175464 577612
rect 175516 577600 175522 577652
rect 183462 577600 183468 577652
rect 183520 577640 183526 577652
rect 232498 577640 232504 577652
rect 183520 577612 232504 577640
rect 183520 577600 183526 577612
rect 232498 577600 232504 577612
rect 232556 577600 232562 577652
rect 235442 577600 235448 577652
rect 235500 577640 235506 577652
rect 242342 577640 242348 577652
rect 235500 577612 242348 577640
rect 235500 577600 235506 577612
rect 242342 577600 242348 577612
rect 242400 577600 242406 577652
rect 249058 577600 249064 577652
rect 249116 577640 249122 577652
rect 259638 577640 259644 577652
rect 249116 577612 259644 577640
rect 249116 577600 249122 577612
rect 259638 577600 259644 577612
rect 259696 577600 259702 577652
rect 280798 577600 280804 577652
rect 280856 577640 280862 577652
rect 296990 577640 296996 577652
rect 280856 577612 296996 577640
rect 280856 577600 280862 577612
rect 296990 577600 296996 577612
rect 297048 577600 297054 577652
rect 68738 577532 68744 577584
rect 68796 577572 68802 577584
rect 105538 577572 105544 577584
rect 68796 577544 105544 577572
rect 68796 577532 68802 577544
rect 105538 577532 105544 577544
rect 105596 577532 105602 577584
rect 133322 577532 133328 577584
rect 133380 577572 133386 577584
rect 187050 577572 187056 577584
rect 133380 577544 187056 577572
rect 133380 577532 133386 577544
rect 187050 577532 187056 577544
rect 187108 577532 187114 577584
rect 195238 577532 195244 577584
rect 195296 577572 195302 577584
rect 212718 577572 212724 577584
rect 195296 577544 212724 577572
rect 195296 577532 195302 577544
rect 212718 577532 212724 577544
rect 212776 577532 212782 577584
rect 222194 577532 222200 577584
rect 222252 577572 222258 577584
rect 273806 577572 273812 577584
rect 222252 577544 273812 577572
rect 222252 577532 222258 577544
rect 273806 577532 273812 577544
rect 273864 577532 273870 577584
rect 280890 577532 280896 577584
rect 280948 577572 280954 577584
rect 322382 577572 322388 577584
rect 280948 577544 322388 577572
rect 280948 577532 280954 577544
rect 322382 577532 322388 577544
rect 322440 577532 322446 577584
rect 71314 577464 71320 577516
rect 71372 577504 71378 577516
rect 108390 577504 108396 577516
rect 71372 577476 108396 577504
rect 71372 577464 71378 577476
rect 108390 577464 108396 577476
rect 108448 577464 108454 577516
rect 110414 577464 110420 577516
rect 110472 577504 110478 577516
rect 121178 577504 121184 577516
rect 110472 577476 121184 577504
rect 110472 577464 110478 577476
rect 121178 577464 121184 577476
rect 121236 577464 121242 577516
rect 134702 577464 134708 577516
rect 134760 577504 134766 577516
rect 207014 577504 207020 577516
rect 134760 577476 207020 577504
rect 134760 577464 134766 577476
rect 207014 577464 207020 577476
rect 207072 577464 207078 577516
rect 217134 577464 217140 577516
rect 217192 577504 217198 577516
rect 223482 577504 223488 577516
rect 217192 577476 223488 577504
rect 217192 577464 217198 577476
rect 223482 577464 223488 577476
rect 223540 577464 223546 577516
rect 231302 577464 231308 577516
rect 231360 577504 231366 577516
rect 239766 577504 239772 577516
rect 231360 577476 239772 577504
rect 231360 577464 231366 577476
rect 239766 577464 239772 577476
rect 239824 577464 239830 577516
rect 257982 577464 257988 577516
rect 258040 577504 258046 577516
rect 324774 577504 324780 577516
rect 258040 577476 324780 577504
rect 258040 577464 258046 577476
rect 324774 577464 324780 577476
rect 324832 577464 324838 577516
rect 202230 577192 202236 577244
rect 202288 577232 202294 577244
rect 204438 577232 204444 577244
rect 202288 577204 204444 577232
rect 202288 577192 202294 577204
rect 204438 577192 204444 577204
rect 204496 577192 204502 577244
rect 269758 577192 269764 577244
rect 269816 577232 269822 577244
rect 271230 577232 271236 577244
rect 269816 577204 271236 577232
rect 269816 577192 269822 577204
rect 271230 577192 271236 577204
rect 271288 577192 271294 577244
rect 242158 576920 242164 576972
rect 242216 576960 242222 576972
rect 248506 576960 248512 576972
rect 242216 576932 248512 576960
rect 242216 576920 242222 576932
rect 248506 576920 248512 576932
rect 248564 576920 248570 576972
rect 64138 576852 64144 576904
rect 64196 576892 64202 576904
rect 64966 576892 64972 576904
rect 64196 576864 64972 576892
rect 64196 576852 64202 576864
rect 64966 576852 64972 576864
rect 65024 576852 65030 576904
rect 199470 576852 199476 576904
rect 199528 576892 199534 576904
rect 201494 576892 201500 576904
rect 199528 576864 201500 576892
rect 199528 576852 199534 576864
rect 201494 576852 201500 576864
rect 201552 576852 201558 576904
rect 244918 576852 244924 576904
rect 244976 576892 244982 576904
rect 250622 576892 250628 576904
rect 244976 576864 250628 576892
rect 244976 576852 244982 576864
rect 250622 576852 250628 576864
rect 250680 576852 250686 576904
rect 282178 576852 282184 576904
rect 282236 576892 282242 576904
rect 288710 576892 288716 576904
rect 282236 576864 288716 576892
rect 282236 576852 282242 576864
rect 288710 576852 288716 576864
rect 288768 576852 288774 576904
rect 160738 576376 160744 576428
rect 160796 576416 160802 576428
rect 212994 576416 213000 576428
rect 160796 576388 213000 576416
rect 160796 576376 160802 576388
rect 212994 576376 213000 576388
rect 213052 576376 213058 576428
rect 122558 576308 122564 576360
rect 122616 576348 122622 576360
rect 211246 576348 211252 576360
rect 122616 576320 211252 576348
rect 122616 576308 122622 576320
rect 211246 576308 211252 576320
rect 211304 576308 211310 576360
rect 228634 576308 228640 576360
rect 228692 576348 228698 576360
rect 300946 576348 300952 576360
rect 228692 576320 300952 576348
rect 228692 576308 228698 576320
rect 300946 576308 300952 576320
rect 301004 576308 301010 576360
rect 57238 576240 57244 576292
rect 57296 576280 57302 576292
rect 79318 576280 79324 576292
rect 57296 576252 79324 576280
rect 57296 576240 57302 576252
rect 79318 576240 79324 576252
rect 79376 576240 79382 576292
rect 91094 576240 91100 576292
rect 91152 576280 91158 576292
rect 96798 576280 96804 576292
rect 91152 576252 96804 576280
rect 91152 576240 91158 576252
rect 96798 576240 96804 576252
rect 96856 576240 96862 576292
rect 100386 576240 100392 576292
rect 100444 576280 100450 576292
rect 123294 576280 123300 576292
rect 100444 576252 123300 576280
rect 100444 576240 100450 576252
rect 123294 576240 123300 576252
rect 123352 576240 123358 576292
rect 206278 576240 206284 576292
rect 206336 576280 206342 576292
rect 302970 576280 302976 576292
rect 206336 576252 302976 576280
rect 206336 576240 206342 576252
rect 302970 576240 302976 576252
rect 303028 576240 303034 576292
rect 65242 576172 65248 576224
rect 65300 576212 65306 576224
rect 122006 576212 122012 576224
rect 65300 576184 122012 576212
rect 65300 576172 65306 576184
rect 122006 576172 122012 576184
rect 122064 576172 122070 576224
rect 180610 576172 180616 576224
rect 180668 576212 180674 576224
rect 300854 576212 300860 576224
rect 180668 576184 300860 576212
rect 180668 576172 180674 576184
rect 300854 576172 300860 576184
rect 300912 576172 300918 576224
rect 3418 576104 3424 576156
rect 3476 576144 3482 576156
rect 323854 576144 323860 576156
rect 3476 576116 323860 576144
rect 3476 576104 3482 576116
rect 323854 576104 323860 576116
rect 323912 576104 323918 576156
rect 128262 574948 128268 575000
rect 128320 574988 128326 575000
rect 211798 574988 211804 575000
rect 128320 574960 211804 574988
rect 128320 574948 128326 574960
rect 211798 574948 211804 574960
rect 211856 574948 211862 575000
rect 266538 574948 266544 575000
rect 266596 574988 266602 575000
rect 322290 574988 322296 575000
rect 266596 574960 322296 574988
rect 266596 574948 266602 574960
rect 322290 574948 322296 574960
rect 322348 574948 322354 575000
rect 58618 574880 58624 574932
rect 58676 574920 58682 574932
rect 91002 574920 91008 574932
rect 58676 574892 91008 574920
rect 58676 574880 58682 574892
rect 91002 574880 91008 574892
rect 91060 574880 91066 574932
rect 187786 574880 187792 574932
rect 187844 574920 187850 574932
rect 302326 574920 302332 574932
rect 187844 574892 302332 574920
rect 187844 574880 187850 574892
rect 302326 574880 302332 574892
rect 302384 574880 302390 574932
rect 70302 574812 70308 574864
rect 70360 574852 70366 574864
rect 122190 574852 122196 574864
rect 70360 574824 122196 574852
rect 70360 574812 70366 574824
rect 122190 574812 122196 574824
rect 122248 574812 122254 574864
rect 181346 574812 181352 574864
rect 181404 574852 181410 574864
rect 301314 574852 301320 574864
rect 181404 574824 301320 574852
rect 181404 574812 181410 574824
rect 301314 574812 301320 574824
rect 301372 574812 301378 574864
rect 4798 574744 4804 574796
rect 4856 574784 4862 574796
rect 321830 574784 321836 574796
rect 4856 574756 321836 574784
rect 4856 574744 4862 574756
rect 321830 574744 321836 574756
rect 321888 574744 321894 574796
rect 204254 573520 204260 573572
rect 204312 573560 204318 573572
rect 239674 573560 239680 573572
rect 204312 573532 239680 573560
rect 204312 573520 204318 573532
rect 239674 573520 239680 573532
rect 239732 573520 239738 573572
rect 59078 573452 59084 573504
rect 59136 573492 59142 573504
rect 92474 573492 92480 573504
rect 59136 573464 92480 573492
rect 59136 573452 59142 573464
rect 92474 573452 92480 573464
rect 92532 573452 92538 573504
rect 177022 573452 177028 573504
rect 177080 573492 177086 573504
rect 217410 573492 217416 573504
rect 177080 573464 217416 573492
rect 177080 573452 177086 573464
rect 217410 573452 217416 573464
rect 217468 573452 217474 573504
rect 240778 573452 240784 573504
rect 240836 573492 240842 573504
rect 320910 573492 320916 573504
rect 240836 573464 320916 573492
rect 240836 573452 240842 573464
rect 320910 573452 320916 573464
rect 320968 573452 320974 573504
rect 59446 573384 59452 573436
rect 59504 573424 59510 573436
rect 76006 573424 76012 573436
rect 59504 573396 76012 573424
rect 59504 573384 59510 573396
rect 76006 573384 76012 573396
rect 76064 573384 76070 573436
rect 80330 573384 80336 573436
rect 80388 573424 80394 573436
rect 120810 573424 120816 573436
rect 80388 573396 120816 573424
rect 80388 573384 80394 573396
rect 120810 573384 120816 573396
rect 120868 573384 120874 573436
rect 126146 573384 126152 573436
rect 126204 573424 126210 573436
rect 211338 573424 211344 573436
rect 126204 573396 211344 573424
rect 126204 573384 126210 573396
rect 211338 573384 211344 573396
rect 211396 573384 211402 573436
rect 216398 573384 216404 573436
rect 216456 573424 216462 573436
rect 301498 573424 301504 573436
rect 216456 573396 301504 573424
rect 216456 573384 216462 573396
rect 301498 573384 301504 573396
rect 301556 573384 301562 573436
rect 64506 573316 64512 573368
rect 64564 573356 64570 573368
rect 122926 573356 122932 573368
rect 64564 573328 122932 573356
rect 64564 573316 64570 573328
rect 122926 573316 122932 573328
rect 122984 573316 122990 573368
rect 181990 573316 181996 573368
rect 182048 573356 182054 573368
rect 301130 573356 301136 573368
rect 182048 573328 301136 573356
rect 182048 573316 182054 573328
rect 301130 573316 301136 573328
rect 301188 573316 301194 573368
rect 68094 572228 68100 572280
rect 68152 572268 68158 572280
rect 121822 572268 121828 572280
rect 68152 572240 121828 572268
rect 68152 572228 68158 572240
rect 121822 572228 121828 572240
rect 121880 572228 121886 572280
rect 189902 572228 189908 572280
rect 189960 572268 189966 572280
rect 239582 572268 239588 572280
rect 189960 572240 239588 572268
rect 189960 572228 189966 572240
rect 239582 572228 239588 572240
rect 239640 572228 239646 572280
rect 139026 572160 139032 572212
rect 139084 572200 139090 572212
rect 213086 572200 213092 572212
rect 139084 572172 213092 572200
rect 139084 572160 139090 572172
rect 213086 572160 213092 572172
rect 213144 572160 213150 572212
rect 121822 572092 121828 572144
rect 121880 572132 121886 572144
rect 211890 572132 211896 572144
rect 121880 572104 211896 572132
rect 121880 572092 121886 572104
rect 211890 572092 211896 572104
rect 211948 572092 211954 572144
rect 267274 572092 267280 572144
rect 267332 572132 267338 572144
rect 313918 572132 313924 572144
rect 267332 572104 313924 572132
rect 267332 572092 267338 572104
rect 313918 572092 313924 572104
rect 313976 572092 313982 572144
rect 70946 572024 70952 572076
rect 71004 572064 71010 572076
rect 121914 572064 121920 572076
rect 71004 572036 121920 572064
rect 71004 572024 71010 572036
rect 121914 572024 121920 572036
rect 121972 572024 121978 572076
rect 209774 572024 209780 572076
rect 209832 572064 209838 572076
rect 301222 572064 301228 572076
rect 209832 572036 301228 572064
rect 209832 572024 209838 572036
rect 301222 572024 301228 572036
rect 301280 572024 301286 572076
rect 65978 571956 65984 572008
rect 66036 571996 66042 572008
rect 123202 571996 123208 572008
rect 66036 571968 123208 571996
rect 66036 571956 66042 571968
rect 123202 571956 123208 571968
rect 123260 571956 123266 572008
rect 147030 571956 147036 572008
rect 147088 571996 147094 572008
rect 169110 571996 169116 572008
rect 147088 571968 169116 571996
rect 147088 571956 147094 571968
rect 169110 571956 169116 571968
rect 169168 571956 169174 572008
rect 194962 571956 194968 572008
rect 195020 571996 195026 572008
rect 302878 571996 302884 572008
rect 195020 571968 302884 571996
rect 195020 571956 195026 571968
rect 302878 571956 302884 571968
rect 302936 571956 302942 572008
rect 268010 571344 268016 571396
rect 268068 571384 268074 571396
rect 321554 571384 321560 571396
rect 268068 571356 321560 571384
rect 268068 571344 268074 571356
rect 321554 571344 321560 571356
rect 321612 571344 321618 571396
rect 192110 570800 192116 570852
rect 192168 570840 192174 570852
rect 238938 570840 238944 570852
rect 192168 570812 238944 570840
rect 192168 570800 192174 570812
rect 238938 570800 238944 570812
rect 238996 570800 239002 570852
rect 269482 570800 269488 570852
rect 269540 570840 269546 570852
rect 317138 570840 317144 570852
rect 269540 570812 317144 570840
rect 269540 570800 269546 570812
rect 317138 570800 317144 570812
rect 317196 570800 317202 570852
rect 136910 570732 136916 570784
rect 136968 570772 136974 570784
rect 213178 570772 213184 570784
rect 136968 570744 213184 570772
rect 136968 570732 136974 570744
rect 213178 570732 213184 570744
rect 213236 570732 213242 570784
rect 253658 570732 253664 570784
rect 253716 570772 253722 570784
rect 323762 570772 323768 570784
rect 253716 570744 323768 570772
rect 253716 570732 253722 570744
rect 323762 570732 323768 570744
rect 323820 570732 323826 570784
rect 57514 570664 57520 570716
rect 57572 570704 57578 570716
rect 87598 570704 87604 570716
rect 57572 570676 87604 570704
rect 57572 570664 57578 570676
rect 87598 570664 87604 570676
rect 87656 570664 87662 570716
rect 89622 570664 89628 570716
rect 89680 570704 89686 570716
rect 104894 570704 104900 570716
rect 89680 570676 104900 570704
rect 89680 570664 89686 570676
rect 104894 570664 104900 570676
rect 104952 570664 104958 570716
rect 119706 570664 119712 570716
rect 119764 570704 119770 570716
rect 154666 570704 154672 570716
rect 119764 570676 154672 570704
rect 119764 570664 119770 570676
rect 154666 570664 154672 570676
rect 154724 570664 154730 570716
rect 197078 570664 197084 570716
rect 197136 570704 197142 570716
rect 302694 570704 302700 570716
rect 197136 570676 302700 570704
rect 197136 570664 197142 570676
rect 302694 570664 302700 570676
rect 302752 570664 302758 570716
rect 78858 570596 78864 570648
rect 78916 570636 78922 570648
rect 123478 570636 123484 570648
rect 78916 570608 123484 570636
rect 78916 570596 78922 570608
rect 123478 570596 123484 570608
rect 123536 570596 123542 570648
rect 185578 570596 185584 570648
rect 185636 570636 185642 570648
rect 293954 570636 293960 570648
rect 185636 570608 293960 570636
rect 185636 570596 185642 570608
rect 293954 570596 293960 570608
rect 294012 570596 294018 570648
rect 81434 569304 81440 569356
rect 81492 569344 81498 569356
rect 90358 569344 90364 569356
rect 81492 569316 90364 569344
rect 81492 569304 81498 569316
rect 90358 569304 90364 569316
rect 90416 569304 90422 569356
rect 98638 569304 98644 569356
rect 98696 569344 98702 569356
rect 123386 569344 123392 569356
rect 98696 569316 123392 569344
rect 98696 569304 98702 569316
rect 123386 569304 123392 569316
rect 123444 569304 123450 569356
rect 204990 569304 204996 569356
rect 205048 569344 205054 569356
rect 239490 569344 239496 569356
rect 205048 569316 239496 569344
rect 205048 569304 205054 569316
rect 239490 569304 239496 569316
rect 239548 569304 239554 569356
rect 274450 569304 274456 569356
rect 274508 569344 274514 569356
rect 322198 569344 322204 569356
rect 274508 569316 322204 569344
rect 274508 569304 274514 569316
rect 322198 569304 322204 569316
rect 322256 569304 322262 569356
rect 80974 569236 80980 569288
rect 81032 569276 81038 569288
rect 121086 569276 121092 569288
rect 81032 569248 121092 569276
rect 81032 569236 81038 569248
rect 121086 569236 121092 569248
rect 121144 569236 121150 569288
rect 178494 569236 178500 569288
rect 178552 569276 178558 569288
rect 216030 569276 216036 569288
rect 178552 569248 216036 569276
rect 178552 569236 178558 569248
rect 216030 569236 216036 569248
rect 216088 569236 216094 569288
rect 250806 569236 250812 569288
rect 250864 569276 250870 569288
rect 323670 569276 323676 569288
rect 250864 569248 323676 569276
rect 250864 569236 250870 569248
rect 323670 569236 323676 569248
rect 323728 569236 323734 569288
rect 57146 569168 57152 569220
rect 57204 569208 57210 569220
rect 103238 569208 103244 569220
rect 57204 569180 103244 569208
rect 57204 569168 57210 569180
rect 103238 569168 103244 569180
rect 103296 569168 103302 569220
rect 124030 569168 124036 569220
rect 124088 569208 124094 569220
rect 211522 569208 211528 569220
rect 124088 569180 211528 569208
rect 124088 569168 124094 569180
rect 211522 569168 211528 569180
rect 211580 569168 211586 569220
rect 229278 569168 229284 569220
rect 229336 569208 229342 569220
rect 303062 569208 303068 569220
rect 229336 569180 303068 569208
rect 229336 569168 229342 569180
rect 303062 569168 303068 569180
rect 303120 569168 303126 569220
rect 199194 567944 199200 567996
rect 199252 567984 199258 567996
rect 232590 567984 232596 567996
rect 199252 567956 232596 567984
rect 199252 567944 199258 567956
rect 232590 567944 232596 567956
rect 232648 567944 232654 567996
rect 263686 567944 263692 567996
rect 263744 567984 263750 567996
rect 311158 567984 311164 567996
rect 263744 567956 311164 567984
rect 263744 567944 263750 567956
rect 311158 567944 311164 567956
rect 311216 567944 311222 567996
rect 78674 567876 78680 567928
rect 78732 567916 78738 567928
rect 115382 567916 115388 567928
rect 78732 567888 115388 567916
rect 78732 567876 78738 567888
rect 115382 567876 115388 567888
rect 115440 567876 115446 567928
rect 147030 567876 147036 567928
rect 147088 567916 147094 567928
rect 212810 567916 212816 567928
rect 147088 567888 212816 567916
rect 147088 567876 147094 567888
rect 212810 567876 212816 567888
rect 212868 567876 212874 567928
rect 247954 567876 247960 567928
rect 248012 567916 248018 567928
rect 324866 567916 324872 567928
rect 248012 567888 324872 567916
rect 248012 567876 248018 567888
rect 324866 567876 324872 567888
rect 324924 567876 324930 567928
rect 57054 567808 57060 567860
rect 57112 567848 57118 567860
rect 101030 567848 101036 567860
rect 57112 567820 101036 567848
rect 57112 567808 57118 567820
rect 101030 567808 101036 567820
rect 101088 567808 101094 567860
rect 205634 567808 205640 567860
rect 205692 567848 205698 567860
rect 285858 567848 285864 567860
rect 205692 567820 285864 567848
rect 205692 567808 205698 567820
rect 285858 567808 285864 567820
rect 285916 567808 285922 567860
rect 3418 567196 3424 567248
rect 3476 567236 3482 567248
rect 321554 567236 321560 567248
rect 3476 567208 321560 567236
rect 3476 567196 3482 567208
rect 321554 567196 321560 567208
rect 321612 567196 321618 567248
rect 177758 566652 177764 566704
rect 177816 566692 177822 566704
rect 244274 566692 244280 566704
rect 177816 566664 244280 566692
rect 177816 566652 177822 566664
rect 244274 566652 244280 566664
rect 244332 566652 244338 566704
rect 259454 566652 259460 566704
rect 259512 566692 259518 566704
rect 312538 566692 312544 566704
rect 259512 566664 312544 566692
rect 259512 566652 259518 566664
rect 312538 566652 312544 566664
rect 312596 566652 312602 566704
rect 128998 566584 129004 566636
rect 129056 566624 129062 566636
rect 211430 566624 211436 566636
rect 129056 566596 211436 566624
rect 129056 566584 129062 566596
rect 211430 566584 211436 566596
rect 211488 566584 211494 566636
rect 250070 566584 250076 566636
rect 250128 566624 250134 566636
rect 314194 566624 314200 566636
rect 250128 566596 314200 566624
rect 250128 566584 250134 566596
rect 314194 566584 314200 566596
rect 314252 566584 314258 566636
rect 86034 566516 86040 566568
rect 86092 566556 86098 566568
rect 121546 566556 121552 566568
rect 86092 566528 121552 566556
rect 86092 566516 86098 566528
rect 121546 566516 121552 566528
rect 121604 566516 121610 566568
rect 151170 566516 151176 566568
rect 151228 566556 151234 566568
rect 163406 566556 163412 566568
rect 151228 566528 163412 566556
rect 151228 566516 151234 566528
rect 163406 566516 163412 566528
rect 163464 566516 163470 566568
rect 191374 566516 191380 566568
rect 191432 566556 191438 566568
rect 277394 566556 277400 566568
rect 191432 566528 277400 566556
rect 191432 566516 191438 566528
rect 277394 566516 277400 566528
rect 277452 566516 277458 566568
rect 279510 566516 279516 566568
rect 279568 566556 279574 566568
rect 307110 566556 307116 566568
rect 279568 566528 307116 566556
rect 279568 566516 279574 566528
rect 307110 566516 307116 566528
rect 307168 566516 307174 566568
rect 58986 566448 58992 566500
rect 59044 566488 59050 566500
rect 102502 566488 102508 566500
rect 59044 566460 102508 566488
rect 59044 566448 59050 566460
rect 102502 566448 102508 566460
rect 102560 566448 102566 566500
rect 160094 566448 160100 566500
rect 160152 566488 160158 566500
rect 172698 566488 172704 566500
rect 160152 566460 172704 566488
rect 160152 566448 160158 566460
rect 172698 566448 172704 566460
rect 172756 566448 172762 566500
rect 198550 566448 198556 566500
rect 198608 566488 198614 566500
rect 289078 566488 289084 566500
rect 198608 566460 289084 566488
rect 198608 566448 198614 566460
rect 289078 566448 289084 566460
rect 289136 566448 289142 566500
rect 202782 565292 202788 565344
rect 202840 565332 202846 565344
rect 256694 565332 256700 565344
rect 202840 565304 256700 565332
rect 202840 565292 202846 565304
rect 256694 565292 256700 565304
rect 256752 565292 256758 565344
rect 152642 565224 152648 565276
rect 152700 565264 152706 565276
rect 212902 565264 212908 565276
rect 152700 565236 212908 565264
rect 152700 565224 152706 565236
rect 212902 565224 212908 565236
rect 212960 565224 212966 565276
rect 275186 565224 275192 565276
rect 275244 565264 275250 565276
rect 316770 565264 316776 565276
rect 275244 565236 316776 565264
rect 275244 565224 275250 565236
rect 316770 565224 316776 565236
rect 316828 565224 316834 565276
rect 124674 565156 124680 565208
rect 124732 565196 124738 565208
rect 210878 565196 210884 565208
rect 124732 565168 210884 565196
rect 124732 565156 124738 565168
rect 210878 565156 210884 565168
rect 210936 565156 210942 565208
rect 246482 565156 246488 565208
rect 246540 565196 246546 565208
rect 305730 565196 305736 565208
rect 246540 565168 305736 565196
rect 246540 565156 246546 565168
rect 305730 565156 305736 565168
rect 305788 565156 305794 565208
rect 71130 565088 71136 565140
rect 71188 565128 71194 565140
rect 105354 565128 105360 565140
rect 71188 565100 105360 565128
rect 71188 565088 71194 565100
rect 105354 565088 105360 565100
rect 105412 565088 105418 565140
rect 149054 565088 149060 565140
rect 149112 565128 149118 565140
rect 161290 565128 161296 565140
rect 149112 565100 161296 565128
rect 149112 565088 149118 565100
rect 161290 565088 161296 565100
rect 161348 565088 161354 565140
rect 179138 565088 179144 565140
rect 179196 565128 179202 565140
rect 291194 565128 291200 565140
rect 179196 565100 291200 565128
rect 179196 565088 179202 565100
rect 291194 565088 291200 565100
rect 291252 565088 291258 565140
rect 193490 563864 193496 563916
rect 193548 563904 193554 563916
rect 235258 563904 235264 563916
rect 193548 563876 235264 563904
rect 193548 563864 193554 563876
rect 235258 563864 235264 563876
rect 235316 563864 235322 563916
rect 245102 563864 245108 563916
rect 245160 563904 245166 563916
rect 318150 563904 318156 563916
rect 245160 563876 318156 563904
rect 245160 563864 245166 563876
rect 318150 563864 318156 563876
rect 318208 563864 318214 563916
rect 82446 563796 82452 563848
rect 82504 563836 82510 563848
rect 116670 563836 116676 563848
rect 82504 563808 116676 563836
rect 82504 563796 82510 563808
rect 116670 563796 116676 563808
rect 116728 563796 116734 563848
rect 142614 563796 142620 563848
rect 142672 563836 142678 563848
rect 211614 563836 211620 563848
rect 142672 563808 211620 563836
rect 142672 563796 142678 563808
rect 211614 563796 211620 563808
rect 211672 563796 211678 563848
rect 242894 563796 242900 563848
rect 242952 563836 242958 563848
rect 320818 563836 320824 563848
rect 242952 563808 320824 563836
rect 242952 563796 242958 563808
rect 320818 563796 320824 563808
rect 320876 563796 320882 563848
rect 62206 563728 62212 563780
rect 62264 563768 62270 563780
rect 109678 563768 109684 563780
rect 62264 563740 109684 563768
rect 62264 563728 62270 563740
rect 109678 563728 109684 563740
rect 109736 563728 109742 563780
rect 131206 563728 131212 563780
rect 131264 563768 131270 563780
rect 192478 563768 192484 563780
rect 131264 563740 192484 563768
rect 131264 563728 131270 563740
rect 192478 563728 192484 563740
rect 192536 563728 192542 563780
rect 192754 563728 192760 563780
rect 192812 563768 192818 563780
rect 280798 563768 280804 563780
rect 192812 563740 280804 563768
rect 192812 563728 192818 563740
rect 280798 563728 280804 563740
rect 280856 563728 280862 563780
rect 71682 563660 71688 563712
rect 71740 563700 71746 563712
rect 121730 563700 121736 563712
rect 71740 563672 121736 563700
rect 71740 563660 71746 563672
rect 121730 563660 121736 563672
rect 121788 563660 121794 563712
rect 187050 563660 187056 563712
rect 187108 563700 187114 563712
rect 302418 563700 302424 563712
rect 187108 563672 302424 563700
rect 187108 563660 187114 563672
rect 302418 563660 302424 563672
rect 302476 563660 302482 563712
rect 40034 562980 40040 563032
rect 40092 563020 40098 563032
rect 321554 563020 321560 563032
rect 40092 562992 321560 563020
rect 40092 562980 40098 562992
rect 321554 562980 321560 562992
rect 321612 562980 321618 563032
rect 207106 562436 207112 562488
rect 207164 562476 207170 562488
rect 229738 562476 229744 562488
rect 207164 562448 229744 562476
rect 207164 562436 207170 562448
rect 229738 562436 229744 562448
rect 229796 562436 229802 562488
rect 88334 562368 88340 562420
rect 88392 562408 88398 562420
rect 104618 562408 104624 562420
rect 88392 562380 104624 562408
rect 88392 562368 88398 562380
rect 104618 562368 104624 562380
rect 104676 562368 104682 562420
rect 158346 562368 158352 562420
rect 158404 562408 158410 562420
rect 213270 562408 213276 562420
rect 158404 562380 213276 562408
rect 158404 562368 158410 562380
rect 213270 562368 213276 562380
rect 213328 562368 213334 562420
rect 57790 562300 57796 562352
rect 57848 562340 57854 562352
rect 116670 562340 116676 562352
rect 57848 562312 116676 562340
rect 57848 562300 57854 562312
rect 116670 562300 116676 562312
rect 116728 562300 116734 562352
rect 147306 562300 147312 562352
rect 147364 562340 147370 562352
rect 174906 562340 174912 562352
rect 147364 562312 174912 562340
rect 147364 562300 147370 562312
rect 174906 562300 174912 562312
rect 174964 562300 174970 562352
rect 189166 562300 189172 562352
rect 189224 562340 189230 562352
rect 282178 562340 282184 562352
rect 189224 562312 282184 562340
rect 189224 562300 189230 562312
rect 282178 562300 282184 562312
rect 282236 562300 282242 562352
rect 169846 562164 169852 562216
rect 169904 562204 169910 562216
rect 170030 562204 170036 562216
rect 169904 562176 170036 562204
rect 169904 562164 169910 562176
rect 170030 562164 170036 562176
rect 170088 562164 170094 562216
rect 121086 561076 121092 561128
rect 121144 561116 121150 561128
rect 199470 561116 199476 561128
rect 121144 561088 199476 561116
rect 121144 561076 121150 561088
rect 199470 561076 199476 561088
rect 199528 561076 199534 561128
rect 206370 561076 206376 561128
rect 206428 561116 206434 561128
rect 262214 561116 262220 561128
rect 206428 561088 262220 561116
rect 206428 561076 206434 561088
rect 262214 561076 262220 561088
rect 262272 561076 262278 561128
rect 76742 561008 76748 561060
rect 76800 561048 76806 561060
rect 116578 561048 116584 561060
rect 76800 561020 116584 561048
rect 76800 561008 76806 561020
rect 116578 561008 116584 561020
rect 116636 561008 116642 561060
rect 129734 561008 129740 561060
rect 129792 561048 129798 561060
rect 212534 561048 212540 561060
rect 129792 561020 212540 561048
rect 129792 561008 129798 561020
rect 212534 561008 212540 561020
rect 212592 561008 212598 561060
rect 251542 561008 251548 561060
rect 251600 561048 251606 561060
rect 323578 561048 323584 561060
rect 251600 561020 323584 561048
rect 251600 561008 251606 561020
rect 323578 561008 323584 561020
rect 323636 561008 323642 561060
rect 63126 560940 63132 560992
rect 63184 560980 63190 560992
rect 110506 560980 110512 560992
rect 63184 560952 110512 560980
rect 63184 560940 63190 560952
rect 110506 560940 110512 560952
rect 110564 560940 110570 560992
rect 182726 560940 182732 560992
rect 182784 560980 182790 560992
rect 300670 560980 300676 560992
rect 182784 560952 300676 560980
rect 182784 560940 182790 560952
rect 300670 560940 300676 560952
rect 300728 560940 300734 560992
rect 217870 559716 217876 559768
rect 217928 559756 217934 559768
rect 273898 559756 273904 559768
rect 217928 559728 273904 559756
rect 217928 559716 217934 559728
rect 273898 559716 273904 559728
rect 273956 559716 273962 559768
rect 73246 559648 73252 559700
rect 73304 559688 73310 559700
rect 106918 559688 106924 559700
rect 73304 559660 106924 559688
rect 73304 559648 73310 559660
rect 106918 559648 106924 559660
rect 106976 559648 106982 559700
rect 197814 559648 197820 559700
rect 197872 559688 197878 559700
rect 217502 559688 217508 559700
rect 197872 559660 217508 559688
rect 197872 559648 197878 559660
rect 217502 559648 217508 559660
rect 217560 559648 217566 559700
rect 256510 559648 256516 559700
rect 256568 559688 256574 559700
rect 316678 559688 316684 559700
rect 256568 559660 316684 559688
rect 256568 559648 256574 559660
rect 316678 559648 316684 559660
rect 316736 559648 316742 559700
rect 69566 559580 69572 559632
rect 69624 559620 69630 559632
rect 114554 559620 114560 559632
rect 69624 559592 114560 559620
rect 69624 559580 69630 559592
rect 114554 559580 114560 559592
rect 114612 559580 114618 559632
rect 120442 559580 120448 559632
rect 120500 559620 120506 559632
rect 144270 559620 144276 559632
rect 120500 559592 144276 559620
rect 120500 559580 120506 559592
rect 144270 559580 144276 559592
rect 144328 559580 144334 559632
rect 148686 559580 148692 559632
rect 148744 559620 148750 559632
rect 160554 559620 160560 559632
rect 148744 559592 160560 559620
rect 148744 559580 148750 559592
rect 160554 559580 160560 559592
rect 160612 559580 160618 559632
rect 184934 559580 184940 559632
rect 184992 559620 184998 559632
rect 235350 559620 235356 559632
rect 184992 559592 235356 559620
rect 184992 559580 184998 559592
rect 235350 559580 235356 559592
rect 235408 559580 235414 559632
rect 260098 559580 260104 559632
rect 260156 559620 260162 559632
rect 321094 559620 321100 559632
rect 260156 559592 321100 559620
rect 260156 559580 260162 559592
rect 321094 559580 321100 559592
rect 321152 559580 321158 559632
rect 58710 559512 58716 559564
rect 58768 559552 58774 559564
rect 111058 559552 111064 559564
rect 58768 559524 111064 559552
rect 58768 559512 58774 559524
rect 111058 559512 111064 559524
rect 111116 559512 111122 559564
rect 140498 559512 140504 559564
rect 140556 559552 140562 559564
rect 197998 559552 198004 559564
rect 140556 559524 198004 559552
rect 140556 559512 140562 559524
rect 197998 559512 198004 559524
rect 198056 559512 198062 559564
rect 202138 559512 202144 559564
rect 202196 559552 202202 559564
rect 302234 559552 302240 559564
rect 202196 559524 302240 559552
rect 202196 559512 202202 559524
rect 302234 559512 302240 559524
rect 302292 559512 302298 559564
rect 148502 558832 148508 558884
rect 148560 558872 148566 558884
rect 149790 558872 149796 558884
rect 148560 558844 149796 558872
rect 148560 558832 148566 558844
rect 149790 558832 149796 558844
rect 149848 558832 149854 558884
rect 208578 558356 208584 558408
rect 208636 558396 208642 558408
rect 238202 558396 238208 558408
rect 208636 558368 238208 558396
rect 208636 558356 208642 558368
rect 238202 558356 238208 558368
rect 238260 558356 238266 558408
rect 148318 558288 148324 558340
rect 148376 558328 148382 558340
rect 172514 558328 172520 558340
rect 148376 558300 172520 558328
rect 148376 558288 148382 558300
rect 172514 558288 172520 558300
rect 172572 558288 172578 558340
rect 190638 558288 190644 558340
rect 190696 558328 190702 558340
rect 238294 558328 238300 558340
rect 190696 558300 238300 558328
rect 190696 558288 190702 558300
rect 238294 558288 238300 558300
rect 238352 558288 238358 558340
rect 283742 558288 283748 558340
rect 283800 558328 283806 558340
rect 312630 558328 312636 558340
rect 283800 558300 312636 558328
rect 283800 558288 283806 558300
rect 312630 558288 312636 558300
rect 312688 558288 312694 558340
rect 147398 558220 147404 558272
rect 147456 558260 147462 558272
rect 169754 558260 169760 558272
rect 147456 558232 169760 558260
rect 147456 558220 147462 558232
rect 169754 558220 169760 558232
rect 169812 558220 169818 558272
rect 171318 558220 171324 558272
rect 171376 558260 171382 558272
rect 210786 558260 210792 558272
rect 171376 558232 210792 558260
rect 171376 558220 171382 558232
rect 210786 558220 210792 558232
rect 210844 558220 210850 558272
rect 212810 558220 212816 558272
rect 212868 558260 212874 558272
rect 269758 558260 269764 558272
rect 212868 558232 269764 558260
rect 212868 558220 212874 558232
rect 269758 558220 269764 558232
rect 269816 558220 269822 558272
rect 271598 558220 271604 558272
rect 271656 558260 271662 558272
rect 309870 558260 309876 558272
rect 271656 558232 309876 558260
rect 271656 558220 271662 558232
rect 309870 558220 309876 558232
rect 309928 558220 309934 558272
rect 58526 558152 58532 558204
rect 58584 558192 58590 558204
rect 108206 558192 108212 558204
rect 58584 558164 108212 558192
rect 58584 558152 58590 558164
rect 108206 558152 108212 558164
rect 108264 558152 108270 558204
rect 131850 558152 131856 558204
rect 131908 558192 131914 558204
rect 142798 558192 142804 558204
rect 131908 558164 142804 558192
rect 131908 558152 131914 558164
rect 142798 558152 142804 558164
rect 142856 558152 142862 558204
rect 144730 558152 144736 558204
rect 144788 558192 144794 558204
rect 165706 558192 165712 558204
rect 144788 558164 165712 558192
rect 144788 558152 144794 558164
rect 165706 558152 165712 558164
rect 165764 558152 165770 558204
rect 168374 558152 168380 558204
rect 168432 558192 168438 558204
rect 210694 558192 210700 558204
rect 168432 558164 210700 558192
rect 168432 558152 168438 558164
rect 210694 558152 210700 558164
rect 210752 558152 210758 558204
rect 212166 558152 212172 558204
rect 212224 558192 212230 558204
rect 302510 558192 302516 558204
rect 212224 558164 302516 558192
rect 212224 558152 212230 558164
rect 302510 558152 302516 558164
rect 302568 558152 302574 558204
rect 287330 557880 287336 557932
rect 287388 557920 287394 557932
rect 316770 557920 316776 557932
rect 287388 557892 316776 557920
rect 287388 557880 287394 557892
rect 316770 557880 316776 557892
rect 316828 557880 316834 557932
rect 283098 557812 283104 557864
rect 283156 557852 283162 557864
rect 319438 557852 319444 557864
rect 283156 557824 319444 557852
rect 283156 557812 283162 557824
rect 319438 557812 319444 557824
rect 319496 557812 319502 557864
rect 284938 557744 284944 557796
rect 284996 557784 285002 557796
rect 322198 557784 322204 557796
rect 284996 557756 322204 557784
rect 284996 557744 285002 557756
rect 322198 557744 322204 557756
rect 322256 557744 322262 557796
rect 252278 557676 252284 557728
rect 252336 557716 252342 557728
rect 321554 557716 321560 557728
rect 252336 557688 321560 557716
rect 252336 557676 252342 557688
rect 321554 557676 321560 557688
rect 321612 557676 321618 557728
rect 248690 557608 248696 557660
rect 248748 557648 248754 557660
rect 319714 557648 319720 557660
rect 248748 557620 319720 557648
rect 248748 557608 248754 557620
rect 319714 557608 319720 557620
rect 319772 557608 319778 557660
rect 237926 557540 237932 557592
rect 237984 557580 237990 557592
rect 322290 557580 322296 557592
rect 237984 557552 322296 557580
rect 237984 557540 237990 557552
rect 322290 557540 322296 557552
rect 322348 557540 322354 557592
rect 146938 557132 146944 557184
rect 146996 557172 147002 557184
rect 148410 557172 148416 557184
rect 146996 557144 148416 557172
rect 146996 557132 147002 557144
rect 148410 557132 148416 557144
rect 148468 557132 148474 557184
rect 147674 556996 147680 557048
rect 147732 557036 147738 557048
rect 191098 557036 191104 557048
rect 147732 557008 191104 557036
rect 147732 556996 147738 557008
rect 191098 556996 191104 557008
rect 191156 556996 191162 557048
rect 211430 556996 211436 557048
rect 211488 557036 211494 557048
rect 220262 557036 220268 557048
rect 211488 557008 220268 557036
rect 211488 556996 211494 557008
rect 220262 556996 220268 557008
rect 220320 556996 220326 557048
rect 176286 556928 176292 556980
rect 176344 556968 176350 556980
rect 222930 556968 222936 556980
rect 176344 556940 222936 556968
rect 176344 556928 176350 556940
rect 222930 556928 222936 556940
rect 222988 556928 222994 556980
rect 188522 556860 188528 556912
rect 188580 556900 188586 556912
rect 253934 556900 253940 556912
rect 188580 556872 253940 556900
rect 188580 556860 188586 556872
rect 253934 556860 253940 556872
rect 253992 556860 253998 556912
rect 282362 556860 282368 556912
rect 282420 556900 282426 556912
rect 308398 556900 308404 556912
rect 282420 556872 308404 556900
rect 282420 556860 282426 556872
rect 308398 556860 308404 556872
rect 308456 556860 308462 556912
rect 94590 556792 94596 556844
rect 94648 556832 94654 556844
rect 123018 556832 123024 556844
rect 94648 556804 123024 556832
rect 94648 556792 94654 556804
rect 123018 556792 123024 556804
rect 123076 556792 123082 556844
rect 127618 556792 127624 556844
rect 127676 556832 127682 556844
rect 202230 556832 202236 556844
rect 127676 556804 202236 556832
rect 127676 556792 127682 556804
rect 202230 556792 202236 556804
rect 202288 556792 202294 556844
rect 207842 556792 207848 556844
rect 207900 556832 207906 556844
rect 233878 556832 233884 556844
rect 207900 556804 233884 556832
rect 207900 556792 207906 556804
rect 233878 556792 233884 556804
rect 233936 556792 233942 556844
rect 270126 556792 270132 556844
rect 270184 556832 270190 556844
rect 311250 556832 311256 556844
rect 270184 556804 311256 556832
rect 270184 556792 270190 556804
rect 311250 556792 311256 556804
rect 311308 556792 311314 556844
rect 291654 556656 291660 556708
rect 291712 556696 291718 556708
rect 316862 556696 316868 556708
rect 291712 556668 316868 556696
rect 291712 556656 291718 556668
rect 316862 556656 316868 556668
rect 316920 556656 316926 556708
rect 285214 556588 285220 556640
rect 285272 556628 285278 556640
rect 316678 556628 316684 556640
rect 285272 556600 316684 556628
rect 285272 556588 285278 556600
rect 316678 556588 316684 556600
rect 316736 556588 316742 556640
rect 255866 556520 255872 556572
rect 255924 556560 255930 556572
rect 304350 556560 304356 556572
rect 255924 556532 304356 556560
rect 255924 556520 255930 556532
rect 304350 556520 304356 556532
rect 304408 556520 304414 556572
rect 273714 556452 273720 556504
rect 273772 556492 273778 556504
rect 323670 556492 323676 556504
rect 273772 556464 323676 556492
rect 273772 556452 273778 556464
rect 323670 556452 323676 556464
rect 323728 556452 323734 556504
rect 264422 556384 264428 556436
rect 264480 556424 264486 556436
rect 320818 556424 320824 556436
rect 264480 556396 320824 556424
rect 264480 556384 264486 556396
rect 320818 556384 320824 556396
rect 320876 556384 320882 556436
rect 265894 556316 265900 556368
rect 265952 556356 265958 556368
rect 324866 556356 324872 556368
rect 265952 556328 324872 556356
rect 265952 556316 265958 556328
rect 324866 556316 324872 556328
rect 324924 556316 324930 556368
rect 263042 556248 263048 556300
rect 263100 556288 263106 556300
rect 323578 556288 323584 556300
rect 263100 556260 323584 556288
rect 263100 556248 263106 556260
rect 323578 556248 323584 556260
rect 323636 556248 323642 556300
rect 135438 556180 135444 556232
rect 135496 556220 135502 556232
rect 140038 556220 140044 556232
rect 135496 556192 140044 556220
rect 135496 556180 135502 556192
rect 140038 556180 140044 556192
rect 140096 556180 140102 556232
rect 148226 556180 148232 556232
rect 148284 556220 148290 556232
rect 149054 556220 149060 556232
rect 148284 556192 149060 556220
rect 148284 556180 148290 556192
rect 149054 556180 149060 556192
rect 149112 556180 149118 556232
rect 254394 556180 254400 556232
rect 254452 556220 254458 556232
rect 318150 556220 318156 556232
rect 254452 556192 318156 556220
rect 254452 556180 254458 556192
rect 318150 556180 318156 556192
rect 318208 556180 318214 556232
rect 136174 556112 136180 556164
rect 136232 556152 136238 556164
rect 144178 556152 144184 556164
rect 136232 556124 144184 556152
rect 136232 556112 136238 556124
rect 144178 556112 144184 556124
rect 144236 556112 144242 556164
rect 169938 556112 169944 556164
rect 169996 556152 170002 556164
rect 173434 556152 173440 556164
rect 169996 556124 173440 556152
rect 169996 556112 170002 556124
rect 173434 556112 173440 556124
rect 173492 556112 173498 556164
rect 54938 556044 54944 556096
rect 54996 556084 55002 556096
rect 67358 556084 67364 556096
rect 54996 556056 67364 556084
rect 54996 556044 55002 556056
rect 67358 556044 67364 556056
rect 67416 556044 67422 556096
rect 71038 556044 71044 556096
rect 71096 556084 71102 556096
rect 77386 556084 77392 556096
rect 71096 556056 77392 556084
rect 71096 556044 71102 556056
rect 77386 556044 77392 556056
rect 77444 556044 77450 556096
rect 108390 556044 108396 556096
rect 108448 556084 108454 556096
rect 114646 556084 114652 556096
rect 108448 556056 114652 556084
rect 108448 556044 108454 556056
rect 114646 556044 114652 556056
rect 114704 556044 114710 556096
rect 151078 556044 151084 556096
rect 151136 556084 151142 556096
rect 153378 556084 153384 556096
rect 151136 556056 153384 556084
rect 151136 556044 151142 556056
rect 153378 556044 153384 556056
rect 153436 556044 153442 556096
rect 55030 555976 55036 556028
rect 55088 556016 55094 556028
rect 79594 556016 79600 556028
rect 55088 555988 79600 556016
rect 55088 555976 55094 555988
rect 79594 555976 79600 555988
rect 79652 555976 79658 556028
rect 54846 555908 54852 555960
rect 54904 555948 54910 555960
rect 88886 555948 88892 555960
rect 54904 555920 88892 555948
rect 54904 555908 54910 555920
rect 88886 555908 88892 555920
rect 88944 555908 88950 555960
rect 203518 555908 203524 555960
rect 203576 555948 203582 555960
rect 217318 555948 217324 555960
rect 203576 555920 217324 555948
rect 203576 555908 203582 555920
rect 217318 555908 217324 555920
rect 217376 555908 217382 555960
rect 60366 555840 60372 555892
rect 60424 555880 60430 555892
rect 95326 555880 95332 555892
rect 60424 555852 95332 555880
rect 60424 555840 60430 555852
rect 95326 555840 95332 555852
rect 95384 555840 95390 555892
rect 118234 555840 118240 555892
rect 118292 555880 118298 555892
rect 126238 555880 126244 555892
rect 118292 555852 126244 555880
rect 118292 555840 118298 555852
rect 126238 555840 126244 555852
rect 126296 555840 126302 555892
rect 201402 555840 201408 555892
rect 201460 555880 201466 555892
rect 215938 555880 215944 555892
rect 201460 555852 215944 555880
rect 201460 555840 201466 555852
rect 215938 555840 215944 555852
rect 215996 555840 216002 555892
rect 225782 555840 225788 555892
rect 225840 555880 225846 555892
rect 235442 555880 235448 555892
rect 225840 555852 235448 555880
rect 225840 555840 225846 555852
rect 235442 555840 235448 555852
rect 235500 555840 235506 555892
rect 56410 555772 56416 555824
rect 56468 555812 56474 555824
rect 83918 555812 83924 555824
rect 56468 555784 83924 555812
rect 56468 555772 56474 555784
rect 83918 555772 83924 555784
rect 83976 555772 83982 555824
rect 85298 555772 85304 555824
rect 85356 555812 85362 555824
rect 120902 555812 120908 555824
rect 85356 555784 120908 555812
rect 85356 555772 85362 555784
rect 120902 555772 120908 555784
rect 120960 555772 120966 555824
rect 157334 555772 157340 555824
rect 157392 555812 157398 555824
rect 166994 555812 167000 555824
rect 157392 555784 167000 555812
rect 157392 555772 157398 555784
rect 166994 555772 167000 555784
rect 167052 555772 167058 555824
rect 186314 555772 186320 555824
rect 186372 555812 186378 555824
rect 206278 555812 206284 555824
rect 186372 555784 206284 555812
rect 186372 555772 186378 555784
rect 206278 555772 206284 555784
rect 206336 555772 206342 555824
rect 209222 555772 209228 555824
rect 209280 555812 209286 555824
rect 220170 555812 220176 555824
rect 209280 555784 220176 555812
rect 209280 555772 209286 555784
rect 220170 555772 220176 555784
rect 220228 555772 220234 555824
rect 221458 555772 221464 555824
rect 221516 555812 221522 555824
rect 231302 555812 231308 555824
rect 221516 555784 231308 555812
rect 221516 555772 221522 555784
rect 231302 555772 231308 555784
rect 231360 555772 231366 555824
rect 55122 555704 55128 555756
rect 55180 555744 55186 555756
rect 93210 555744 93216 555756
rect 55180 555716 93216 555744
rect 55180 555704 55186 555716
rect 93210 555704 93216 555716
rect 93268 555704 93274 555756
rect 114002 555704 114008 555756
rect 114060 555744 114066 555756
rect 122834 555744 122840 555756
rect 114060 555716 122840 555744
rect 114060 555704 114066 555716
rect 122834 555704 122840 555716
rect 122892 555704 122898 555756
rect 146110 555704 146116 555756
rect 146168 555744 146174 555756
rect 156966 555744 156972 555756
rect 146168 555716 156972 555744
rect 146168 555704 146174 555716
rect 156966 555704 156972 555716
rect 157024 555704 157030 555756
rect 199930 555704 199936 555756
rect 199988 555744 199994 555756
rect 220078 555744 220084 555756
rect 199988 555716 220084 555744
rect 199988 555704 199994 555716
rect 220078 555704 220084 555716
rect 220136 555704 220142 555756
rect 230750 555704 230756 555756
rect 230808 555744 230814 555756
rect 244918 555744 244924 555756
rect 230808 555716 244924 555744
rect 230808 555704 230814 555716
rect 244918 555704 244924 555716
rect 244976 555704 244982 555756
rect 278038 555704 278044 555756
rect 278096 555744 278102 555756
rect 300302 555744 300308 555756
rect 278096 555716 300308 555744
rect 278096 555704 278102 555716
rect 300302 555704 300308 555716
rect 300360 555704 300366 555756
rect 59262 555636 59268 555688
rect 59320 555676 59326 555688
rect 99650 555676 99656 555688
rect 59320 555648 99656 555676
rect 59320 555636 59326 555648
rect 99650 555636 99656 555648
rect 99708 555636 99714 555688
rect 106826 555636 106832 555688
rect 106884 555676 106890 555688
rect 124306 555676 124312 555688
rect 106884 555648 124312 555676
rect 106884 555636 106890 555648
rect 124306 555636 124312 555648
rect 124364 555636 124370 555688
rect 147490 555636 147496 555688
rect 147548 555676 147554 555688
rect 157702 555676 157708 555688
rect 147548 555648 157708 555676
rect 147548 555636 147554 555648
rect 157702 555636 157708 555648
rect 157760 555636 157766 555688
rect 169754 555636 169760 555688
rect 169812 555676 169818 555688
rect 175550 555676 175556 555688
rect 169812 555648 175556 555676
rect 169812 555636 169818 555648
rect 175550 555636 175556 555648
rect 175608 555636 175614 555688
rect 194226 555636 194232 555688
rect 194284 555676 194290 555688
rect 214558 555676 214564 555688
rect 194284 555648 214564 555676
rect 194284 555636 194290 555648
rect 214558 555636 214564 555648
rect 214616 555636 214622 555688
rect 225046 555636 225052 555688
rect 225104 555676 225110 555688
rect 242158 555676 242164 555688
rect 225104 555648 242164 555676
rect 225104 555636 225110 555648
rect 242158 555636 242164 555648
rect 242216 555636 242222 555688
rect 270862 555636 270868 555688
rect 270920 555676 270926 555688
rect 324682 555676 324688 555688
rect 270920 555648 324688 555676
rect 270920 555636 270926 555648
rect 324682 555636 324688 555648
rect 324740 555636 324746 555688
rect 56502 555568 56508 555620
rect 56560 555608 56566 555620
rect 98914 555608 98920 555620
rect 56560 555580 98920 555608
rect 56560 555568 56566 555580
rect 98914 555568 98920 555580
rect 98972 555568 98978 555620
rect 103974 555568 103980 555620
rect 104032 555608 104038 555620
rect 124214 555608 124220 555620
rect 104032 555580 124220 555608
rect 104032 555568 104038 555580
rect 124214 555568 124220 555580
rect 124272 555568 124278 555620
rect 151998 555568 152004 555620
rect 152056 555608 152062 555620
rect 167730 555608 167736 555620
rect 152056 555580 167736 555608
rect 152056 555568 152062 555580
rect 167730 555568 167736 555580
rect 167788 555568 167794 555620
rect 170582 555568 170588 555620
rect 170640 555608 170646 555620
rect 199378 555608 199384 555620
rect 170640 555580 199384 555608
rect 170640 555568 170646 555580
rect 199378 555568 199384 555580
rect 199436 555568 199442 555620
rect 209958 555568 209964 555620
rect 210016 555608 210022 555620
rect 231210 555608 231216 555620
rect 210016 555580 231216 555608
rect 210016 555568 210022 555580
rect 231210 555568 231216 555580
rect 231268 555568 231274 555620
rect 231486 555568 231492 555620
rect 231544 555608 231550 555620
rect 249058 555608 249064 555620
rect 231544 555580 249064 555608
rect 231544 555568 231550 555580
rect 249058 555568 249064 555580
rect 249116 555568 249122 555620
rect 252922 555568 252928 555620
rect 252980 555608 252986 555620
rect 323762 555608 323768 555620
rect 252980 555580 323768 555608
rect 252980 555568 252986 555580
rect 323762 555568 323768 555580
rect 323820 555568 323826 555620
rect 61654 555500 61660 555552
rect 61712 555540 61718 555552
rect 64138 555540 64144 555552
rect 61712 555512 64144 555540
rect 61712 555500 61718 555512
rect 64138 555500 64144 555512
rect 64196 555500 64202 555552
rect 73798 555540 73804 555552
rect 64340 555512 73804 555540
rect 56318 555364 56324 555416
rect 56376 555404 56382 555416
rect 64340 555404 64368 555512
rect 73798 555500 73804 555512
rect 73856 555500 73862 555552
rect 78122 555500 78128 555552
rect 78180 555540 78186 555552
rect 121454 555540 121460 555552
rect 78180 555512 121460 555540
rect 78180 555500 78186 555512
rect 121454 555500 121460 555512
rect 121512 555500 121518 555552
rect 138290 555500 138296 555552
rect 138348 555540 138354 555552
rect 147030 555540 147036 555552
rect 138348 555512 147036 555540
rect 138348 555500 138354 555512
rect 147030 555500 147036 555512
rect 147088 555500 147094 555552
rect 147582 555500 147588 555552
rect 147640 555540 147646 555552
rect 171962 555540 171968 555552
rect 147640 555512 171968 555540
rect 147640 555500 147646 555512
rect 171962 555500 171968 555512
rect 172020 555500 172026 555552
rect 195606 555500 195612 555552
rect 195664 555540 195670 555552
rect 238110 555540 238116 555552
rect 195664 555512 238116 555540
rect 195664 555500 195670 555512
rect 238110 555500 238116 555512
rect 238168 555500 238174 555552
rect 261570 555500 261576 555552
rect 261628 555540 261634 555552
rect 286318 555540 286324 555552
rect 261628 555512 286324 555540
rect 261628 555500 261634 555512
rect 286318 555500 286324 555512
rect 286376 555500 286382 555552
rect 298646 555500 298652 555552
rect 298704 555540 298710 555552
rect 302050 555540 302056 555552
rect 298704 555512 302056 555540
rect 298704 555500 298710 555512
rect 302050 555500 302056 555512
rect 302108 555500 302114 555552
rect 116854 555472 116860 555484
rect 56376 555376 64368 555404
rect 64846 555444 116860 555472
rect 56376 555364 56382 555376
rect 61378 555296 61384 555348
rect 61436 555336 61442 555348
rect 64846 555336 64874 555444
rect 116854 555432 116860 555444
rect 116912 555432 116918 555484
rect 118970 555432 118976 555484
rect 119028 555472 119034 555484
rect 129090 555472 129096 555484
rect 119028 555444 129096 555472
rect 119028 555432 119034 555444
rect 129090 555432 129096 555444
rect 129148 555432 129154 555484
rect 144086 555432 144092 555484
rect 144144 555472 144150 555484
rect 195238 555472 195244 555484
rect 144144 555444 195244 555472
rect 144144 555432 144150 555444
rect 195238 555432 195244 555444
rect 195296 555432 195302 555484
rect 213546 555432 213552 555484
rect 213604 555472 213610 555484
rect 236638 555472 236644 555484
rect 213604 555444 236644 555472
rect 213604 555432 213610 555444
rect 236638 555432 236644 555444
rect 236696 555432 236702 555484
rect 237190 555432 237196 555484
rect 237248 555472 237254 555484
rect 284938 555472 284944 555484
rect 237248 555444 284944 555472
rect 237248 555432 237254 555444
rect 284938 555432 284944 555444
rect 284996 555432 285002 555484
rect 299566 555432 299572 555484
rect 299624 555472 299630 555484
rect 318058 555472 318064 555484
rect 299624 555444 318064 555472
rect 299624 555432 299630 555444
rect 318058 555432 318064 555444
rect 318116 555432 318122 555484
rect 72418 555364 72424 555416
rect 72476 555404 72482 555416
rect 73154 555404 73160 555416
rect 72476 555376 73160 555404
rect 72476 555364 72482 555376
rect 73154 555364 73160 555376
rect 73212 555364 73218 555416
rect 113266 555364 113272 555416
rect 113324 555404 113330 555416
rect 119338 555404 119344 555416
rect 113324 555376 119344 555404
rect 113324 555364 113330 555376
rect 119338 555364 119344 555376
rect 119396 555364 119402 555416
rect 242250 555364 242256 555416
rect 242308 555404 242314 555416
rect 324130 555404 324136 555416
rect 242308 555376 324136 555404
rect 242308 555364 242314 555376
rect 324130 555364 324136 555376
rect 324188 555364 324194 555416
rect 61436 555308 64874 555336
rect 61436 555296 61442 555308
rect 276566 555296 276572 555348
rect 276624 555336 276630 555348
rect 300394 555336 300400 555348
rect 276624 555308 300400 555336
rect 276624 555296 276630 555308
rect 300394 555296 300400 555308
rect 300452 555296 300458 555348
rect 79318 555228 79324 555280
rect 79376 555268 79382 555280
rect 81710 555268 81716 555280
rect 79376 555240 81716 555268
rect 79376 555228 79382 555240
rect 81710 555228 81716 555240
rect 81768 555228 81774 555280
rect 87598 555228 87604 555280
rect 87656 555268 87662 555280
rect 91738 555268 91744 555280
rect 87656 555240 91744 555268
rect 87656 555228 87662 555240
rect 91738 555228 91744 555240
rect 91796 555228 91802 555280
rect 96062 555228 96068 555280
rect 96120 555268 96126 555280
rect 98638 555268 98644 555280
rect 96120 555240 98644 555268
rect 96120 555228 96126 555240
rect 98638 555228 98644 555240
rect 98696 555228 98702 555280
rect 104158 555228 104164 555280
rect 104216 555268 104222 555280
rect 106090 555268 106096 555280
rect 104216 555240 106096 555268
rect 104216 555228 104222 555240
rect 106090 555228 106096 555240
rect 106148 555228 106154 555280
rect 108298 555228 108304 555280
rect 108356 555268 108362 555280
rect 111794 555268 111800 555280
rect 108356 555240 111800 555268
rect 108356 555228 108362 555240
rect 111794 555228 111800 555240
rect 111852 555228 111858 555280
rect 115198 555228 115204 555280
rect 115256 555268 115262 555280
rect 116118 555268 116124 555280
rect 115256 555240 116124 555268
rect 115256 555228 115262 555240
rect 116118 555228 116124 555240
rect 116176 555228 116182 555280
rect 116670 555228 116676 555280
rect 116728 555268 116734 555280
rect 117590 555268 117596 555280
rect 116728 555240 117596 555268
rect 116728 555228 116734 555240
rect 117590 555228 117596 555240
rect 117648 555228 117654 555280
rect 144914 555228 144920 555280
rect 144972 555268 144978 555280
rect 146202 555268 146208 555280
rect 144972 555240 146208 555268
rect 144972 555228 144978 555240
rect 146202 555228 146208 555240
rect 146260 555228 146266 555280
rect 149882 555228 149888 555280
rect 149940 555268 149946 555280
rect 151262 555268 151268 555280
rect 149940 555240 151268 555268
rect 149940 555228 149946 555240
rect 151262 555228 151268 555240
rect 151320 555228 151326 555280
rect 154114 555228 154120 555280
rect 154172 555268 154178 555280
rect 160738 555268 160744 555280
rect 154172 555240 160744 555268
rect 154172 555228 154178 555240
rect 160738 555228 160744 555240
rect 160796 555228 160802 555280
rect 219986 555228 219992 555280
rect 220044 555268 220050 555280
rect 228358 555268 228364 555280
rect 220044 555240 228364 555268
rect 220044 555228 220050 555240
rect 228358 555228 228364 555240
rect 228416 555228 228422 555280
rect 230014 555228 230020 555280
rect 230072 555268 230078 555280
rect 231118 555268 231124 555280
rect 230072 555240 231124 555268
rect 230072 555228 230078 555240
rect 231118 555228 231124 555240
rect 231176 555228 231182 555280
rect 277302 555228 277308 555280
rect 277360 555268 277366 555280
rect 277360 555240 298784 555268
rect 277360 555228 277366 555240
rect 105538 555160 105544 555212
rect 105596 555200 105602 555212
rect 108942 555200 108948 555212
rect 105596 555172 108948 555200
rect 105596 555160 105602 555172
rect 108942 555160 108948 555172
rect 109000 555160 109006 555212
rect 275922 555160 275928 555212
rect 275980 555200 275986 555212
rect 298646 555200 298652 555212
rect 275980 555172 298652 555200
rect 275980 555160 275986 555172
rect 298646 555160 298652 555172
rect 298704 555160 298710 555212
rect 298756 555200 298784 555240
rect 298830 555228 298836 555280
rect 298888 555268 298894 555280
rect 304258 555268 304264 555280
rect 298888 555240 304264 555268
rect 298888 555228 298894 555240
rect 304258 555228 304264 555240
rect 304316 555228 304322 555280
rect 301866 555200 301872 555212
rect 298756 555172 301872 555200
rect 301866 555160 301872 555172
rect 301924 555160 301930 555212
rect 290918 555092 290924 555144
rect 290976 555132 290982 555144
rect 322474 555132 322480 555144
rect 290976 555104 322480 555132
rect 290976 555092 290982 555104
rect 322474 555092 322480 555104
rect 322532 555092 322538 555144
rect 280154 555024 280160 555076
rect 280212 555064 280218 555076
rect 322658 555064 322664 555076
rect 280212 555036 322664 555064
rect 280212 555024 280218 555036
rect 322658 555024 322664 555036
rect 322716 555024 322722 555076
rect 257246 554956 257252 555008
rect 257304 554996 257310 555008
rect 300486 554996 300492 555008
rect 257304 554968 300492 554996
rect 257304 554956 257310 554968
rect 300486 554956 300492 554968
rect 300544 554956 300550 555008
rect 265158 554888 265164 554940
rect 265216 554928 265222 554940
rect 274634 554928 274640 554940
rect 265216 554900 274640 554928
rect 265216 554888 265222 554900
rect 274634 554888 274640 554900
rect 274692 554888 274698 554940
rect 301498 554928 301504 554940
rect 296686 554900 301504 554928
rect 281626 554820 281632 554872
rect 281684 554860 281690 554872
rect 296686 554860 296714 554900
rect 301498 554888 301504 554900
rect 301556 554888 301562 554940
rect 301590 554860 301596 554872
rect 281684 554832 296714 554860
rect 296748 554832 301596 554860
rect 281684 554820 281690 554832
rect 295978 554752 295984 554804
rect 296036 554792 296042 554804
rect 296748 554792 296776 554832
rect 301590 554820 301596 554832
rect 301648 554820 301654 554872
rect 296036 554764 296776 554792
rect 296036 554752 296042 554764
rect 296806 554752 296812 554804
rect 296864 554792 296870 554804
rect 300118 554792 300124 554804
rect 296864 554764 300124 554792
rect 296864 554752 296870 554764
rect 300118 554752 300124 554764
rect 300176 554752 300182 554804
rect 240042 554276 240048 554328
rect 240100 554316 240106 554328
rect 303062 554316 303068 554328
rect 240100 554288 303068 554316
rect 240100 554276 240106 554288
rect 303062 554276 303068 554288
rect 303120 554276 303126 554328
rect 236454 554208 236460 554260
rect 236512 554248 236518 554260
rect 321646 554248 321652 554260
rect 236512 554220 321652 554248
rect 236512 554208 236518 554220
rect 321646 554208 321652 554220
rect 321704 554208 321710 554260
rect 235810 554140 235816 554192
rect 235868 554180 235874 554192
rect 324038 554180 324044 554192
rect 235868 554152 324044 554180
rect 235868 554140 235874 554152
rect 324038 554140 324044 554152
rect 324096 554140 324102 554192
rect 268746 554072 268752 554124
rect 268804 554112 268810 554124
rect 302970 554112 302976 554124
rect 268804 554084 302976 554112
rect 268804 554072 268810 554084
rect 302970 554072 302976 554084
rect 303028 554072 303034 554124
rect 274634 554004 274640 554056
rect 274692 554044 274698 554056
rect 324314 554044 324320 554056
rect 274692 554016 324320 554044
rect 274692 554004 274698 554016
rect 324314 554004 324320 554016
rect 324372 554004 324378 554056
rect 260834 553936 260840 553988
rect 260892 553976 260898 553988
rect 305638 553976 305644 553988
rect 260892 553948 305644 553976
rect 260892 553936 260898 553948
rect 305638 553936 305644 553948
rect 305696 553936 305702 553988
rect 272334 553868 272340 553920
rect 272392 553908 272398 553920
rect 324590 553908 324596 553920
rect 272392 553880 324596 553908
rect 272392 553868 272398 553880
rect 324590 553868 324596 553880
rect 324648 553868 324654 553920
rect 247218 553800 247224 553852
rect 247276 553840 247282 553852
rect 301774 553840 301780 553852
rect 247276 553812 301780 553840
rect 247276 553800 247282 553812
rect 301774 553800 301780 553812
rect 301832 553800 301838 553852
rect 243630 553732 243636 553784
rect 243688 553772 243694 553784
rect 300670 553772 300676 553784
rect 243688 553744 300676 553772
rect 243688 553732 243694 553744
rect 300670 553732 300676 553744
rect 300728 553732 300734 553784
rect 262306 553664 262312 553716
rect 262364 553704 262370 553716
rect 324774 553704 324780 553716
rect 262364 553676 324780 553704
rect 262364 553664 262370 553676
rect 324774 553664 324780 553676
rect 324832 553664 324838 553716
rect 284478 553596 284484 553648
rect 284536 553636 284542 553648
rect 319530 553636 319536 553648
rect 284536 553608 319536 553636
rect 284536 553596 284542 553608
rect 319530 553596 319536 553608
rect 319588 553596 319594 553648
rect 244366 553528 244372 553580
rect 244424 553568 244430 553580
rect 322566 553568 322572 553580
rect 244424 553540 322572 553568
rect 244424 553528 244430 553540
rect 322566 553528 322572 553540
rect 322624 553528 322630 553580
rect 278774 553460 278780 553512
rect 278832 553500 278838 553512
rect 299382 553500 299388 553512
rect 278832 553472 299388 553500
rect 278832 553460 278838 553472
rect 299382 553460 299388 553472
rect 299440 553460 299446 553512
rect 273070 553392 273076 553444
rect 273128 553432 273134 553444
rect 301682 553432 301688 553444
rect 273128 553404 301688 553432
rect 273128 553392 273134 553404
rect 301682 553392 301688 553404
rect 301740 553392 301746 553444
rect 299382 553324 299388 553376
rect 299440 553364 299446 553376
rect 321554 553364 321560 553376
rect 299440 553336 321560 553364
rect 299440 553324 299446 553336
rect 321554 553324 321560 553336
rect 321612 553324 321618 553376
rect 3510 553052 3516 553104
rect 3568 553092 3574 553104
rect 322750 553092 322756 553104
rect 3568 553064 322756 553092
rect 3568 553052 3574 553064
rect 322750 553052 322756 553064
rect 322808 553052 322814 553104
rect 302234 545096 302240 545148
rect 302292 545136 302298 545148
rect 304258 545136 304264 545148
rect 302292 545108 304264 545136
rect 302292 545096 302298 545108
rect 304258 545096 304264 545108
rect 304316 545096 304322 545148
rect 300670 543668 300676 543720
rect 300728 543708 300734 543720
rect 321554 543708 321560 543720
rect 300728 543680 321560 543708
rect 300728 543668 300734 543680
rect 321554 543668 321560 543680
rect 321612 543668 321618 543720
rect 436830 543192 436836 543244
rect 436888 543192 436894 543244
rect 436278 543056 436284 543108
rect 436336 543056 436342 543108
rect 436296 542892 436324 543056
rect 436848 543040 436876 543192
rect 436830 542988 436836 543040
rect 436888 542988 436894 543040
rect 436646 542892 436652 542904
rect 436296 542864 436652 542892
rect 436646 542852 436652 542864
rect 436704 542852 436710 542904
rect 303062 539520 303068 539572
rect 303120 539560 303126 539572
rect 321554 539560 321560 539572
rect 303120 539532 321560 539560
rect 303120 539520 303126 539532
rect 321554 539520 321560 539532
rect 321612 539520 321618 539572
rect 324130 535372 324136 535424
rect 324188 535412 324194 535424
rect 436554 535412 436560 535424
rect 324188 535384 436560 535412
rect 324188 535372 324194 535384
rect 436554 535372 436560 535384
rect 436612 535372 436618 535424
rect 324314 534556 324320 534608
rect 324372 534596 324378 534608
rect 325142 534596 325148 534608
rect 324372 534568 325148 534596
rect 324372 534556 324378 534568
rect 325142 534556 325148 534568
rect 325200 534556 325206 534608
rect 300210 534012 300216 534064
rect 300268 534052 300274 534064
rect 436278 534052 436284 534064
rect 300268 534024 436284 534052
rect 300268 534012 300274 534024
rect 436278 534012 436284 534024
rect 436336 534012 436342 534064
rect 300302 533944 300308 533996
rect 300360 533984 300366 533996
rect 436094 533984 436100 533996
rect 300360 533956 436100 533984
rect 300360 533944 300366 533956
rect 436094 533944 436100 533956
rect 436152 533944 436158 533996
rect 300486 533876 300492 533928
rect 300544 533916 300550 533928
rect 436830 533916 436836 533928
rect 300544 533888 436836 533916
rect 300544 533876 300550 533888
rect 436830 533876 436836 533888
rect 436888 533876 436894 533928
rect 301866 533808 301872 533860
rect 301924 533848 301930 533860
rect 436370 533848 436376 533860
rect 301924 533820 436376 533848
rect 301924 533808 301930 533820
rect 436370 533808 436376 533820
rect 436428 533808 436434 533860
rect 319714 533740 319720 533792
rect 319772 533780 319778 533792
rect 433334 533780 433340 533792
rect 319772 533752 433340 533780
rect 319772 533740 319778 533752
rect 433334 533740 433340 533752
rect 433392 533740 433398 533792
rect 322658 533672 322664 533724
rect 322716 533712 322722 533724
rect 434622 533712 434628 533724
rect 322716 533684 434628 533712
rect 322716 533672 322722 533684
rect 434622 533672 434628 533684
rect 434680 533672 434686 533724
rect 323762 533604 323768 533656
rect 323820 533644 323826 533656
rect 436738 533644 436744 533656
rect 323820 533616 436744 533644
rect 323820 533604 323826 533616
rect 436738 533604 436744 533616
rect 436796 533604 436802 533656
rect 323946 533536 323952 533588
rect 324004 533576 324010 533588
rect 436922 533576 436928 533588
rect 324004 533548 436928 533576
rect 324004 533536 324010 533548
rect 436922 533536 436928 533548
rect 436980 533536 436986 533588
rect 324682 533468 324688 533520
rect 324740 533508 324746 533520
rect 436646 533508 436652 533520
rect 324740 533480 436652 533508
rect 324740 533468 324746 533480
rect 436646 533468 436652 533480
rect 436704 533468 436710 533520
rect 322290 533400 322296 533452
rect 322348 533440 322354 533452
rect 433794 533440 433800 533452
rect 322348 533412 433800 533440
rect 322348 533400 322354 533412
rect 433794 533400 433800 533412
rect 433852 533400 433858 533452
rect 302050 532856 302056 532908
rect 302108 532896 302114 532908
rect 356238 532896 356244 532908
rect 302108 532868 356244 532896
rect 302108 532856 302114 532868
rect 356238 532856 356244 532868
rect 356296 532856 356302 532908
rect 307018 532788 307024 532840
rect 307076 532828 307082 532840
rect 374270 532828 374276 532840
rect 307076 532800 374276 532828
rect 307076 532788 307082 532800
rect 374270 532788 374276 532800
rect 374328 532788 374334 532840
rect 300394 532720 300400 532772
rect 300452 532760 300458 532772
rect 419994 532760 420000 532772
rect 300452 532732 420000 532760
rect 300452 532720 300458 532732
rect 419994 532720 420000 532732
rect 420052 532720 420058 532772
rect 324038 532652 324044 532704
rect 324096 532692 324102 532704
rect 338206 532692 338212 532704
rect 324096 532664 338212 532692
rect 324096 532652 324102 532664
rect 338206 532652 338212 532664
rect 338264 532652 338270 532704
rect 322566 532584 322572 532636
rect 322624 532624 322630 532636
rect 424502 532624 424508 532636
rect 322624 532596 424508 532624
rect 322624 532584 322630 532596
rect 424502 532584 424508 532596
rect 424560 532584 424566 532636
rect 324774 532516 324780 532568
rect 324832 532556 324838 532568
rect 334066 532556 334072 532568
rect 324832 532528 334072 532556
rect 324832 532516 324838 532528
rect 334066 532516 334072 532528
rect 334124 532516 334130 532568
rect 302970 532448 302976 532500
rect 303028 532488 303034 532500
rect 393314 532488 393320 532500
rect 303028 532460 393320 532488
rect 303028 532448 303034 532460
rect 393314 532448 393320 532460
rect 393372 532448 393378 532500
rect 323578 532380 323584 532432
rect 323636 532420 323642 532432
rect 406470 532420 406476 532432
rect 323636 532392 406476 532420
rect 323636 532380 323642 532392
rect 406470 532380 406476 532392
rect 406528 532380 406534 532432
rect 323670 532312 323676 532364
rect 323728 532352 323734 532364
rect 401962 532352 401968 532364
rect 323728 532324 401968 532352
rect 323728 532312 323734 532324
rect 401962 532312 401968 532324
rect 402020 532312 402026 532364
rect 301682 532244 301688 532296
rect 301740 532284 301746 532296
rect 369854 532284 369860 532296
rect 301740 532256 369860 532284
rect 301740 532244 301746 532256
rect 369854 532244 369860 532256
rect 369912 532244 369918 532296
rect 324866 532176 324872 532228
rect 324924 532216 324930 532228
rect 388438 532216 388444 532228
rect 324924 532188 388444 532216
rect 324924 532176 324930 532188
rect 388438 532176 388444 532188
rect 388496 532176 388502 532228
rect 301774 532108 301780 532160
rect 301832 532148 301838 532160
rect 365254 532148 365260 532160
rect 301832 532120 365260 532148
rect 301832 532108 301838 532120
rect 365254 532108 365260 532120
rect 365312 532108 365318 532160
rect 320818 532040 320824 532092
rect 320876 532080 320882 532092
rect 379514 532080 379520 532092
rect 320876 532052 379520 532080
rect 320876 532040 320882 532052
rect 379514 532040 379520 532052
rect 379572 532040 379578 532092
rect 318150 531972 318156 532024
rect 318208 532012 318214 532024
rect 351914 532012 351920 532024
rect 318208 531984 351920 532012
rect 318208 531972 318214 531984
rect 351914 531972 351920 531984
rect 351972 531972 351978 532024
rect 305638 531904 305644 531956
rect 305696 531944 305702 531956
rect 347222 531944 347228 531956
rect 305696 531916 347228 531944
rect 305696 531904 305702 531916
rect 347222 531904 347228 531916
rect 347280 531904 347286 531956
rect 304350 531836 304356 531888
rect 304408 531876 304414 531888
rect 411346 531876 411352 531888
rect 304408 531848 411352 531876
rect 304408 531836 304414 531848
rect 411346 531836 411352 531848
rect 411404 531836 411410 531888
rect 324590 531768 324596 531820
rect 324648 531808 324654 531820
rect 415486 531808 415492 531820
rect 324648 531780 415492 531808
rect 324648 531768 324654 531780
rect 415486 531768 415492 531780
rect 415544 531768 415550 531820
rect 302878 531224 302884 531276
rect 302936 531264 302942 531276
rect 495434 531264 495440 531276
rect 302936 531236 495440 531264
rect 302936 531224 302942 531236
rect 495434 531224 495440 531236
rect 495492 531224 495498 531276
rect 322382 531156 322388 531208
rect 322440 531196 322446 531208
rect 512178 531196 512184 531208
rect 322440 531168 512184 531196
rect 322440 531156 322446 531168
rect 512178 531156 512184 531168
rect 512236 531156 512242 531208
rect 322474 531088 322480 531140
rect 322532 531128 322538 531140
rect 488534 531128 488540 531140
rect 322532 531100 488540 531128
rect 322532 531088 322538 531100
rect 488534 531088 488540 531100
rect 488592 531088 488598 531140
rect 300118 531020 300124 531072
rect 300176 531060 300182 531072
rect 459554 531060 459560 531072
rect 300176 531032 459560 531060
rect 300176 531020 300182 531032
rect 459554 531020 459560 531032
rect 459612 531020 459618 531072
rect 316770 530952 316776 531004
rect 316828 530992 316834 531004
rect 476114 530992 476120 531004
rect 316828 530964 476120 530992
rect 316828 530952 316834 530964
rect 476114 530952 476120 530964
rect 476172 530952 476178 531004
rect 301590 530884 301596 530936
rect 301648 530924 301654 530936
rect 457438 530924 457444 530936
rect 301648 530896 457444 530924
rect 301648 530884 301654 530896
rect 457438 530884 457444 530896
rect 457496 530884 457502 530936
rect 316862 530816 316868 530868
rect 316920 530856 316926 530868
rect 457622 530856 457628 530868
rect 316920 530828 457628 530856
rect 316920 530816 316926 530828
rect 457622 530816 457628 530828
rect 457680 530816 457686 530868
rect 301498 530748 301504 530800
rect 301556 530788 301562 530800
rect 436462 530788 436468 530800
rect 301556 530760 436468 530788
rect 301556 530748 301562 530760
rect 436462 530748 436468 530760
rect 436520 530748 436526 530800
rect 302418 529932 302424 529984
rect 302476 529972 302482 529984
rect 520918 529972 520924 529984
rect 302476 529944 520924 529972
rect 302476 529932 302482 529944
rect 520918 529932 520924 529944
rect 520976 529932 520982 529984
rect 316954 529864 316960 529916
rect 317012 529904 317018 529916
rect 512270 529904 512276 529916
rect 317012 529876 512276 529904
rect 317012 529864 317018 529876
rect 512270 529864 512276 529876
rect 512328 529864 512334 529916
rect 319622 529796 319628 529848
rect 319680 529836 319686 529848
rect 500954 529836 500960 529848
rect 319680 529808 500960 529836
rect 319680 529796 319686 529808
rect 500954 529796 500960 529808
rect 501012 529796 501018 529848
rect 316678 529728 316684 529780
rect 316736 529768 316742 529780
rect 470594 529768 470600 529780
rect 316736 529740 470600 529768
rect 316736 529728 316742 529740
rect 470594 529728 470600 529740
rect 470652 529728 470658 529780
rect 319806 529660 319812 529712
rect 319864 529700 319870 529712
rect 465074 529700 465080 529712
rect 319864 529672 465080 529700
rect 319864 529660 319870 529672
rect 465074 529660 465080 529672
rect 465132 529660 465138 529712
rect 319438 529592 319444 529644
rect 319496 529632 319502 529644
rect 433518 529632 433524 529644
rect 319496 529604 433524 529632
rect 319496 529592 319502 529604
rect 433518 529592 433524 529604
rect 433576 529592 433582 529644
rect 319530 529524 319536 529576
rect 319588 529564 319594 529576
rect 433702 529564 433708 529576
rect 319588 529536 433708 529564
rect 319588 529524 319594 529536
rect 433702 529524 433708 529536
rect 433760 529524 433766 529576
rect 322198 529456 322204 529508
rect 322256 529496 322262 529508
rect 433426 529496 433432 529508
rect 322256 529468 433432 529496
rect 322256 529456 322262 529468
rect 433426 529456 433432 529468
rect 433484 529456 433490 529508
rect 329742 529388 329748 529440
rect 329800 529428 329806 529440
rect 434714 529428 434720 529440
rect 329800 529400 434720 529428
rect 329800 529388 329806 529400
rect 434714 529388 434720 529400
rect 434772 529388 434778 529440
rect 363598 527824 363604 527876
rect 363656 527864 363662 527876
rect 506474 527864 506480 527876
rect 363656 527836 506480 527864
rect 363656 527824 363662 527836
rect 506474 527824 506480 527836
rect 506532 527824 506538 527876
rect 53742 521704 53748 521756
rect 53800 521744 53806 521756
rect 57698 521744 57704 521756
rect 53800 521716 57704 521744
rect 53800 521704 53806 521716
rect 57698 521704 57704 521716
rect 57756 521704 57762 521756
rect 302878 499536 302884 499588
rect 302936 499576 302942 499588
rect 518158 499576 518164 499588
rect 302936 499548 518164 499576
rect 302936 499536 302942 499548
rect 518158 499536 518164 499548
rect 518216 499536 518222 499588
rect 304258 494708 304264 494760
rect 304316 494748 304322 494760
rect 580258 494748 580264 494760
rect 304316 494720 580264 494748
rect 304316 494708 304322 494720
rect 580258 494708 580264 494720
rect 580316 494708 580322 494760
rect 49418 492124 49424 492176
rect 49476 492164 49482 492176
rect 82170 492164 82176 492176
rect 49476 492136 82176 492164
rect 49476 492124 49482 492136
rect 82170 492124 82176 492136
rect 82228 492124 82234 492176
rect 50982 492056 50988 492108
rect 51040 492096 51046 492108
rect 84378 492096 84384 492108
rect 51040 492068 84384 492096
rect 51040 492056 51046 492068
rect 84378 492056 84384 492068
rect 84436 492056 84442 492108
rect 140774 492056 140780 492108
rect 140832 492096 140838 492108
rect 198918 492096 198924 492108
rect 140832 492068 198924 492096
rect 140832 492056 140838 492068
rect 198918 492056 198924 492068
rect 198976 492056 198982 492108
rect 51902 491988 51908 492040
rect 51960 492028 51966 492040
rect 99374 492028 99380 492040
rect 51960 492000 99380 492028
rect 51960 491988 51966 492000
rect 99374 491988 99380 492000
rect 99432 491988 99438 492040
rect 109034 491988 109040 492040
rect 109092 492028 109098 492040
rect 197446 492028 197452 492040
rect 109092 492000 197452 492028
rect 109092 491988 109098 492000
rect 197446 491988 197452 492000
rect 197504 491988 197510 492040
rect 15838 491920 15844 491972
rect 15896 491960 15902 491972
rect 383654 491960 383660 491972
rect 15896 491932 383660 491960
rect 15896 491920 15902 491932
rect 383654 491920 383660 491932
rect 383712 491920 383718 491972
rect 214006 491512 214012 491564
rect 214064 491552 214070 491564
rect 214926 491552 214932 491564
rect 214064 491524 214932 491552
rect 214064 491512 214070 491524
rect 214926 491512 214932 491524
rect 214984 491512 214990 491564
rect 59354 491444 59360 491496
rect 59412 491484 59418 491496
rect 60274 491484 60280 491496
rect 59412 491456 60280 491484
rect 59412 491444 59418 491456
rect 60274 491444 60280 491456
rect 60332 491444 60338 491496
rect 204438 491444 204444 491496
rect 204496 491484 204502 491496
rect 204806 491484 204812 491496
rect 204496 491456 204812 491484
rect 204496 491444 204502 491456
rect 204806 491444 204812 491456
rect 204864 491444 204870 491496
rect 207014 491444 207020 491496
rect 207072 491484 207078 491496
rect 207750 491484 207756 491496
rect 207072 491456 207756 491484
rect 207072 491444 207078 491456
rect 207750 491444 207756 491456
rect 207808 491444 207814 491496
rect 209774 491444 209780 491496
rect 209832 491484 209838 491496
rect 210510 491484 210516 491496
rect 209832 491456 210516 491484
rect 209832 491444 209838 491456
rect 210510 491444 210516 491456
rect 210568 491444 210574 491496
rect 213914 491444 213920 491496
rect 213972 491484 213978 491496
rect 214374 491484 214380 491496
rect 213972 491456 214380 491484
rect 213972 491444 213978 491456
rect 214374 491444 214380 491456
rect 214432 491444 214438 491496
rect 215294 491444 215300 491496
rect 215352 491484 215358 491496
rect 216214 491484 216220 491496
rect 215352 491456 216220 491484
rect 215352 491444 215358 491456
rect 216214 491444 216220 491456
rect 216272 491444 216278 491496
rect 219894 491444 219900 491496
rect 219952 491484 219958 491496
rect 220078 491484 220084 491496
rect 219952 491456 220084 491484
rect 219952 491444 219958 491456
rect 220078 491444 220084 491456
rect 220136 491444 220142 491496
rect 64138 491240 64144 491292
rect 64196 491280 64202 491292
rect 86218 491280 86224 491292
rect 64196 491252 86224 491280
rect 64196 491240 64202 491252
rect 86218 491240 86224 491252
rect 86276 491240 86282 491292
rect 153470 491240 153476 491292
rect 153528 491280 153534 491292
rect 212534 491280 212540 491292
rect 153528 491252 212540 491280
rect 153528 491240 153534 491252
rect 212534 491240 212540 491252
rect 212592 491240 212598 491292
rect 213822 491240 213828 491292
rect 213880 491280 213886 491292
rect 219250 491280 219256 491292
rect 213880 491252 219256 491280
rect 213880 491240 213886 491252
rect 219250 491240 219256 491252
rect 219308 491240 219314 491292
rect 68278 491172 68284 491224
rect 68336 491212 68342 491224
rect 95326 491212 95332 491224
rect 68336 491184 95332 491212
rect 68336 491172 68342 491184
rect 95326 491172 95332 491184
rect 95384 491172 95390 491224
rect 150894 491172 150900 491224
rect 150952 491212 150958 491224
rect 150952 491184 201908 491212
rect 150952 491172 150958 491184
rect 62850 491104 62856 491156
rect 62908 491144 62914 491156
rect 91370 491144 91376 491156
rect 62908 491116 91376 491144
rect 62908 491104 62914 491116
rect 91370 491104 91376 491116
rect 91428 491104 91434 491156
rect 152182 491104 152188 491156
rect 152240 491144 152246 491156
rect 152240 491116 201816 491144
rect 152240 491104 152246 491116
rect 72418 491036 72424 491088
rect 72476 491076 72482 491088
rect 103330 491076 103336 491088
rect 72476 491048 103336 491076
rect 72476 491036 72482 491048
rect 103330 491036 103336 491048
rect 103388 491036 103394 491088
rect 149514 491036 149520 491088
rect 149572 491076 149578 491088
rect 201586 491076 201592 491088
rect 149572 491048 201592 491076
rect 149572 491036 149578 491048
rect 201586 491036 201592 491048
rect 201644 491036 201650 491088
rect 50890 490968 50896 491020
rect 50948 491008 50954 491020
rect 68922 491008 68928 491020
rect 50948 490980 68928 491008
rect 50948 490968 50954 490980
rect 68922 490968 68928 490980
rect 68980 490968 68986 491020
rect 72510 490968 72516 491020
rect 72568 491008 72574 491020
rect 104618 491008 104624 491020
rect 72568 490980 104624 491008
rect 72568 490968 72574 490980
rect 104618 490968 104624 490980
rect 104676 490968 104682 491020
rect 157886 490968 157892 491020
rect 157944 491008 157950 491020
rect 201678 491008 201684 491020
rect 157944 490980 201684 491008
rect 157944 490968 157950 490980
rect 201678 490968 201684 490980
rect 201736 490968 201742 491020
rect 52270 490900 52276 490952
rect 52328 490940 52334 490952
rect 84838 490940 84844 490952
rect 52328 490912 84844 490940
rect 52328 490900 52334 490912
rect 84838 490900 84844 490912
rect 84896 490900 84902 490952
rect 149974 490900 149980 490952
rect 150032 490940 150038 490952
rect 200758 490940 200764 490952
rect 150032 490912 200764 490940
rect 150032 490900 150038 490912
rect 200758 490900 200764 490912
rect 200816 490900 200822 490952
rect 201788 490940 201816 491116
rect 201880 491076 201908 491184
rect 201954 491172 201960 491224
rect 202012 491212 202018 491224
rect 206646 491212 206652 491224
rect 202012 491184 206652 491212
rect 202012 491172 202018 491184
rect 206646 491172 206652 491184
rect 206704 491172 206710 491224
rect 211614 491172 211620 491224
rect 211672 491212 211678 491224
rect 218146 491212 218152 491224
rect 211672 491184 218152 491212
rect 211672 491172 211678 491184
rect 218146 491172 218152 491184
rect 218204 491172 218210 491224
rect 289998 491172 290004 491224
rect 290056 491212 290062 491224
rect 356974 491212 356980 491224
rect 290056 491184 356980 491212
rect 290056 491172 290062 491184
rect 356974 491172 356980 491184
rect 357032 491172 357038 491224
rect 248598 491104 248604 491156
rect 248656 491144 248662 491156
rect 361114 491144 361120 491156
rect 248656 491116 361120 491144
rect 248656 491104 248662 491116
rect 361114 491104 361120 491116
rect 361172 491104 361178 491156
rect 205634 491076 205640 491088
rect 201880 491048 205640 491076
rect 205634 491036 205640 491048
rect 205692 491036 205698 491088
rect 240686 491036 240692 491088
rect 240744 491076 240750 491088
rect 356790 491076 356796 491088
rect 240744 491048 356796 491076
rect 240744 491036 240750 491048
rect 356790 491036 356796 491048
rect 356848 491036 356854 491088
rect 239398 490968 239404 491020
rect 239456 491008 239462 491020
rect 356698 491008 356704 491020
rect 239456 490980 356704 491008
rect 239456 490968 239462 490980
rect 356698 490968 356704 490980
rect 356756 490968 356762 491020
rect 204254 490940 204260 490952
rect 201788 490912 204260 490940
rect 204254 490900 204260 490912
rect 204312 490900 204318 490952
rect 238938 490900 238944 490952
rect 238996 490940 239002 490952
rect 358262 490940 358268 490952
rect 238996 490912 358268 490940
rect 238996 490900 239002 490912
rect 358262 490900 358268 490912
rect 358320 490900 358326 490952
rect 53558 490832 53564 490884
rect 53616 490872 53622 490884
rect 86126 490872 86132 490884
rect 53616 490844 86132 490872
rect 53616 490832 53622 490844
rect 86126 490832 86132 490844
rect 86184 490832 86190 490884
rect 156598 490832 156604 490884
rect 156656 490872 156662 490884
rect 205634 490872 205640 490884
rect 156656 490844 205640 490872
rect 156656 490832 156662 490844
rect 205634 490832 205640 490844
rect 205692 490832 205698 490884
rect 207934 490832 207940 490884
rect 207992 490872 207998 490884
rect 217410 490872 217416 490884
rect 207992 490844 217416 490872
rect 207992 490832 207998 490844
rect 217410 490832 217416 490844
rect 217468 490832 217474 490884
rect 237650 490832 237656 490884
rect 237708 490872 237714 490884
rect 365162 490872 365168 490884
rect 237708 490844 365168 490872
rect 237708 490832 237714 490844
rect 365162 490832 365168 490844
rect 365220 490832 365226 490884
rect 59078 490764 59084 490816
rect 59136 490804 59142 490816
rect 91830 490804 91836 490816
rect 59136 490776 91836 490804
rect 59136 490764 59142 490776
rect 91830 490764 91836 490776
rect 91888 490764 91894 490816
rect 155310 490764 155316 490816
rect 155368 490804 155374 490816
rect 209038 490804 209044 490816
rect 155368 490776 209044 490804
rect 155368 490764 155374 490776
rect 209038 490764 209044 490776
rect 209096 490764 209102 490816
rect 233234 490764 233240 490816
rect 233292 490804 233298 490816
rect 363690 490804 363696 490816
rect 233292 490776 363696 490804
rect 233292 490764 233298 490776
rect 363690 490764 363696 490776
rect 363748 490764 363754 490816
rect 55122 490696 55128 490748
rect 55180 490736 55186 490748
rect 89162 490736 89168 490748
rect 55180 490708 89168 490736
rect 55180 490696 55186 490708
rect 89162 490696 89168 490708
rect 89220 490696 89226 490748
rect 139394 490696 139400 490748
rect 139452 490736 139458 490748
rect 193950 490736 193956 490748
rect 139452 490708 193956 490736
rect 139452 490696 139458 490708
rect 193950 490696 193956 490708
rect 194008 490696 194014 490748
rect 194870 490696 194876 490748
rect 194928 490736 194934 490748
rect 196802 490736 196808 490748
rect 194928 490708 196808 490736
rect 194928 490696 194934 490708
rect 196802 490696 196808 490708
rect 196860 490696 196866 490748
rect 206554 490696 206560 490748
rect 206612 490736 206618 490748
rect 217778 490736 217784 490748
rect 206612 490708 217784 490736
rect 206612 490696 206618 490708
rect 217778 490696 217784 490708
rect 217836 490696 217842 490748
rect 225322 490696 225328 490748
rect 225380 490736 225386 490748
rect 358170 490736 358176 490748
rect 225380 490708 358176 490736
rect 225380 490696 225386 490708
rect 358170 490696 358176 490708
rect 358228 490696 358234 490748
rect 49050 490628 49056 490680
rect 49108 490668 49114 490680
rect 97166 490668 97172 490680
rect 49108 490640 97172 490668
rect 49108 490628 49114 490640
rect 97166 490628 97172 490640
rect 97224 490628 97230 490680
rect 138934 490628 138940 490680
rect 138992 490668 138998 490680
rect 193858 490668 193864 490680
rect 138992 490640 193864 490668
rect 138992 490628 138998 490640
rect 193858 490628 193864 490640
rect 193916 490628 193922 490680
rect 195330 490628 195336 490680
rect 195388 490668 195394 490680
rect 199378 490668 199384 490680
rect 195388 490640 199384 490668
rect 195388 490628 195394 490640
rect 199378 490628 199384 490640
rect 199436 490628 199442 490680
rect 201678 490628 201684 490680
rect 201736 490668 201742 490680
rect 208394 490668 208400 490680
rect 201736 490640 208400 490668
rect 201736 490628 201742 490640
rect 208394 490628 208400 490640
rect 208452 490628 208458 490680
rect 209406 490628 209412 490680
rect 209464 490668 209470 490680
rect 210050 490668 210056 490680
rect 209464 490640 210056 490668
rect 209464 490628 209470 490640
rect 210050 490628 210056 490640
rect 210108 490628 210114 490680
rect 223574 490628 223580 490680
rect 223632 490668 223638 490680
rect 360930 490668 360936 490680
rect 223632 490640 360936 490668
rect 223632 490628 223638 490640
rect 360930 490628 360936 490640
rect 360988 490628 360994 490680
rect 41046 490560 41052 490612
rect 41104 490600 41110 490612
rect 100202 490600 100208 490612
rect 41104 490572 100208 490600
rect 41104 490560 41110 490572
rect 100202 490560 100208 490572
rect 100260 490560 100266 490612
rect 110322 490560 110328 490612
rect 110380 490600 110386 490612
rect 180058 490600 180064 490612
rect 110380 490572 180064 490600
rect 110380 490560 110386 490572
rect 180058 490560 180064 490572
rect 180116 490560 180122 490612
rect 200666 490560 200672 490612
rect 200724 490600 200730 490612
rect 217410 490600 217416 490612
rect 200724 490572 217416 490600
rect 200724 490560 200730 490572
rect 217410 490560 217416 490572
rect 217468 490560 217474 490612
rect 223114 490560 223120 490612
rect 223172 490600 223178 490612
rect 374638 490600 374644 490612
rect 223172 490572 374644 490600
rect 223172 490560 223178 490572
rect 374638 490560 374644 490572
rect 374696 490560 374702 490612
rect 58526 490492 58532 490544
rect 58584 490532 58590 490544
rect 81250 490532 81256 490544
rect 58584 490504 81256 490532
rect 58584 490492 58590 490504
rect 81250 490492 81256 490504
rect 81308 490492 81314 490544
rect 157426 490492 157432 490544
rect 157484 490532 157490 490544
rect 204254 490532 204260 490544
rect 157484 490504 204260 490532
rect 157484 490492 157490 490504
rect 204254 490492 204260 490504
rect 204312 490492 204318 490544
rect 53650 490424 53656 490476
rect 53708 490464 53714 490476
rect 74258 490464 74264 490476
rect 53708 490436 74264 490464
rect 53708 490424 53714 490436
rect 74258 490424 74264 490436
rect 74316 490424 74322 490476
rect 154390 490424 154396 490476
rect 154448 490464 154454 490476
rect 200574 490464 200580 490476
rect 154448 490436 200580 490464
rect 154448 490424 154454 490436
rect 200574 490424 200580 490436
rect 200632 490424 200638 490476
rect 204070 490424 204076 490476
rect 204128 490464 204134 490476
rect 219158 490464 219164 490476
rect 204128 490436 219164 490464
rect 204128 490424 204134 490436
rect 219158 490424 219164 490436
rect 219216 490424 219222 490476
rect 56318 490356 56324 490408
rect 56376 490396 56382 490408
rect 71774 490396 71780 490408
rect 56376 490368 71780 490396
rect 56376 490356 56382 490368
rect 71774 490356 71780 490368
rect 71832 490356 71838 490408
rect 153102 490356 153108 490408
rect 153160 490396 153166 490408
rect 197354 490396 197360 490408
rect 153160 490368 197360 490396
rect 153160 490356 153166 490368
rect 197354 490356 197360 490368
rect 197412 490356 197418 490408
rect 68370 490288 68376 490340
rect 68428 490328 68434 490340
rect 85206 490328 85212 490340
rect 68428 490300 85212 490328
rect 68428 490288 68434 490300
rect 85206 490288 85212 490300
rect 85264 490288 85270 490340
rect 203242 490288 203248 490340
rect 203300 490328 203306 490340
rect 212258 490328 212264 490340
rect 203300 490300 212264 490328
rect 203300 490288 203306 490300
rect 212258 490288 212264 490300
rect 212316 490288 212322 490340
rect 67726 489948 67732 490000
rect 67784 489988 67790 490000
rect 68186 489988 68192 490000
rect 67784 489960 68192 489988
rect 67784 489948 67790 489960
rect 68186 489948 68192 489960
rect 68244 489948 68250 490000
rect 218698 489948 218704 490000
rect 218756 489988 218762 490000
rect 219618 489988 219624 490000
rect 218756 489960 219624 489988
rect 218756 489948 218762 489960
rect 219618 489948 219624 489960
rect 219676 489948 219682 490000
rect 50062 489880 50068 489932
rect 50120 489920 50126 489932
rect 72234 489920 72240 489932
rect 50120 489892 72240 489920
rect 50120 489880 50126 489892
rect 72234 489880 72240 489892
rect 72292 489880 72298 489932
rect 208578 489880 208584 489932
rect 208636 489920 208642 489932
rect 211246 489920 211252 489932
rect 208636 489892 211252 489920
rect 208636 489880 208642 489892
rect 211246 489880 211252 489892
rect 211304 489880 211310 489932
rect 283834 489336 283840 489388
rect 283892 489376 283898 489388
rect 359734 489376 359740 489388
rect 283892 489348 359740 489376
rect 283892 489336 283898 489348
rect 359734 489336 359740 489348
rect 359792 489336 359798 489388
rect 257890 489268 257896 489320
rect 257948 489308 257954 489320
rect 373534 489308 373540 489320
rect 257948 489280 373540 489308
rect 257948 489268 257954 489280
rect 373534 489268 373540 489280
rect 373592 489268 373598 489320
rect 167638 489200 167644 489252
rect 167696 489240 167702 489252
rect 210510 489240 210516 489252
rect 167696 489212 210516 489240
rect 167696 489200 167702 489212
rect 210510 489200 210516 489212
rect 210568 489200 210574 489252
rect 242066 489200 242072 489252
rect 242124 489240 242130 489252
rect 361022 489240 361028 489252
rect 242124 489212 361028 489240
rect 242124 489200 242130 489212
rect 361022 489200 361028 489212
rect 361080 489200 361086 489252
rect 59446 489132 59452 489184
rect 59504 489172 59510 489184
rect 160738 489172 160744 489184
rect 59504 489144 160744 489172
rect 59504 489132 59510 489144
rect 160738 489132 160744 489144
rect 160796 489132 160802 489184
rect 164050 489132 164056 489184
rect 164108 489172 164114 489184
rect 215938 489172 215944 489184
rect 164108 489144 215944 489172
rect 164108 489132 164114 489144
rect 215938 489132 215944 489144
rect 215996 489132 216002 489184
rect 222194 489132 222200 489184
rect 222252 489172 222258 489184
rect 376018 489172 376024 489184
rect 222252 489144 376024 489172
rect 222252 489132 222258 489144
rect 376018 489132 376024 489144
rect 376076 489132 376082 489184
rect 47946 488452 47952 488504
rect 48004 488492 48010 488504
rect 97994 488492 98000 488504
rect 48004 488464 98000 488492
rect 48004 488452 48010 488464
rect 97994 488452 98000 488464
rect 98052 488452 98058 488504
rect 59722 488384 59728 488436
rect 59780 488424 59786 488436
rect 119614 488424 119620 488436
rect 59780 488396 119620 488424
rect 59780 488384 59786 488396
rect 119614 488384 119620 488396
rect 119672 488384 119678 488436
rect 48038 488316 48044 488368
rect 48096 488356 48102 488368
rect 111702 488356 111708 488368
rect 48096 488328 111708 488356
rect 48096 488316 48102 488328
rect 111702 488316 111708 488328
rect 111760 488316 111766 488368
rect 46382 488248 46388 488300
rect 46440 488288 46446 488300
rect 111242 488288 111248 488300
rect 46440 488260 111248 488288
rect 46440 488248 46446 488260
rect 111242 488248 111248 488260
rect 111300 488248 111306 488300
rect 160094 488248 160100 488300
rect 160152 488288 160158 488300
rect 209130 488288 209136 488300
rect 160152 488260 209136 488288
rect 160152 488248 160158 488260
rect 209130 488248 209136 488260
rect 209188 488248 209194 488300
rect 50522 488180 50528 488232
rect 50580 488220 50586 488232
rect 116026 488220 116032 488232
rect 50580 488192 116032 488220
rect 50580 488180 50586 488192
rect 116026 488180 116032 488192
rect 116084 488180 116090 488232
rect 138566 488180 138572 488232
rect 138624 488220 138630 488232
rect 196986 488220 196992 488232
rect 138624 488192 196992 488220
rect 138624 488180 138630 488192
rect 196986 488180 196992 488192
rect 197044 488180 197050 488232
rect 46290 488112 46296 488164
rect 46348 488152 46354 488164
rect 112070 488152 112076 488164
rect 46348 488124 112076 488152
rect 46348 488112 46354 488124
rect 112070 488112 112076 488124
rect 112128 488112 112134 488164
rect 137646 488112 137652 488164
rect 137704 488152 137710 488164
rect 197722 488152 197728 488164
rect 137704 488124 197728 488152
rect 137704 488112 137710 488124
rect 197722 488112 197728 488124
rect 197780 488112 197786 488164
rect 48958 488044 48964 488096
rect 49016 488084 49022 488096
rect 115198 488084 115204 488096
rect 49016 488056 115204 488084
rect 49016 488044 49022 488056
rect 115198 488044 115204 488056
rect 115256 488044 115262 488096
rect 136726 488044 136732 488096
rect 136784 488084 136790 488096
rect 197630 488084 197636 488096
rect 136784 488056 197636 488084
rect 136784 488044 136790 488056
rect 197630 488044 197636 488056
rect 197688 488044 197694 488096
rect 46842 487976 46848 488028
rect 46900 488016 46906 488028
rect 115658 488016 115664 488028
rect 46900 487988 115664 488016
rect 46900 487976 46906 487988
rect 115658 487976 115664 487988
rect 115716 487976 115722 488028
rect 136358 487976 136364 488028
rect 136416 488016 136422 488028
rect 198090 488016 198096 488028
rect 136416 487988 198096 488016
rect 136416 487976 136422 487988
rect 198090 487976 198096 487988
rect 198148 487976 198154 488028
rect 59354 487908 59360 487960
rect 59412 487948 59418 487960
rect 133138 487948 133144 487960
rect 59412 487920 133144 487948
rect 59412 487908 59418 487920
rect 133138 487908 133144 487920
rect 133196 487908 133202 487960
rect 138106 487908 138112 487960
rect 138164 487948 138170 487960
rect 200298 487948 200304 487960
rect 138164 487920 200304 487948
rect 138164 487908 138170 487920
rect 200298 487908 200304 487920
rect 200356 487908 200362 487960
rect 256970 487908 256976 487960
rect 257028 487948 257034 487960
rect 367922 487948 367928 487960
rect 257028 487920 367928 487948
rect 257028 487908 257034 487920
rect 367922 487908 367928 487920
rect 367980 487908 367986 487960
rect 56410 487840 56416 487892
rect 56468 487880 56474 487892
rect 131942 487880 131948 487892
rect 56468 487852 131948 487880
rect 56468 487840 56474 487852
rect 131942 487840 131948 487852
rect 132000 487840 132006 487892
rect 135438 487840 135444 487892
rect 135496 487880 135502 487892
rect 198182 487880 198188 487892
rect 135496 487852 198188 487880
rect 135496 487840 135502 487852
rect 198182 487840 198188 487852
rect 198240 487840 198246 487892
rect 246850 487840 246856 487892
rect 246908 487880 246914 487892
rect 363782 487880 363788 487892
rect 246908 487852 363788 487880
rect 246908 487840 246914 487852
rect 363782 487840 363788 487852
rect 363840 487840 363846 487892
rect 48866 487772 48872 487824
rect 48924 487812 48930 487824
rect 134610 487812 134616 487824
rect 48924 487784 134616 487812
rect 48924 487772 48930 487784
rect 134610 487772 134616 487784
rect 134668 487772 134674 487824
rect 144730 487772 144736 487824
rect 144788 487812 144794 487824
rect 218698 487812 218704 487824
rect 144788 487784 218704 487812
rect 144788 487772 144794 487784
rect 218698 487772 218704 487784
rect 218756 487772 218762 487824
rect 236730 487772 236736 487824
rect 236788 487812 236794 487824
rect 370498 487812 370504 487824
rect 236788 487784 370504 487812
rect 236788 487772 236794 487784
rect 370498 487772 370504 487784
rect 370556 487772 370562 487824
rect 50430 487704 50436 487756
rect 50488 487744 50494 487756
rect 97534 487744 97540 487756
rect 50488 487716 97540 487744
rect 50488 487704 50494 487716
rect 97534 487704 97540 487716
rect 97592 487704 97598 487756
rect 51810 487636 51816 487688
rect 51868 487676 51874 487688
rect 98454 487676 98460 487688
rect 51868 487648 98460 487676
rect 51868 487636 51874 487648
rect 98454 487636 98460 487648
rect 98512 487636 98518 487688
rect 54846 487568 54852 487620
rect 54904 487608 54910 487620
rect 96798 487608 96804 487620
rect 54904 487580 96804 487608
rect 54904 487568 54910 487580
rect 96798 487568 96804 487580
rect 96856 487568 96862 487620
rect 177298 486548 177304 486600
rect 177356 486588 177362 486600
rect 203702 486588 203708 486600
rect 177356 486560 203708 486588
rect 177356 486548 177362 486560
rect 203702 486548 203708 486560
rect 203760 486548 203766 486600
rect 260926 486548 260932 486600
rect 260984 486588 260990 486600
rect 366726 486588 366732 486600
rect 260984 486560 366732 486588
rect 260984 486548 260990 486560
rect 366726 486548 366732 486560
rect 366784 486548 366790 486600
rect 164510 486480 164516 486532
rect 164568 486520 164574 486532
rect 211798 486520 211804 486532
rect 164568 486492 211804 486520
rect 164568 486480 164574 486492
rect 211798 486480 211804 486492
rect 211856 486480 211862 486532
rect 242434 486480 242440 486532
rect 242492 486520 242498 486532
rect 363874 486520 363880 486532
rect 242492 486492 363880 486520
rect 242492 486480 242498 486492
rect 363874 486480 363880 486492
rect 363932 486480 363938 486532
rect 144270 486412 144276 486464
rect 144328 486452 144334 486464
rect 213270 486452 213276 486464
rect 144328 486424 213276 486452
rect 144328 486412 144334 486424
rect 213270 486412 213276 486424
rect 213328 486412 213334 486464
rect 247770 486412 247776 486464
rect 247828 486452 247834 486464
rect 374822 486452 374828 486464
rect 247828 486424 374828 486452
rect 247828 486412 247834 486424
rect 374822 486412 374828 486424
rect 374880 486412 374886 486464
rect 57146 485732 57152 485784
rect 57204 485772 57210 485784
rect 132402 485772 132408 485784
rect 57204 485744 132408 485772
rect 57204 485732 57210 485744
rect 132402 485732 132408 485744
rect 132460 485732 132466 485784
rect 58618 485664 58624 485716
rect 58676 485704 58682 485716
rect 132770 485704 132776 485716
rect 58676 485676 132776 485704
rect 58676 485664 58682 485676
rect 132770 485664 132776 485676
rect 132828 485664 132834 485716
rect 44082 485596 44088 485648
rect 44140 485636 44146 485648
rect 119154 485636 119160 485648
rect 44140 485608 119160 485636
rect 44140 485596 44146 485608
rect 119154 485596 119160 485608
rect 119212 485596 119218 485648
rect 54478 485528 54484 485580
rect 54536 485568 54542 485580
rect 129734 485568 129740 485580
rect 54536 485540 129740 485568
rect 54536 485528 54542 485540
rect 129734 485528 129740 485540
rect 129792 485528 129798 485580
rect 57882 485460 57888 485512
rect 57940 485500 57946 485512
rect 135898 485500 135904 485512
rect 57940 485472 135904 485500
rect 57940 485460 57946 485472
rect 135898 485460 135904 485472
rect 135956 485460 135962 485512
rect 47762 485392 47768 485444
rect 47820 485432 47826 485444
rect 129274 485432 129280 485444
rect 47820 485404 129280 485432
rect 47820 485392 47826 485404
rect 129274 485392 129280 485404
rect 129332 485392 129338 485444
rect 47854 485324 47860 485376
rect 47912 485364 47918 485376
rect 131022 485364 131028 485376
rect 47912 485336 131028 485364
rect 47912 485324 47918 485336
rect 131022 485324 131028 485336
rect 131080 485324 131086 485376
rect 50154 485256 50160 485308
rect 50212 485296 50218 485308
rect 131482 485296 131488 485308
rect 50212 485268 131488 485296
rect 50212 485256 50218 485268
rect 131482 485256 131488 485268
rect 131540 485256 131546 485308
rect 44634 485188 44640 485240
rect 44692 485228 44698 485240
rect 130194 485228 130200 485240
rect 44692 485200 130200 485228
rect 44692 485188 44698 485200
rect 130194 485188 130200 485200
rect 130252 485188 130258 485240
rect 284294 485188 284300 485240
rect 284352 485228 284358 485240
rect 359826 485228 359832 485240
rect 284352 485200 359832 485228
rect 284352 485188 284358 485200
rect 359826 485188 359832 485200
rect 359884 485188 359890 485240
rect 44818 485120 44824 485172
rect 44876 485160 44882 485172
rect 130562 485160 130568 485172
rect 44876 485132 130568 485160
rect 44876 485120 44882 485132
rect 130562 485120 130568 485132
rect 130620 485120 130626 485172
rect 261386 485120 261392 485172
rect 261444 485160 261450 485172
rect 368014 485160 368020 485172
rect 261444 485132 368020 485160
rect 261444 485120 261450 485132
rect 368014 485120 368020 485132
rect 368072 485120 368078 485172
rect 46198 485052 46204 485104
rect 46256 485092 46262 485104
rect 133230 485092 133236 485104
rect 46256 485064 133236 485092
rect 46256 485052 46262 485064
rect 133230 485052 133236 485064
rect 133288 485052 133294 485104
rect 159634 485052 159640 485104
rect 159692 485092 159698 485104
rect 214558 485092 214564 485104
rect 159692 485064 214564 485092
rect 159692 485052 159698 485064
rect 214558 485052 214564 485064
rect 214616 485052 214622 485104
rect 242894 485052 242900 485104
rect 242952 485092 242958 485104
rect 369118 485092 369124 485104
rect 242952 485064 369124 485092
rect 242952 485052 242958 485064
rect 369118 485052 369124 485064
rect 369176 485052 369182 485104
rect 46750 484984 46756 485036
rect 46808 485024 46814 485036
rect 116946 485024 116952 485036
rect 46808 484996 116952 485024
rect 46808 484984 46814 484996
rect 116946 484984 116952 484996
rect 117004 484984 117010 485036
rect 48222 484916 48228 484968
rect 48280 484956 48286 484968
rect 117866 484956 117872 484968
rect 48280 484928 117872 484956
rect 48280 484916 48286 484928
rect 117866 484916 117872 484928
rect 117924 484916 117930 484968
rect 58802 484848 58808 484900
rect 58860 484888 58866 484900
rect 110782 484888 110788 484900
rect 58860 484860 110788 484888
rect 58860 484848 58866 484860
rect 110782 484848 110788 484860
rect 110840 484848 110846 484900
rect 292206 484304 292212 484356
rect 292264 484344 292270 484356
rect 368198 484344 368204 484356
rect 292264 484316 368204 484344
rect 292264 484304 292270 484316
rect 368198 484304 368204 484316
rect 368256 484304 368262 484356
rect 270218 484236 270224 484288
rect 270276 484276 270282 484288
rect 357066 484276 357072 484288
rect 270276 484248 357072 484276
rect 270276 484236 270282 484248
rect 357066 484236 357072 484248
rect 357124 484236 357130 484288
rect 269758 484168 269764 484220
rect 269816 484208 269822 484220
rect 358722 484208 358728 484220
rect 269816 484180 358728 484208
rect 269816 484168 269822 484180
rect 358722 484168 358728 484180
rect 358780 484168 358786 484220
rect 280798 484100 280804 484152
rect 280856 484140 280862 484152
rect 374454 484140 374460 484152
rect 280856 484112 374460 484140
rect 280856 484100 280862 484112
rect 374454 484100 374460 484112
rect 374512 484100 374518 484152
rect 281258 484032 281264 484084
rect 281316 484072 281322 484084
rect 376570 484072 376576 484084
rect 281316 484044 376576 484072
rect 281316 484032 281322 484044
rect 376570 484032 376576 484044
rect 376628 484032 376634 484084
rect 268930 483964 268936 484016
rect 268988 484004 268994 484016
rect 370958 484004 370964 484016
rect 268988 483976 370964 484004
rect 268988 483964 268994 483976
rect 370958 483964 370964 483976
rect 371016 483964 371022 484016
rect 268470 483896 268476 483948
rect 268528 483936 268534 483948
rect 377306 483936 377312 483948
rect 268528 483908 377312 483936
rect 268528 483896 268534 483908
rect 377306 483896 377312 483908
rect 377364 483896 377370 483948
rect 260558 483828 260564 483880
rect 260616 483868 260622 483880
rect 369394 483868 369400 483880
rect 260616 483840 369400 483868
rect 260616 483828 260622 483840
rect 369394 483828 369400 483840
rect 369452 483828 369458 483880
rect 243354 483760 243360 483812
rect 243412 483800 243418 483812
rect 366542 483800 366548 483812
rect 243412 483772 366548 483800
rect 243412 483760 243418 483772
rect 366542 483760 366548 483772
rect 366600 483760 366606 483812
rect 205450 483692 205456 483744
rect 205508 483732 205514 483744
rect 217318 483732 217324 483744
rect 205508 483704 217324 483732
rect 205508 483692 205514 483704
rect 217318 483692 217324 483704
rect 217376 483692 217382 483744
rect 231854 483692 231860 483744
rect 231912 483732 231918 483744
rect 366450 483732 366456 483744
rect 231912 483704 366456 483732
rect 231912 483692 231918 483704
rect 366450 483692 366456 483704
rect 366508 483692 366514 483744
rect 58710 483624 58716 483676
rect 58768 483664 58774 483676
rect 96246 483664 96252 483676
rect 58768 483636 96252 483664
rect 58768 483624 58774 483636
rect 96246 483624 96252 483636
rect 96304 483624 96310 483676
rect 184290 483624 184296 483676
rect 184348 483664 184354 483676
rect 214834 483664 214840 483676
rect 184348 483636 214840 483664
rect 184348 483624 184354 483636
rect 214834 483624 214840 483636
rect 214892 483624 214898 483676
rect 238478 483624 238484 483676
rect 238536 483664 238542 483676
rect 378778 483664 378784 483676
rect 238536 483636 378784 483664
rect 238536 483624 238542 483636
rect 378778 483624 378784 483636
rect 378836 483624 378842 483676
rect 57698 482944 57704 482996
rect 57756 482984 57762 482996
rect 114278 482984 114284 482996
rect 57756 482956 114284 482984
rect 57756 482944 57762 482956
rect 114278 482944 114284 482956
rect 114336 482944 114342 482996
rect 59630 482876 59636 482928
rect 59688 482916 59694 482928
rect 127986 482916 127992 482928
rect 59688 482888 127992 482916
rect 59688 482876 59694 482888
rect 127986 482876 127992 482888
rect 128044 482876 128050 482928
rect 58434 482808 58440 482860
rect 58492 482848 58498 482860
rect 128814 482848 128820 482860
rect 58492 482820 128820 482848
rect 58492 482808 58498 482820
rect 128814 482808 128820 482820
rect 128872 482808 128878 482860
rect 50338 482740 50344 482792
rect 50396 482780 50402 482792
rect 126238 482780 126244 482792
rect 50396 482752 126244 482780
rect 50396 482740 50402 482752
rect 126238 482740 126244 482752
rect 126296 482740 126302 482792
rect 43622 482672 43628 482724
rect 43680 482712 43686 482724
rect 123570 482712 123576 482724
rect 43680 482684 123576 482712
rect 43680 482672 43686 482684
rect 123570 482672 123576 482684
rect 123628 482672 123634 482724
rect 43806 482604 43812 482656
rect 43864 482644 43870 482656
rect 124398 482644 124404 482656
rect 43864 482616 124404 482644
rect 43864 482604 43870 482616
rect 124398 482604 124404 482616
rect 124456 482604 124462 482656
rect 43898 482536 43904 482588
rect 43956 482576 43962 482588
rect 124858 482576 124864 482588
rect 43956 482548 124864 482576
rect 43956 482536 43962 482548
rect 124858 482536 124864 482548
rect 124916 482536 124922 482588
rect 43714 482468 43720 482520
rect 43772 482508 43778 482520
rect 125778 482508 125784 482520
rect 43772 482480 125784 482508
rect 43772 482468 43778 482480
rect 125778 482468 125784 482480
rect 125836 482468 125842 482520
rect 40954 482400 40960 482452
rect 41012 482440 41018 482452
rect 123110 482440 123116 482452
rect 41012 482412 123116 482440
rect 41012 482400 41018 482412
rect 123110 482400 123116 482412
rect 123168 482400 123174 482452
rect 253014 482400 253020 482452
rect 253072 482440 253078 482452
rect 375006 482440 375012 482452
rect 253072 482412 375012 482440
rect 253072 482400 253078 482412
rect 375006 482400 375012 482412
rect 375064 482400 375070 482452
rect 48774 482332 48780 482384
rect 48832 482372 48838 482384
rect 133690 482372 133696 482384
rect 48832 482344 133696 482372
rect 48832 482332 48838 482344
rect 133690 482332 133696 482344
rect 133748 482332 133754 482384
rect 245102 482332 245108 482384
rect 245160 482372 245166 482384
rect 370590 482372 370596 482384
rect 245160 482344 370596 482372
rect 245160 482332 245166 482344
rect 370590 482332 370596 482344
rect 370648 482332 370654 482384
rect 43254 482264 43260 482316
rect 43312 482304 43318 482316
rect 143810 482304 143816 482316
rect 43312 482276 143816 482304
rect 43312 482264 43318 482276
rect 143810 482264 143816 482276
rect 143868 482264 143874 482316
rect 171962 482264 171968 482316
rect 172020 482304 172026 482316
rect 203518 482304 203524 482316
rect 172020 482276 203524 482304
rect 172020 482264 172026 482276
rect 203518 482264 203524 482276
rect 203576 482264 203582 482316
rect 239858 482264 239864 482316
rect 239916 482304 239922 482316
rect 378870 482304 378876 482316
rect 239916 482276 378876 482304
rect 239916 482264 239922 482276
rect 378870 482264 378876 482276
rect 378928 482264 378934 482316
rect 292666 481448 292672 481500
rect 292724 481488 292730 481500
rect 357986 481488 357992 481500
rect 292724 481460 357992 481488
rect 292724 481448 292730 481460
rect 357986 481448 357992 481460
rect 358044 481448 358050 481500
rect 291838 481380 291844 481432
rect 291896 481420 291902 481432
rect 365622 481420 365628 481432
rect 291896 481392 365628 481420
rect 291896 481380 291902 481392
rect 365622 481380 365628 481392
rect 365680 481380 365686 481432
rect 289630 481312 289636 481364
rect 289688 481352 289694 481364
rect 368382 481352 368388 481364
rect 289688 481324 368388 481352
rect 289688 481312 289694 481324
rect 368382 481312 368388 481324
rect 368440 481312 368446 481364
rect 279050 481244 279056 481296
rect 279108 481284 279114 481296
rect 360838 481284 360844 481296
rect 279108 481256 360844 481284
rect 279108 481244 279114 481256
rect 360838 481244 360844 481256
rect 360896 481244 360902 481296
rect 279510 481176 279516 481228
rect 279568 481216 279574 481228
rect 364150 481216 364156 481228
rect 279568 481188 364156 481216
rect 279568 481176 279574 481188
rect 364150 481176 364156 481188
rect 364208 481176 364214 481228
rect 279878 481108 279884 481160
rect 279936 481148 279942 481160
rect 367002 481148 367008 481160
rect 279936 481120 367008 481148
rect 279936 481108 279942 481120
rect 367002 481108 367008 481120
rect 367060 481108 367066 481160
rect 274634 481040 274640 481092
rect 274692 481080 274698 481092
rect 364886 481080 364892 481092
rect 274692 481052 364892 481080
rect 274692 481040 274698 481052
rect 364886 481040 364892 481052
rect 364944 481040 364950 481092
rect 177758 480972 177764 481024
rect 177816 481012 177822 481024
rect 202322 481012 202328 481024
rect 177816 480984 202328 481012
rect 177816 480972 177822 480984
rect 202322 480972 202328 480984
rect 202380 480972 202386 481024
rect 275094 480972 275100 481024
rect 275152 481012 275158 481024
rect 367646 481012 367652 481024
rect 275152 480984 367652 481012
rect 275152 480972 275158 480984
rect 367646 480972 367652 480984
rect 367704 480972 367710 481024
rect 162302 480904 162308 480956
rect 162360 480944 162366 480956
rect 204898 480944 204904 480956
rect 162360 480916 204904 480944
rect 162360 480904 162366 480916
rect 204898 480904 204904 480916
rect 204956 480904 204962 480956
rect 258810 480904 258816 480956
rect 258868 480944 258874 480956
rect 365438 480944 365444 480956
rect 258868 480916 365444 480944
rect 258868 480904 258874 480916
rect 365438 480904 365444 480916
rect 365496 480904 365502 480956
rect 254394 479680 254400 479732
rect 254452 479720 254458 479732
rect 373626 479720 373632 479732
rect 254452 479692 373632 479720
rect 254452 479680 254458 479692
rect 373626 479680 373632 479692
rect 373684 479680 373690 479732
rect 176378 479612 176384 479664
rect 176436 479652 176442 479664
rect 209498 479652 209504 479664
rect 176436 479624 209504 479652
rect 176436 479612 176442 479624
rect 209498 479612 209504 479624
rect 209556 479612 209562 479664
rect 238110 479612 238116 479664
rect 238168 479652 238174 479664
rect 376110 479652 376116 479664
rect 238168 479624 376116 479652
rect 238168 479612 238174 479624
rect 376110 479612 376116 479624
rect 376168 479612 376174 479664
rect 166258 479544 166264 479596
rect 166316 479584 166322 479596
rect 213362 479584 213368 479596
rect 166316 479556 213368 479584
rect 166316 479544 166322 479556
rect 213362 479544 213368 479556
rect 213420 479544 213426 479596
rect 227898 479544 227904 479596
rect 227956 479584 227962 479596
rect 367738 479584 367744 479596
rect 227956 479556 367744 479584
rect 227956 479544 227962 479556
rect 367738 479544 367744 479556
rect 367796 479544 367802 479596
rect 3510 479476 3516 479528
rect 3568 479516 3574 479528
rect 309778 479516 309784 479528
rect 3568 479488 309784 479516
rect 3568 479476 3574 479488
rect 309778 479476 309784 479488
rect 309836 479476 309842 479528
rect 291378 478796 291384 478848
rect 291436 478836 291442 478848
rect 362678 478836 362684 478848
rect 291436 478808 362684 478836
rect 291436 478796 291442 478808
rect 362678 478796 362684 478808
rect 362736 478796 362742 478848
rect 289170 478728 289176 478780
rect 289228 478768 289234 478780
rect 360746 478768 360752 478780
rect 289228 478740 360752 478768
rect 289228 478728 289234 478740
rect 360746 478728 360752 478740
rect 360804 478728 360810 478780
rect 278590 478660 278596 478712
rect 278648 478700 278654 478712
rect 357158 478700 357164 478712
rect 278648 478672 357164 478700
rect 278648 478660 278654 478672
rect 357158 478660 357164 478672
rect 357216 478660 357222 478712
rect 278130 478592 278136 478644
rect 278188 478632 278194 478644
rect 362770 478632 362776 478644
rect 278188 478604 362776 478632
rect 278188 478592 278194 478604
rect 362770 478592 362776 478604
rect 362828 478592 362834 478644
rect 273714 478524 273720 478576
rect 273772 478564 273778 478576
rect 360654 478564 360660 478576
rect 273772 478536 360660 478564
rect 273772 478524 273778 478536
rect 360654 478524 360660 478536
rect 360712 478524 360718 478576
rect 273254 478456 273260 478508
rect 273312 478496 273318 478508
rect 364242 478496 364248 478508
rect 273312 478468 364248 478496
rect 273312 478456 273318 478468
rect 364242 478456 364248 478468
rect 364300 478456 364306 478508
rect 256142 478388 256148 478440
rect 256200 478428 256206 478440
rect 356882 478428 356888 478440
rect 256200 478400 356888 478428
rect 256200 478388 256206 478400
rect 356882 478388 356888 478400
rect 356940 478388 356946 478440
rect 256602 478320 256608 478372
rect 256660 478360 256666 478372
rect 358446 478360 358452 478372
rect 256660 478332 358452 478360
rect 256660 478320 256666 478332
rect 358446 478320 358452 478332
rect 358504 478320 358510 478372
rect 260098 478252 260104 478304
rect 260156 478292 260162 478304
rect 362494 478292 362500 478304
rect 260156 478264 362500 478292
rect 260156 478252 260162 478264
rect 362494 478252 362500 478264
rect 362552 478252 362558 478304
rect 159266 478184 159272 478236
rect 159324 478224 159330 478236
rect 204990 478224 204996 478236
rect 159324 478196 204996 478224
rect 159324 478184 159330 478196
rect 204990 478184 204996 478196
rect 205048 478184 205054 478236
rect 246022 478184 246028 478236
rect 246080 478224 246086 478236
rect 369210 478224 369216 478236
rect 246080 478196 369216 478224
rect 246080 478184 246086 478196
rect 369210 478184 369216 478196
rect 369268 478184 369274 478236
rect 3602 478116 3608 478168
rect 3660 478156 3666 478168
rect 434806 478156 434812 478168
rect 3660 478128 434812 478156
rect 3660 478116 3666 478128
rect 434806 478116 434812 478128
rect 434864 478116 434870 478168
rect 178586 476892 178592 476944
rect 178644 476932 178650 476944
rect 200850 476932 200856 476944
rect 178644 476904 200856 476932
rect 178644 476892 178650 476904
rect 200850 476892 200856 476904
rect 200908 476892 200914 476944
rect 259638 476892 259644 476944
rect 259696 476932 259702 476944
rect 370866 476932 370872 476944
rect 259696 476904 370872 476932
rect 259696 476892 259702 476904
rect 370866 476892 370872 476904
rect 370924 476892 370930 476944
rect 163222 476824 163228 476876
rect 163280 476864 163286 476876
rect 210602 476864 210608 476876
rect 163280 476836 210608 476864
rect 163280 476824 163286 476836
rect 210602 476824 210608 476836
rect 210660 476824 210666 476876
rect 244642 476824 244648 476876
rect 244700 476864 244706 476876
rect 371878 476864 371884 476876
rect 244700 476836 371884 476864
rect 244700 476824 244706 476836
rect 371878 476824 371884 476836
rect 371936 476824 371942 476876
rect 62758 476756 62764 476808
rect 62816 476796 62822 476808
rect 199102 476796 199108 476808
rect 62816 476768 199108 476796
rect 62816 476756 62822 476768
rect 199102 476756 199108 476768
rect 199160 476756 199166 476808
rect 232774 476756 232780 476808
rect 232832 476796 232838 476808
rect 364978 476796 364984 476808
rect 232832 476768 364984 476796
rect 232832 476756 232838 476768
rect 364978 476756 364984 476768
rect 365036 476756 365042 476808
rect 290918 475804 290924 475856
rect 290976 475844 290982 475856
rect 361390 475844 361396 475856
rect 290976 475816 361396 475844
rect 290976 475804 290982 475816
rect 361390 475804 361396 475816
rect 361448 475804 361454 475856
rect 285674 475736 285680 475788
rect 285732 475776 285738 475788
rect 358078 475776 358084 475788
rect 285732 475748 358084 475776
rect 285732 475736 285738 475748
rect 358078 475736 358084 475748
rect 358136 475736 358142 475788
rect 277670 475668 277676 475720
rect 277728 475708 277734 475720
rect 364794 475708 364800 475720
rect 277728 475680 364800 475708
rect 277728 475668 277734 475680
rect 364794 475668 364800 475680
rect 364852 475668 364858 475720
rect 266262 475600 266268 475652
rect 266320 475640 266326 475652
rect 358538 475640 358544 475652
rect 266320 475612 358544 475640
rect 266320 475600 266326 475612
rect 358538 475600 358544 475612
rect 358596 475600 358602 475652
rect 272886 475532 272892 475584
rect 272944 475572 272950 475584
rect 366266 475572 366272 475584
rect 272944 475544 366272 475572
rect 272944 475532 272950 475544
rect 366266 475532 366272 475544
rect 366324 475532 366330 475584
rect 170674 475464 170680 475516
rect 170732 475504 170738 475516
rect 211890 475504 211896 475516
rect 170732 475476 211896 475504
rect 170732 475464 170738 475476
rect 211890 475464 211896 475476
rect 211948 475464 211954 475516
rect 253934 475464 253940 475516
rect 253992 475504 253998 475516
rect 361206 475504 361212 475516
rect 253992 475476 361212 475504
rect 253992 475464 253998 475476
rect 361206 475464 361212 475476
rect 361264 475464 361270 475516
rect 148226 475396 148232 475448
rect 148284 475436 148290 475448
rect 213178 475436 213184 475448
rect 148284 475408 213184 475436
rect 148284 475396 148290 475408
rect 213178 475396 213184 475408
rect 213236 475396 213242 475448
rect 265342 475396 265348 475448
rect 265400 475436 265406 475448
rect 376294 475436 376300 475448
rect 265400 475408 376300 475436
rect 265400 475396 265406 475408
rect 376294 475396 376300 475408
rect 376352 475396 376358 475448
rect 61930 475328 61936 475380
rect 61988 475368 61994 475380
rect 199194 475368 199200 475380
rect 61988 475340 199200 475368
rect 61988 475328 61994 475340
rect 199194 475328 199200 475340
rect 199252 475328 199258 475380
rect 245562 475328 245568 475380
rect 245620 475368 245626 475380
rect 362310 475368 362316 475380
rect 245620 475340 362316 475368
rect 245620 475328 245626 475340
rect 362310 475328 362316 475340
rect 362368 475328 362374 475380
rect 43346 474648 43352 474700
rect 43404 474688 43410 474700
rect 72510 474688 72516 474700
rect 43404 474660 72516 474688
rect 43404 474648 43410 474660
rect 72510 474648 72516 474660
rect 72568 474648 72574 474700
rect 51718 474580 51724 474632
rect 51776 474620 51782 474632
rect 99742 474620 99748 474632
rect 51776 474592 99748 474620
rect 51776 474580 51782 474592
rect 99742 474580 99748 474592
rect 99800 474580 99806 474632
rect 50246 474512 50252 474564
rect 50304 474552 50310 474564
rect 98914 474552 98920 474564
rect 50304 474524 98920 474552
rect 50304 474512 50310 474524
rect 98914 474512 98920 474524
rect 98972 474512 98978 474564
rect 51626 474444 51632 474496
rect 51684 474484 51690 474496
rect 100662 474484 100668 474496
rect 51684 474456 100668 474484
rect 51684 474444 51690 474456
rect 100662 474444 100668 474456
rect 100720 474444 100726 474496
rect 45186 474376 45192 474428
rect 45244 474416 45250 474428
rect 105078 474416 105084 474428
rect 45244 474388 105084 474416
rect 45244 474376 45250 474388
rect 105078 474376 105084 474388
rect 105136 474376 105142 474428
rect 45094 474308 45100 474360
rect 45152 474348 45158 474360
rect 105906 474348 105912 474360
rect 45152 474320 105912 474348
rect 45152 474308 45158 474320
rect 105906 474308 105912 474320
rect 105964 474308 105970 474360
rect 43530 474240 43536 474292
rect 43588 474280 43594 474292
rect 103698 474280 103704 474292
rect 43588 474252 103704 474280
rect 43588 474240 43594 474252
rect 103698 474240 103704 474252
rect 103756 474240 103762 474292
rect 193950 474240 193956 474292
rect 194008 474280 194014 474292
rect 205726 474280 205732 474292
rect 194008 474252 205732 474280
rect 194008 474240 194014 474252
rect 205726 474240 205732 474252
rect 205784 474240 205790 474292
rect 45002 474172 45008 474224
rect 45060 474212 45066 474224
rect 105538 474212 105544 474224
rect 45060 474184 105544 474212
rect 45060 474172 45066 474184
rect 105538 474172 105544 474184
rect 105596 474172 105602 474224
rect 186130 474172 186136 474224
rect 186188 474212 186194 474224
rect 213546 474212 213552 474224
rect 186188 474184 213552 474212
rect 186188 474172 186194 474184
rect 213546 474172 213552 474184
rect 213604 474172 213610 474224
rect 287790 474172 287796 474224
rect 287848 474212 287854 474224
rect 369026 474212 369032 474224
rect 287848 474184 369032 474212
rect 287848 474172 287854 474184
rect 369026 474172 369032 474184
rect 369084 474172 369090 474224
rect 45370 474104 45376 474156
rect 45428 474144 45434 474156
rect 106366 474144 106372 474156
rect 45428 474116 106372 474144
rect 45428 474104 45434 474116
rect 106366 474104 106372 474116
rect 106424 474104 106430 474156
rect 139854 474104 139860 474156
rect 139912 474144 139918 474156
rect 207290 474144 207296 474156
rect 139912 474116 207296 474144
rect 139912 474104 139918 474116
rect 207290 474104 207296 474116
rect 207348 474104 207354 474156
rect 259178 474104 259184 474156
rect 259236 474144 259242 474156
rect 372062 474144 372068 474156
rect 259236 474116 372068 474144
rect 259236 474104 259242 474116
rect 372062 474104 372068 474116
rect 372120 474104 372126 474156
rect 45278 474036 45284 474088
rect 45336 474076 45342 474088
rect 106826 474076 106832 474088
rect 45336 474048 106832 474076
rect 45336 474036 45342 474048
rect 106826 474036 106832 474048
rect 106884 474036 106890 474088
rect 127526 474036 127532 474088
rect 127584 474076 127590 474088
rect 204346 474076 204352 474088
rect 127584 474048 204352 474076
rect 127584 474036 127590 474048
rect 204346 474036 204352 474048
rect 204404 474036 204410 474088
rect 237190 474036 237196 474088
rect 237248 474076 237254 474088
rect 362402 474076 362408 474088
rect 237248 474048 362408 474076
rect 237248 474036 237254 474048
rect 362402 474036 362408 474048
rect 362460 474036 362466 474088
rect 61470 473968 61476 474020
rect 61528 474008 61534 474020
rect 199470 474008 199476 474020
rect 61528 473980 199476 474008
rect 61528 473968 61534 473980
rect 199470 473968 199476 473980
rect 199528 473968 199534 474020
rect 248230 473968 248236 474020
rect 248288 474008 248294 474020
rect 376202 474008 376208 474020
rect 248288 473980 376208 474008
rect 248288 473968 248294 473980
rect 376202 473968 376208 473980
rect 376260 473968 376266 474020
rect 43438 473900 43444 473952
rect 43496 473940 43502 473952
rect 72418 473940 72424 473952
rect 43496 473912 72424 473940
rect 43496 473900 43502 473912
rect 72418 473900 72424 473912
rect 72476 473900 72482 473952
rect 264054 473220 264060 473272
rect 264112 473260 264118 473272
rect 362586 473260 362592 473272
rect 264112 473232 362592 473260
rect 264112 473220 264118 473232
rect 362586 473220 362592 473232
rect 362644 473220 362650 473272
rect 264514 473152 264520 473204
rect 264572 473192 264578 473204
rect 363966 473192 363972 473204
rect 264572 473164 363972 473192
rect 264572 473152 264578 473164
rect 363966 473152 363972 473164
rect 364024 473152 364030 473204
rect 265802 473084 265808 473136
rect 265860 473124 265866 473136
rect 365530 473124 365536 473136
rect 265860 473096 365536 473124
rect 265860 473084 265866 473096
rect 365530 473084 365536 473096
rect 365588 473084 365594 473136
rect 267550 473016 267556 473068
rect 267608 473056 267614 473068
rect 375190 473056 375196 473068
rect 267608 473028 375196 473056
rect 267608 473016 267614 473028
rect 375190 473016 375196 473028
rect 375248 473016 375254 473068
rect 264974 472948 264980 473000
rect 265032 472988 265038 473000
rect 373718 472988 373724 473000
rect 265032 472960 373724 472988
rect 265032 472948 265038 472960
rect 373718 472948 373724 472960
rect 373776 472948 373782 473000
rect 261846 472880 261852 472932
rect 261904 472920 261910 472932
rect 376386 472920 376392 472932
rect 261904 472892 376392 472920
rect 261904 472880 261910 472892
rect 376386 472880 376392 472892
rect 376444 472880 376450 472932
rect 187418 472812 187424 472864
rect 187476 472852 187482 472864
rect 207750 472852 207756 472864
rect 187476 472824 207756 472852
rect 187476 472812 187482 472824
rect 207750 472812 207756 472824
rect 207808 472812 207814 472864
rect 241606 472812 241612 472864
rect 241664 472852 241670 472864
rect 370682 472852 370688 472864
rect 241664 472824 370688 472852
rect 241664 472812 241670 472824
rect 370682 472812 370688 472824
rect 370740 472812 370746 472864
rect 176010 472744 176016 472796
rect 176068 472784 176074 472796
rect 205082 472784 205088 472796
rect 176068 472756 205088 472784
rect 176068 472744 176074 472756
rect 205082 472744 205088 472756
rect 205140 472744 205146 472796
rect 205910 472744 205916 472796
rect 205968 472784 205974 472796
rect 217686 472784 217692 472796
rect 205968 472756 217692 472784
rect 205968 472744 205974 472756
rect 217686 472744 217692 472756
rect 217744 472744 217750 472796
rect 227070 472744 227076 472796
rect 227128 472784 227134 472796
rect 362218 472784 362224 472796
rect 227128 472756 362224 472784
rect 227128 472744 227134 472756
rect 362218 472744 362224 472756
rect 362276 472744 362282 472796
rect 176838 472676 176844 472728
rect 176896 472716 176902 472728
rect 210694 472716 210700 472728
rect 176896 472688 210700 472716
rect 176896 472676 176902 472688
rect 210694 472676 210700 472688
rect 210752 472676 210758 472728
rect 222654 472676 222660 472728
rect 222712 472716 222718 472728
rect 365070 472716 365076 472728
rect 222712 472688 365076 472716
rect 222712 472676 222718 472688
rect 365070 472676 365076 472688
rect 365128 472676 365134 472728
rect 57606 472608 57612 472660
rect 57664 472648 57670 472660
rect 113910 472648 113916 472660
rect 57664 472620 113916 472648
rect 57664 472608 57670 472620
rect 113910 472608 113916 472620
rect 113968 472608 113974 472660
rect 161014 472608 161020 472660
rect 161072 472648 161078 472660
rect 206278 472648 206284 472660
rect 161072 472620 206284 472648
rect 161072 472608 161078 472620
rect 206278 472608 206284 472620
rect 206336 472608 206342 472660
rect 227530 472608 227536 472660
rect 227588 472648 227594 472660
rect 374730 472648 374736 472660
rect 227588 472620 374736 472648
rect 227588 472608 227594 472620
rect 374730 472608 374736 472620
rect 374788 472608 374794 472660
rect 50982 471928 50988 471980
rect 51040 471968 51046 471980
rect 82998 471968 83004 471980
rect 51040 471940 83004 471968
rect 51040 471928 51046 471940
rect 82998 471928 83004 471940
rect 83056 471928 83062 471980
rect 193122 471928 193128 471980
rect 193180 471968 193186 471980
rect 214926 471968 214932 471980
rect 193180 471940 214932 471968
rect 193180 471928 193186 471940
rect 214926 471928 214932 471940
rect 214984 471928 214990 471980
rect 53466 471860 53472 471912
rect 53524 471900 53530 471912
rect 85666 471900 85672 471912
rect 53524 471872 85672 471900
rect 53524 471860 53530 471872
rect 85666 471860 85672 471872
rect 85724 471860 85730 471912
rect 190914 471860 190920 471912
rect 190972 471900 190978 471912
rect 215846 471900 215852 471912
rect 190972 471872 215852 471900
rect 190972 471860 190978 471872
rect 215846 471860 215852 471872
rect 215904 471860 215910 471912
rect 299750 471860 299756 471912
rect 299808 471900 299814 471912
rect 373074 471900 373080 471912
rect 299808 471872 373080 471900
rect 299808 471860 299814 471872
rect 373074 471860 373080 471872
rect 373132 471860 373138 471912
rect 56318 471792 56324 471844
rect 56376 471832 56382 471844
rect 90082 471832 90088 471844
rect 56376 471804 90088 471832
rect 56376 471792 56382 471804
rect 90082 471792 90088 471804
rect 90140 471792 90146 471844
rect 183002 471792 183008 471844
rect 183060 471832 183066 471844
rect 216122 471832 216128 471844
rect 183060 471804 216128 471832
rect 183060 471792 183066 471804
rect 216122 471792 216128 471804
rect 216180 471792 216186 471844
rect 294874 471792 294880 471844
rect 294932 471832 294938 471844
rect 372430 471832 372436 471844
rect 294932 471804 372436 471832
rect 294932 471792 294938 471804
rect 372430 471792 372436 471804
rect 372488 471792 372494 471844
rect 49326 471724 49332 471776
rect 49384 471764 49390 471776
rect 83458 471764 83464 471776
rect 49384 471736 83464 471764
rect 49384 471724 49390 471736
rect 83458 471724 83464 471736
rect 83516 471724 83522 471776
rect 175090 471724 175096 471776
rect 175148 471764 175154 471776
rect 212074 471764 212080 471776
rect 175148 471736 212080 471764
rect 175148 471724 175154 471736
rect 212074 471724 212080 471736
rect 212132 471724 212138 471776
rect 286042 471724 286048 471776
rect 286100 471764 286106 471776
rect 366174 471764 366180 471776
rect 286100 471736 366180 471764
rect 286100 471724 286106 471736
rect 366174 471724 366180 471736
rect 366232 471724 366238 471776
rect 58894 471656 58900 471708
rect 58952 471696 58958 471708
rect 95786 471696 95792 471708
rect 58952 471668 95792 471696
rect 58952 471656 58958 471668
rect 95786 471656 95792 471668
rect 95844 471656 95850 471708
rect 179046 471656 179052 471708
rect 179104 471696 179110 471708
rect 216766 471696 216772 471708
rect 179104 471668 216772 471696
rect 179104 471656 179110 471668
rect 216766 471656 216772 471668
rect 216824 471656 216830 471708
rect 293586 471656 293592 471708
rect 293644 471696 293650 471708
rect 375926 471696 375932 471708
rect 293644 471668 375932 471696
rect 293644 471656 293650 471668
rect 375926 471656 375932 471668
rect 375984 471656 375990 471708
rect 56870 471588 56876 471640
rect 56928 471628 56934 471640
rect 102870 471628 102876 471640
rect 56928 471600 102876 471628
rect 56928 471588 56934 471600
rect 102870 471588 102876 471600
rect 102928 471588 102934 471640
rect 140314 471588 140320 471640
rect 140372 471628 140378 471640
rect 196894 471628 196900 471640
rect 140372 471600 196900 471628
rect 140372 471588 140378 471600
rect 196894 471588 196900 471600
rect 196952 471588 196958 471640
rect 287422 471588 287428 471640
rect 287480 471628 287486 471640
rect 370406 471628 370412 471640
rect 287480 471600 370412 471628
rect 287480 471588 287486 471600
rect 370406 471588 370412 471600
rect 370464 471588 370470 471640
rect 54662 471520 54668 471572
rect 54720 471560 54726 471572
rect 102410 471560 102416 471572
rect 54720 471532 102416 471560
rect 54720 471520 54726 471532
rect 102410 471520 102416 471532
rect 102468 471520 102474 471572
rect 141142 471520 141148 471572
rect 141200 471560 141206 471572
rect 200390 471560 200396 471572
rect 141200 471532 200396 471560
rect 141200 471520 141206 471532
rect 200390 471520 200396 471532
rect 200448 471520 200454 471572
rect 286502 471520 286508 471572
rect 286560 471560 286566 471572
rect 369762 471560 369768 471572
rect 286560 471532 369768 471560
rect 286560 471520 286566 471532
rect 369762 471520 369768 471532
rect 369820 471520 369826 471572
rect 53190 471452 53196 471504
rect 53248 471492 53254 471504
rect 101122 471492 101128 471504
rect 53248 471464 101128 471492
rect 53248 471452 53254 471464
rect 101122 471452 101128 471464
rect 101180 471452 101186 471504
rect 141602 471452 141608 471504
rect 141660 471492 141666 471504
rect 204622 471492 204628 471504
rect 141660 471464 204628 471492
rect 141660 471452 141666 471464
rect 204622 471452 204628 471464
rect 204680 471452 204686 471504
rect 286962 471452 286968 471504
rect 287020 471492 287026 471504
rect 375282 471492 375288 471504
rect 287020 471464 375288 471492
rect 287020 471452 287026 471464
rect 375282 471452 375288 471464
rect 375340 471452 375346 471504
rect 52822 471384 52828 471436
rect 52880 471424 52886 471436
rect 101490 471424 101496 471436
rect 52880 471396 101496 471424
rect 52880 471384 52886 471396
rect 101490 471384 101496 471396
rect 101548 471384 101554 471436
rect 142062 471384 142068 471436
rect 142120 471424 142126 471436
rect 205818 471424 205824 471436
rect 142120 471396 205824 471424
rect 142120 471384 142126 471396
rect 205818 471384 205824 471396
rect 205876 471384 205882 471436
rect 282546 471384 282552 471436
rect 282604 471424 282610 471436
rect 374546 471424 374552 471436
rect 282604 471396 374552 471424
rect 282604 471384 282610 471396
rect 374546 471384 374552 471396
rect 374604 471384 374610 471436
rect 56686 471316 56692 471368
rect 56744 471356 56750 471368
rect 114738 471356 114744 471368
rect 56744 471328 114744 471356
rect 56744 471316 56750 471328
rect 114738 471316 114744 471328
rect 114796 471316 114802 471368
rect 127066 471316 127072 471368
rect 127124 471356 127130 471368
rect 202874 471356 202880 471368
rect 127124 471328 202880 471356
rect 127124 471316 127130 471328
rect 202874 471316 202880 471328
rect 202932 471316 202938 471368
rect 271506 471316 271512 471368
rect 271564 471356 271570 471368
rect 371786 471356 371792 471368
rect 271564 471328 371792 471356
rect 271564 471316 271570 471328
rect 371786 471316 371792 471328
rect 371844 471316 371850 471368
rect 42610 471248 42616 471300
rect 42668 471288 42674 471300
rect 104158 471288 104164 471300
rect 42668 471260 104164 471288
rect 42668 471248 42674 471260
rect 104158 471248 104164 471260
rect 104216 471248 104222 471300
rect 109494 471248 109500 471300
rect 109552 471288 109558 471300
rect 202966 471288 202972 471300
rect 109552 471260 202972 471288
rect 109552 471248 109558 471260
rect 202966 471248 202972 471260
rect 203024 471248 203030 471300
rect 271138 471248 271144 471300
rect 271196 471288 271202 471300
rect 373166 471288 373172 471300
rect 271196 471260 373172 471288
rect 271196 471248 271202 471260
rect 373166 471248 373172 471260
rect 373224 471248 373230 471300
rect 52086 471180 52092 471232
rect 52144 471220 52150 471232
rect 83918 471220 83924 471232
rect 52144 471192 83924 471220
rect 52144 471180 52150 471192
rect 83918 471180 83924 471192
rect 83976 471180 83982 471232
rect 191374 471180 191380 471232
rect 191432 471220 191438 471232
rect 210234 471220 210240 471232
rect 191432 471192 210240 471220
rect 191432 471180 191438 471192
rect 210234 471180 210240 471192
rect 210292 471180 210298 471232
rect 44726 471112 44732 471164
rect 44784 471152 44790 471164
rect 65426 471152 65432 471164
rect 44784 471124 65432 471152
rect 44784 471112 44790 471124
rect 65426 471112 65432 471124
rect 65484 471112 65490 471164
rect 188706 471112 188712 471164
rect 188764 471152 188770 471164
rect 200758 471152 200764 471164
rect 188764 471124 200764 471152
rect 188764 471112 188770 471124
rect 200758 471112 200764 471124
rect 200816 471112 200822 471164
rect 47670 471044 47676 471096
rect 47728 471084 47734 471096
rect 64966 471084 64972 471096
rect 47728 471056 64972 471084
rect 47728 471044 47734 471056
rect 64966 471044 64972 471056
rect 65024 471044 65030 471096
rect 193858 470568 193864 470620
rect 193916 470608 193922 470620
rect 201862 470608 201868 470620
rect 193916 470580 201868 470608
rect 193916 470568 193922 470580
rect 201862 470568 201868 470580
rect 201920 470568 201926 470620
rect 283466 470500 283472 470552
rect 283524 470540 283530 470552
rect 360010 470540 360016 470552
rect 283524 470512 360016 470540
rect 283524 470500 283530 470512
rect 360010 470500 360016 470512
rect 360068 470500 360074 470552
rect 283006 470432 283012 470484
rect 283064 470472 283070 470484
rect 359918 470472 359924 470484
rect 283064 470444 359924 470472
rect 283064 470432 283070 470444
rect 359918 470432 359924 470444
rect 359976 470432 359982 470484
rect 281626 470364 281632 470416
rect 281684 470404 281690 470416
rect 359642 470404 359648 470416
rect 281684 470376 359648 470404
rect 281684 470364 281690 470376
rect 359642 470364 359648 470376
rect 359700 470364 359706 470416
rect 298002 470296 298008 470348
rect 298060 470336 298066 470348
rect 378226 470336 378232 470348
rect 298060 470308 378232 470336
rect 298060 470296 298066 470308
rect 378226 470296 378232 470308
rect 378284 470296 378290 470348
rect 293126 470228 293132 470280
rect 293184 470268 293190 470280
rect 376754 470268 376760 470280
rect 293184 470240 376760 470268
rect 293184 470228 293190 470240
rect 376754 470228 376760 470240
rect 376812 470228 376818 470280
rect 293954 470160 293960 470212
rect 294012 470200 294018 470212
rect 379238 470200 379244 470212
rect 294012 470172 379244 470200
rect 294012 470160 294018 470172
rect 379238 470160 379244 470172
rect 379296 470160 379302 470212
rect 284754 470092 284760 470144
rect 284812 470132 284818 470144
rect 377398 470132 377404 470144
rect 284812 470104 377404 470132
rect 284812 470092 284818 470104
rect 377398 470092 377404 470104
rect 377456 470092 377462 470144
rect 175550 470024 175556 470076
rect 175608 470064 175614 470076
rect 210786 470064 210792 470076
rect 175608 470036 210792 470064
rect 175608 470024 175614 470036
rect 210786 470024 210792 470036
rect 210844 470024 210850 470076
rect 282086 470024 282092 470076
rect 282144 470064 282150 470076
rect 379974 470064 379980 470076
rect 282144 470036 379980 470064
rect 282144 470024 282150 470036
rect 379974 470024 379980 470036
rect 380032 470024 380038 470076
rect 173802 469956 173808 470008
rect 173860 469996 173866 470008
rect 209406 469996 209412 470008
rect 173860 469968 209412 469996
rect 173860 469956 173866 469968
rect 209406 469956 209412 469968
rect 209464 469956 209470 470008
rect 250806 469956 250812 470008
rect 250864 469996 250870 470008
rect 365254 469996 365260 470008
rect 250864 469968 365260 469996
rect 250864 469956 250870 469968
rect 365254 469956 365260 469968
rect 365312 469956 365318 470008
rect 178126 469888 178132 469940
rect 178184 469928 178190 469940
rect 215202 469928 215208 469940
rect 178184 469900 215208 469928
rect 178184 469888 178190 469900
rect 215202 469888 215208 469900
rect 215260 469888 215266 469940
rect 251266 469888 251272 469940
rect 251324 469928 251330 469940
rect 373350 469928 373356 469940
rect 251324 469900 373356 469928
rect 251324 469888 251330 469900
rect 373350 469888 373356 469900
rect 373408 469888 373414 469940
rect 57514 469820 57520 469872
rect 57572 469860 57578 469872
rect 112990 469860 112996 469872
rect 57572 469832 112996 469860
rect 57572 469820 57578 469832
rect 112990 469820 112996 469832
rect 113048 469820 113054 469872
rect 161474 469820 161480 469872
rect 161532 469860 161538 469872
rect 207658 469860 207664 469872
rect 161532 469832 207664 469860
rect 161532 469820 161538 469832
rect 207658 469820 207664 469832
rect 207716 469820 207722 469872
rect 240226 469820 240232 469872
rect 240284 469860 240290 469872
rect 366634 469860 366640 469872
rect 240284 469832 366640 469860
rect 240284 469820 240290 469832
rect 366634 469820 366640 469832
rect 366692 469820 366698 469872
rect 295794 469752 295800 469804
rect 295852 469792 295858 469804
rect 357250 469792 357256 469804
rect 295852 469764 357256 469792
rect 295852 469752 295858 469764
rect 357250 469752 357256 469764
rect 357308 469752 357314 469804
rect 56042 469140 56048 469192
rect 56100 469180 56106 469192
rect 81710 469180 81716 469192
rect 56100 469152 81716 469180
rect 56100 469140 56106 469152
rect 81710 469140 81716 469152
rect 81768 469140 81774 469192
rect 186498 469140 186504 469192
rect 186556 469180 186562 469192
rect 206462 469180 206468 469192
rect 186556 469152 206468 469180
rect 186556 469140 186562 469152
rect 206462 469140 206468 469152
rect 206520 469140 206526 469192
rect 269298 469140 269304 469192
rect 269356 469180 269362 469192
rect 359458 469180 359464 469192
rect 269356 469152 359464 469180
rect 269356 469140 269362 469152
rect 359458 469140 359464 469152
rect 359516 469140 359522 469192
rect 56134 469072 56140 469124
rect 56192 469112 56198 469124
rect 87874 469112 87880 469124
rect 56192 469084 87880 469112
rect 56192 469072 56198 469084
rect 87874 469072 87880 469084
rect 87932 469072 87938 469124
rect 181714 469072 181720 469124
rect 181772 469112 181778 469124
rect 203794 469112 203800 469124
rect 181772 469084 203800 469112
rect 181772 469072 181778 469084
rect 203794 469072 203800 469084
rect 203852 469072 203858 469124
rect 277302 469072 277308 469124
rect 277360 469112 277366 469124
rect 367554 469112 367560 469124
rect 277360 469084 367560 469112
rect 277360 469072 277366 469084
rect 367554 469072 367560 469084
rect 367612 469072 367618 469124
rect 55030 469004 55036 469056
rect 55088 469044 55094 469056
rect 87046 469044 87052 469056
rect 55088 469016 87052 469044
rect 55088 469004 55094 469016
rect 87046 469004 87052 469016
rect 87104 469004 87110 469056
rect 192662 469004 192668 469056
rect 192720 469044 192726 469056
rect 217962 469044 217968 469056
rect 192720 469016 217968 469044
rect 192720 469004 192726 469016
rect 217962 469004 217968 469016
rect 218020 469004 218026 469056
rect 266722 469004 266728 469056
rect 266780 469044 266786 469056
rect 358630 469044 358636 469056
rect 266780 469016 358636 469044
rect 266780 469004 266786 469016
rect 358630 469004 358636 469016
rect 358688 469004 358694 469056
rect 55950 468936 55956 468988
rect 56008 468976 56014 468988
rect 88794 468976 88800 468988
rect 56008 468948 88800 468976
rect 56008 468936 56014 468948
rect 88794 468936 88800 468948
rect 88852 468936 88858 468988
rect 190454 468936 190460 468988
rect 190512 468976 190518 468988
rect 217502 468976 217508 468988
rect 190512 468948 217508 468976
rect 190512 468936 190518 468948
rect 217502 468936 217508 468948
rect 217560 468936 217566 468988
rect 267090 468936 267096 468988
rect 267148 468976 267154 468988
rect 359550 468976 359556 468988
rect 267148 468948 359556 468976
rect 267148 468936 267154 468948
rect 359550 468936 359556 468948
rect 359608 468936 359614 468988
rect 55858 468868 55864 468920
rect 55916 468908 55922 468920
rect 89622 468908 89628 468920
rect 55916 468880 89628 468908
rect 55916 468868 55922 468880
rect 89622 468868 89628 468880
rect 89680 468868 89686 468920
rect 189626 468868 189632 468920
rect 189684 468908 189690 468920
rect 217594 468908 217600 468920
rect 189684 468880 217600 468908
rect 189684 468868 189690 468880
rect 217594 468868 217600 468880
rect 217652 468868 217658 468920
rect 285214 468868 285220 468920
rect 285272 468908 285278 468920
rect 377766 468908 377772 468920
rect 285272 468880 377772 468908
rect 285272 468868 285278 468880
rect 377766 468868 377772 468880
rect 377824 468868 377830 468920
rect 54938 468800 54944 468852
rect 54996 468840 55002 468852
rect 88334 468840 88340 468852
rect 54996 468812 88340 468840
rect 54996 468800 55002 468812
rect 88334 468800 88340 468812
rect 88392 468800 88398 468852
rect 168466 468800 168472 468852
rect 168524 468840 168530 468852
rect 209314 468840 209320 468852
rect 168524 468812 209320 468840
rect 168524 468800 168530 468812
rect 209314 468800 209320 468812
rect 209372 468800 209378 468852
rect 275462 468800 275468 468852
rect 275520 468840 275526 468852
rect 370314 468840 370320 468852
rect 275520 468812 370320 468840
rect 275520 468800 275526 468812
rect 370314 468800 370320 468812
rect 370372 468800 370378 468852
rect 51994 468732 52000 468784
rect 52052 468772 52058 468784
rect 86586 468772 86592 468784
rect 52052 468744 86592 468772
rect 52052 468732 52058 468744
rect 86586 468732 86592 468744
rect 86644 468732 86650 468784
rect 169386 468732 169392 468784
rect 169444 468772 169450 468784
rect 211982 468772 211988 468784
rect 169444 468744 211988 468772
rect 169444 468732 169450 468744
rect 211982 468732 211988 468744
rect 212040 468732 212046 468784
rect 272426 468732 272432 468784
rect 272484 468772 272490 468784
rect 368842 468772 368848 468784
rect 272484 468744 368848 468772
rect 272484 468732 272490 468744
rect 368842 468732 368848 468744
rect 368900 468732 368906 468784
rect 57330 468664 57336 468716
rect 57388 468704 57394 468716
rect 113450 468704 113456 468716
rect 57388 468676 113456 468704
rect 57388 468664 57394 468676
rect 113450 468664 113456 468676
rect 113508 468664 113514 468716
rect 170214 468664 170220 468716
rect 170272 468704 170278 468716
rect 213454 468704 213460 468716
rect 170272 468676 213460 468704
rect 170272 468664 170278 468676
rect 213454 468664 213460 468676
rect 213512 468664 213518 468716
rect 271966 468664 271972 468716
rect 272024 468704 272030 468716
rect 372246 468704 372252 468716
rect 272024 468676 372252 468704
rect 272024 468664 272030 468676
rect 372246 468664 372252 468676
rect 372304 468664 372310 468716
rect 53374 468596 53380 468648
rect 53432 468636 53438 468648
rect 87414 468636 87420 468648
rect 53432 468608 87420 468636
rect 53432 468596 53438 468608
rect 87414 468596 87420 468608
rect 87472 468596 87478 468648
rect 109862 468596 109868 468648
rect 109920 468636 109926 468648
rect 197446 468636 197452 468648
rect 109920 468608 197452 468636
rect 109920 468596 109926 468608
rect 197446 468596 197452 468608
rect 197504 468596 197510 468648
rect 268010 468596 268016 468648
rect 268068 468636 268074 468648
rect 377214 468636 377220 468648
rect 268068 468608 377220 468636
rect 268068 468596 268074 468608
rect 377214 468596 377220 468608
rect 377272 468596 377278 468648
rect 53282 468528 53288 468580
rect 53340 468568 53346 468580
rect 94038 468568 94044 468580
rect 53340 468540 94044 468568
rect 53340 468528 53346 468540
rect 94038 468528 94044 468540
rect 94096 468528 94102 468580
rect 108114 468528 108120 468580
rect 108172 468568 108178 468580
rect 200114 468568 200120 468580
rect 108172 468540 200120 468568
rect 108172 468528 108178 468540
rect 200114 468528 200120 468540
rect 200172 468528 200178 468580
rect 255222 468528 255228 468580
rect 255280 468568 255286 468580
rect 366818 468568 366824 468580
rect 255280 468540 366824 468568
rect 255280 468528 255286 468540
rect 366818 468528 366824 468540
rect 366876 468528 366882 468580
rect 49234 468460 49240 468512
rect 49292 468500 49298 468512
rect 94498 468500 94504 468512
rect 49292 468472 94504 468500
rect 49292 468460 49298 468472
rect 94498 468460 94504 468472
rect 94556 468460 94562 468512
rect 108574 468460 108580 468512
rect 108632 468500 108638 468512
rect 201678 468500 201684 468512
rect 108632 468472 201684 468500
rect 108632 468460 108638 468472
rect 201678 468460 201684 468472
rect 201736 468460 201742 468512
rect 254762 468460 254768 468512
rect 254820 468500 254826 468512
rect 375098 468500 375104 468512
rect 254820 468472 375104 468500
rect 254820 468460 254826 468472
rect 375098 468460 375104 468472
rect 375156 468460 375162 468512
rect 49970 468392 49976 468444
rect 50028 468432 50034 468444
rect 68370 468432 68376 468444
rect 50028 468404 68376 468432
rect 50028 468392 50034 468404
rect 68370 468392 68376 468404
rect 68428 468392 68434 468444
rect 193582 468392 193588 468444
rect 193640 468432 193646 468444
rect 213086 468432 213092 468444
rect 193640 468404 213092 468432
rect 193640 468392 193646 468404
rect 213086 468392 213092 468404
rect 213144 468392 213150 468444
rect 298830 468392 298836 468444
rect 298888 468432 298894 468444
rect 378134 468432 378140 468444
rect 298888 468404 378140 468432
rect 298888 468392 298894 468404
rect 378134 468392 378140 468404
rect 378192 468392 378198 468444
rect 46106 468324 46112 468376
rect 46164 468364 46170 468376
rect 64506 468364 64512 468376
rect 46164 468336 64512 468364
rect 46164 468324 46170 468336
rect 64506 468324 64512 468336
rect 64564 468324 64570 468376
rect 183922 468324 183928 468376
rect 183980 468364 183986 468376
rect 200942 468364 200948 468376
rect 183980 468336 200948 468364
rect 183980 468324 183986 468336
rect 200942 468324 200948 468336
rect 201000 468324 201006 468376
rect 290458 468324 290464 468376
rect 290516 468364 290522 468376
rect 363506 468364 363512 468376
rect 290516 468336 363512 468364
rect 290516 468324 290522 468336
rect 363506 468324 363512 468336
rect 363564 468324 363570 468376
rect 59998 468256 60004 468308
rect 60056 468296 60062 468308
rect 67726 468296 67732 468308
rect 60056 468268 67732 468296
rect 60056 468256 60062 468268
rect 67726 468256 67732 468268
rect 67784 468256 67790 468308
rect 197262 468256 197268 468308
rect 197320 468296 197326 468308
rect 209774 468296 209780 468308
rect 197320 468268 209780 468296
rect 197320 468256 197326 468268
rect 209774 468256 209780 468268
rect 209832 468256 209838 468308
rect 133138 467780 133144 467832
rect 133196 467820 133202 467832
rect 178034 467820 178040 467832
rect 133196 467792 178040 467820
rect 133196 467780 133202 467792
rect 178034 467780 178040 467792
rect 178092 467780 178098 467832
rect 296622 467780 296628 467832
rect 296680 467820 296686 467832
rect 360562 467820 360568 467832
rect 296680 467792 360568 467820
rect 296680 467780 296686 467792
rect 360562 467780 360568 467792
rect 360620 467780 360626 467832
rect 160738 467712 160744 467764
rect 160796 467752 160802 467764
rect 179414 467752 179420 467764
rect 160796 467724 179420 467752
rect 160796 467712 160802 467724
rect 179414 467712 179420 467724
rect 179472 467712 179478 467764
rect 299290 467712 299296 467764
rect 299348 467752 299354 467764
rect 371234 467752 371240 467764
rect 299348 467724 371240 467752
rect 299348 467712 299354 467724
rect 371234 467712 371240 467724
rect 371292 467712 371298 467764
rect 288250 467644 288256 467696
rect 288308 467684 288314 467696
rect 375834 467684 375840 467696
rect 288308 467656 375840 467684
rect 288308 467644 288314 467656
rect 375834 467644 375840 467656
rect 375892 467644 375898 467696
rect 262306 467576 262312 467628
rect 262364 467616 262370 467628
rect 364058 467616 364064 467628
rect 262364 467588 364064 467616
rect 262364 467576 262370 467588
rect 364058 467576 364064 467588
rect 364116 467576 364122 467628
rect 42518 467508 42524 467560
rect 42576 467548 42582 467560
rect 61010 467548 61016 467560
rect 42576 467520 61016 467548
rect 42576 467508 42582 467520
rect 61010 467508 61016 467520
rect 61068 467508 61074 467560
rect 270678 467508 270684 467560
rect 270736 467548 270742 467560
rect 377122 467548 377128 467560
rect 270736 467520 377128 467548
rect 270736 467508 270742 467520
rect 377122 467508 377128 467520
rect 377180 467508 377186 467560
rect 40862 467440 40868 467492
rect 40920 467480 40926 467492
rect 62298 467480 62304 467492
rect 40920 467452 62304 467480
rect 40920 467440 40926 467452
rect 62298 467440 62304 467452
rect 62356 467440 62362 467492
rect 190086 467440 190092 467492
rect 190144 467480 190150 467492
rect 208026 467480 208032 467492
rect 190144 467452 208032 467480
rect 190144 467440 190150 467452
rect 208026 467440 208032 467452
rect 208084 467440 208090 467492
rect 252186 467440 252192 467492
rect 252244 467480 252250 467492
rect 361298 467480 361304 467492
rect 252244 467452 361304 467480
rect 252244 467440 252250 467452
rect 361298 467440 361304 467452
rect 361356 467440 361362 467492
rect 41138 467372 41144 467424
rect 41196 467412 41202 467424
rect 68278 467412 68284 467424
rect 41196 467384 68284 467412
rect 41196 467372 41202 467384
rect 68278 467372 68284 467384
rect 68336 467372 68342 467424
rect 185210 467372 185216 467424
rect 185268 467412 185274 467424
rect 212166 467412 212172 467424
rect 185268 467384 212172 467412
rect 185268 467372 185274 467384
rect 212166 467372 212172 467384
rect 212224 467372 212230 467424
rect 251726 467372 251732 467424
rect 251784 467412 251790 467424
rect 365346 467412 365352 467424
rect 251784 467384 365352 467412
rect 251784 467372 251790 467384
rect 365346 467372 365352 467384
rect 365404 467372 365410 467424
rect 41230 467304 41236 467356
rect 41288 467344 41294 467356
rect 72878 467344 72884 467356
rect 41288 467316 72884 467344
rect 41288 467304 41294 467316
rect 72878 467304 72884 467316
rect 72936 467304 72942 467356
rect 182174 467304 182180 467356
rect 182232 467344 182238 467356
rect 209590 467344 209596 467356
rect 182232 467316 209596 467344
rect 182232 467304 182238 467316
rect 209590 467304 209596 467316
rect 209648 467304 209654 467356
rect 249518 467304 249524 467356
rect 249576 467344 249582 467356
rect 367830 467344 367836 467356
rect 249576 467316 367836 467344
rect 249576 467304 249582 467316
rect 367830 467304 367836 467316
rect 367888 467304 367894 467356
rect 42702 467236 42708 467288
rect 42760 467276 42766 467288
rect 94958 467276 94964 467288
rect 42760 467248 94964 467276
rect 42760 467236 42766 467248
rect 94958 467236 94964 467248
rect 95016 467236 95022 467288
rect 188338 467236 188344 467288
rect 188396 467276 188402 467288
rect 216214 467276 216220 467288
rect 188396 467248 216220 467276
rect 188396 467236 188402 467248
rect 216214 467236 216220 467248
rect 216272 467236 216278 467288
rect 249978 467236 249984 467288
rect 250036 467276 250042 467288
rect 369302 467276 369308 467288
rect 250036 467248 369308 467276
rect 250036 467236 250042 467248
rect 369302 467236 369308 467248
rect 369360 467236 369366 467288
rect 57422 467168 57428 467220
rect 57480 467208 57486 467220
rect 112530 467208 112536 467220
rect 57480 467180 112536 467208
rect 57480 467168 57486 467180
rect 112530 467168 112536 467180
rect 112588 467168 112594 467220
rect 171594 467168 171600 467220
rect 171652 467208 171658 467220
rect 214742 467208 214748 467220
rect 171652 467180 214748 467208
rect 171652 467168 171658 467180
rect 214742 467168 214748 467180
rect 214800 467168 214806 467220
rect 250438 467168 250444 467220
rect 250496 467208 250502 467220
rect 371970 467208 371976 467220
rect 250496 467180 371976 467208
rect 250496 467168 250502 467180
rect 371970 467168 371976 467180
rect 372028 467168 372034 467220
rect 44910 467100 44916 467152
rect 44968 467140 44974 467152
rect 107286 467140 107292 467152
rect 44968 467112 107292 467140
rect 44968 467100 44974 467112
rect 107286 467100 107292 467112
rect 107344 467100 107350 467152
rect 165430 467100 165436 467152
rect 165488 467140 165494 467152
rect 218882 467140 218888 467152
rect 165488 467112 218888 467140
rect 165488 467100 165494 467112
rect 218882 467100 218888 467112
rect 218940 467100 218946 467152
rect 249058 467100 249064 467152
rect 249116 467140 249122 467152
rect 370774 467140 370780 467152
rect 249116 467112 370780 467140
rect 249116 467100 249122 467112
rect 370774 467100 370780 467112
rect 370832 467100 370838 467152
rect 59262 467032 59268 467084
rect 59320 467072 59326 467084
rect 67174 467072 67180 467084
rect 59320 467044 67180 467072
rect 59320 467032 59326 467044
rect 67174 467032 67180 467044
rect 67232 467032 67238 467084
rect 498470 466664 498476 466676
rect 489886 466636 498476 466664
rect 178034 466556 178040 466608
rect 178092 466596 178098 466608
rect 204530 466596 204536 466608
rect 178092 466568 204536 466596
rect 178092 466556 178098 466568
rect 204530 466556 204536 466568
rect 204588 466596 204594 466608
rect 338482 466596 338488 466608
rect 204588 466568 338488 466596
rect 204588 466556 204594 466568
rect 338482 466556 338488 466568
rect 338540 466596 338546 466608
rect 361574 466596 361580 466608
rect 338540 466568 361580 466596
rect 338540 466556 338546 466568
rect 361574 466556 361580 466568
rect 361632 466596 361638 466608
rect 489886 466596 489914 466636
rect 498470 466624 498476 466636
rect 498528 466664 498534 466676
rect 499482 466664 499488 466676
rect 498528 466636 499488 466664
rect 498528 466624 498534 466636
rect 499482 466624 499488 466636
rect 499540 466624 499546 466676
rect 499758 466596 499764 466608
rect 361632 466568 489914 466596
rect 496096 466568 499764 466596
rect 361632 466556 361638 466568
rect 179414 466488 179420 466540
rect 179472 466528 179478 466540
rect 201770 466528 201776 466540
rect 179472 466500 201776 466528
rect 179472 466488 179478 466500
rect 201770 466488 201776 466500
rect 201828 466528 201834 466540
rect 339770 466528 339776 466540
rect 201828 466500 339776 466528
rect 201828 466488 201834 466500
rect 339770 466488 339776 466500
rect 339828 466528 339834 466540
rect 362954 466528 362960 466540
rect 339828 466500 362960 466528
rect 339828 466488 339834 466500
rect 362954 466488 362960 466500
rect 363012 466528 363018 466540
rect 363012 466500 364334 466528
rect 363012 466488 363018 466500
rect 190914 466420 190920 466472
rect 190972 466460 190978 466472
rect 210418 466460 210424 466472
rect 190972 466432 210424 466460
rect 190972 466420 190978 466432
rect 210418 466420 210424 466432
rect 210476 466420 210482 466472
rect 350994 466420 351000 466472
rect 351052 466460 351058 466472
rect 358814 466460 358820 466472
rect 351052 466432 358820 466460
rect 351052 466420 351058 466432
rect 358814 466420 358820 466432
rect 358872 466420 358878 466472
rect 364306 466460 364334 466500
rect 496096 466460 496124 466568
rect 499758 466556 499764 466568
rect 499816 466596 499822 466608
rect 517882 466596 517888 466608
rect 499816 466568 517888 466596
rect 499816 466556 499822 466568
rect 517882 466556 517888 466568
rect 517940 466556 517946 466608
rect 499482 466488 499488 466540
rect 499540 466528 499546 466540
rect 499540 466500 509234 466528
rect 499540 466488 499546 466500
rect 364306 466432 496124 466460
rect 509206 466460 509234 466500
rect 510890 466488 510896 466540
rect 510948 466528 510954 466540
rect 517514 466528 517520 466540
rect 510948 466500 517520 466528
rect 510948 466488 510954 466500
rect 517514 466488 517520 466500
rect 517572 466488 517578 466540
rect 517790 466460 517796 466472
rect 509206 466432 517796 466460
rect 517790 466420 517796 466432
rect 517848 466420 517854 466472
rect 50706 466352 50712 466404
rect 50764 466392 50770 466404
rect 79502 466392 79508 466404
rect 50764 466364 79508 466392
rect 50764 466352 50770 466364
rect 79502 466352 79508 466364
rect 79560 466352 79566 466404
rect 194042 466352 194048 466404
rect 194100 466392 194106 466404
rect 212902 466392 212908 466404
rect 194100 466364 212908 466392
rect 194100 466352 194106 466364
rect 212902 466352 212908 466364
rect 212960 466352 212966 466404
rect 213822 466352 213828 466404
rect 213880 466392 213886 466404
rect 221366 466392 221372 466404
rect 213880 466364 221372 466392
rect 213880 466352 213886 466364
rect 221366 466352 221372 466364
rect 221424 466352 221430 466404
rect 280338 466352 280344 466404
rect 280396 466392 280402 466404
rect 368934 466392 368940 466404
rect 280396 466364 368940 466392
rect 280396 466352 280402 466364
rect 368934 466352 368940 466364
rect 368992 466352 368998 466404
rect 180334 466284 180340 466336
rect 180392 466324 180398 466336
rect 207842 466324 207848 466336
rect 180392 466296 207848 466324
rect 180392 466284 180398 466296
rect 207842 466284 207848 466296
rect 207900 466284 207906 466336
rect 275922 466284 275928 466336
rect 275980 466324 275986 466336
rect 372982 466324 372988 466336
rect 275980 466296 372988 466324
rect 275980 466284 275986 466296
rect 372982 466284 372988 466296
rect 373040 466284 373046 466336
rect 174170 466216 174176 466268
rect 174228 466256 174234 466268
rect 203886 466256 203892 466268
rect 174228 466228 203892 466256
rect 174228 466216 174234 466228
rect 203886 466216 203892 466228
rect 203944 466216 203950 466268
rect 263134 466216 263140 466268
rect 263192 466256 263198 466268
rect 369486 466256 369492 466268
rect 263192 466228 369492 466256
rect 263192 466216 263198 466228
rect 369486 466216 369492 466228
rect 369544 466216 369550 466268
rect 54386 466148 54392 466200
rect 54444 466188 54450 466200
rect 63218 466188 63224 466200
rect 54444 466160 63224 466188
rect 54444 466148 54450 466160
rect 63218 466148 63224 466160
rect 63276 466148 63282 466200
rect 168006 466148 168012 466200
rect 168064 466188 168070 466200
rect 203610 466188 203616 466200
rect 168064 466160 203616 466188
rect 168064 466148 168070 466160
rect 203610 466148 203616 466160
rect 203668 466148 203674 466200
rect 263594 466148 263600 466200
rect 263652 466188 263658 466200
rect 372154 466188 372160 466200
rect 263652 466160 372160 466188
rect 263652 466148 263658 466160
rect 372154 466148 372160 466160
rect 372212 466148 372218 466200
rect 59170 466080 59176 466132
rect 59228 466120 59234 466132
rect 67634 466120 67640 466132
rect 59228 466092 67640 466120
rect 59228 466080 59234 466092
rect 67634 466080 67640 466092
rect 67692 466080 67698 466132
rect 179506 466080 179512 466132
rect 179564 466120 179570 466132
rect 216306 466120 216312 466132
rect 179564 466092 216312 466120
rect 179564 466080 179570 466092
rect 216306 466080 216312 466092
rect 216364 466080 216370 466132
rect 257430 466080 257436 466132
rect 257488 466120 257494 466132
rect 366910 466120 366916 466132
rect 257488 466092 366916 466120
rect 257488 466080 257494 466092
rect 366910 466080 366916 466092
rect 366968 466080 366974 466132
rect 54294 466012 54300 466064
rect 54352 466052 54358 466064
rect 63678 466052 63684 466064
rect 54352 466024 63684 466052
rect 54352 466012 54358 466024
rect 63678 466012 63684 466024
rect 63736 466012 63742 466064
rect 166718 466012 166724 466064
rect 166776 466052 166782 466064
rect 206370 466052 206376 466064
rect 166776 466024 206376 466052
rect 166776 466012 166782 466024
rect 206370 466012 206376 466024
rect 206428 466012 206434 466064
rect 258350 466012 258356 466064
rect 258408 466052 258414 466064
rect 368106 466052 368112 466064
rect 258408 466024 368112 466052
rect 258408 466012 258414 466024
rect 368106 466012 368112 466024
rect 368164 466012 368170 466064
rect 51534 465944 51540 465996
rect 51592 465984 51598 465996
rect 66714 465984 66720 465996
rect 51592 465956 66720 465984
rect 51592 465944 51598 465956
rect 66714 465944 66720 465956
rect 66772 465944 66778 465996
rect 174630 465944 174636 465996
rect 174688 465984 174694 465996
rect 219158 465984 219164 465996
rect 174688 465956 219164 465984
rect 174688 465944 174694 465956
rect 219158 465944 219164 465956
rect 219216 465944 219222 465996
rect 243814 465944 243820 465996
rect 243872 465984 243878 465996
rect 358354 465984 358360 465996
rect 243872 465956 358360 465984
rect 243872 465944 243878 465956
rect 358354 465944 358360 465956
rect 358412 465944 358418 465996
rect 55582 465876 55588 465928
rect 55640 465916 55646 465928
rect 75546 465916 75552 465928
rect 55640 465888 75552 465916
rect 55640 465876 55646 465888
rect 75546 465876 75552 465888
rect 75604 465876 75610 465928
rect 164970 465876 164976 465928
rect 165028 465916 165034 465928
rect 214650 465916 214656 465928
rect 165028 465888 214656 465916
rect 165028 465876 165034 465888
rect 214650 465876 214656 465888
rect 214708 465876 214714 465928
rect 262766 465876 262772 465928
rect 262824 465916 262830 465928
rect 379054 465916 379060 465928
rect 262824 465888 379060 465916
rect 262824 465876 262830 465888
rect 379054 465876 379060 465888
rect 379112 465876 379118 465928
rect 49510 465808 49516 465860
rect 49568 465848 49574 465860
rect 71130 465848 71136 465860
rect 49568 465820 71136 465848
rect 49568 465808 49574 465820
rect 71130 465808 71136 465820
rect 71188 465808 71194 465860
rect 143350 465808 143356 465860
rect 143408 465848 143414 465860
rect 200482 465848 200488 465860
rect 143408 465820 200488 465848
rect 143408 465808 143414 465820
rect 200482 465808 200488 465820
rect 200540 465808 200546 465860
rect 244274 465808 244280 465860
rect 244332 465848 244338 465860
rect 373442 465848 373448 465860
rect 244332 465820 373448 465848
rect 244332 465808 244338 465820
rect 373442 465808 373448 465820
rect 373500 465808 373506 465860
rect 50798 465740 50804 465792
rect 50856 465780 50862 465792
rect 50982 465780 50988 465792
rect 50856 465752 50988 465780
rect 50856 465740 50862 465752
rect 50982 465740 50988 465752
rect 51040 465740 51046 465792
rect 93578 465780 93584 465792
rect 51184 465752 93584 465780
rect 50614 465672 50620 465724
rect 50672 465712 50678 465724
rect 51184 465712 51212 465752
rect 93578 465740 93584 465752
rect 93636 465740 93642 465792
rect 142522 465740 142528 465792
rect 142580 465780 142586 465792
rect 207106 465780 207112 465792
rect 142580 465752 207112 465780
rect 142580 465740 142586 465752
rect 207106 465740 207112 465752
rect 207164 465740 207170 465792
rect 212442 465740 212448 465792
rect 212500 465780 212506 465792
rect 221734 465780 221740 465792
rect 212500 465752 221740 465780
rect 212500 465740 212506 465752
rect 221734 465740 221740 465752
rect 221792 465740 221798 465792
rect 246390 465740 246396 465792
rect 246448 465780 246454 465792
rect 378962 465780 378968 465792
rect 246448 465752 378968 465780
rect 246448 465740 246454 465752
rect 378962 465740 378968 465752
rect 379020 465740 379026 465792
rect 71774 465712 71780 465724
rect 50672 465684 51212 465712
rect 55186 465684 71780 465712
rect 50672 465672 50678 465684
rect 49602 465604 49608 465656
rect 49660 465644 49666 465656
rect 55186 465644 55214 465684
rect 71774 465672 71780 465684
rect 71832 465672 71838 465724
rect 86218 465672 86224 465724
rect 86276 465712 86282 465724
rect 198734 465712 198740 465724
rect 86276 465684 198740 465712
rect 86276 465672 86282 465684
rect 198734 465672 198740 465684
rect 198792 465672 198798 465724
rect 205542 465672 205548 465724
rect 205600 465712 205606 465724
rect 220906 465712 220912 465724
rect 205600 465684 220912 465712
rect 205600 465672 205606 465684
rect 220906 465672 220912 465684
rect 220964 465672 220970 465724
rect 241146 465672 241152 465724
rect 241204 465712 241210 465724
rect 374914 465712 374920 465724
rect 241204 465684 374920 465712
rect 241204 465672 241210 465684
rect 374914 465672 374920 465684
rect 374972 465672 374978 465724
rect 49660 465616 55214 465644
rect 49660 465604 49666 465616
rect 59814 465604 59820 465656
rect 59872 465644 59878 465656
rect 62850 465644 62856 465656
rect 59872 465616 62856 465644
rect 59872 465604 59878 465616
rect 62850 465604 62856 465616
rect 62908 465604 62914 465656
rect 187878 465604 187884 465656
rect 187936 465644 187942 465656
rect 202506 465644 202512 465656
rect 187936 465616 202512 465644
rect 187936 465604 187942 465616
rect 202506 465604 202512 465616
rect 202564 465604 202570 465656
rect 274174 465604 274180 465656
rect 274232 465644 274238 465656
rect 362126 465644 362132 465656
rect 274232 465616 362132 465644
rect 274232 465604 274238 465616
rect 362126 465604 362132 465616
rect 362184 465604 362190 465656
rect 189166 465536 189172 465588
rect 189224 465576 189230 465588
rect 202138 465576 202144 465588
rect 189224 465548 202144 465576
rect 189224 465536 189230 465548
rect 202138 465536 202144 465548
rect 202196 465536 202202 465588
rect 297082 465536 297088 465588
rect 297140 465576 297146 465588
rect 362862 465576 362868 465588
rect 297140 465548 362868 465576
rect 297140 465536 297146 465548
rect 362862 465536 362868 465548
rect 362920 465536 362926 465588
rect 195790 465468 195796 465520
rect 195848 465508 195854 465520
rect 206738 465508 206744 465520
rect 195848 465480 206744 465508
rect 195848 465468 195854 465480
rect 206738 465468 206744 465480
rect 206796 465468 206802 465520
rect 198734 465060 198740 465112
rect 198792 465100 198798 465112
rect 358906 465100 358912 465112
rect 198792 465072 358912 465100
rect 198792 465060 198798 465072
rect 358906 465060 358912 465072
rect 358964 465100 358970 465112
rect 518894 465100 518900 465112
rect 358964 465072 518900 465100
rect 358964 465060 358970 465072
rect 518894 465060 518900 465072
rect 518952 465060 518958 465112
rect 196986 464992 196992 465044
rect 197044 465032 197050 465044
rect 200574 465032 200580 465044
rect 197044 465004 200580 465032
rect 197044 464992 197050 465004
rect 200574 464992 200580 465004
rect 200632 464992 200638 465044
rect 58986 464720 58992 464772
rect 59044 464760 59050 464772
rect 93210 464760 93216 464772
rect 59044 464732 93216 464760
rect 59044 464720 59050 464732
rect 93210 464720 93216 464732
rect 93268 464720 93274 464772
rect 192294 464720 192300 464772
rect 192352 464760 192358 464772
rect 208946 464760 208952 464772
rect 192352 464732 208952 464760
rect 192352 464720 192358 464732
rect 208946 464720 208952 464732
rect 209004 464720 209010 464772
rect 49970 464652 49976 464704
rect 50028 464692 50034 464704
rect 50706 464692 50712 464704
rect 50028 464664 50712 464692
rect 50028 464652 50034 464664
rect 50706 464652 50712 464664
rect 50764 464652 50770 464704
rect 53006 464652 53012 464704
rect 53064 464692 53070 464704
rect 101950 464692 101956 464704
rect 53064 464664 101956 464692
rect 53064 464652 53070 464664
rect 101950 464652 101956 464664
rect 102008 464652 102014 464704
rect 191834 464652 191840 464704
rect 191892 464692 191898 464704
rect 211614 464692 211620 464704
rect 191892 464664 211620 464692
rect 191892 464652 191898 464664
rect 211614 464652 211620 464664
rect 211672 464652 211678 464704
rect 55766 464584 55772 464636
rect 55824 464624 55830 464636
rect 122650 464624 122656 464636
rect 55824 464596 122656 464624
rect 55824 464584 55830 464596
rect 122650 464584 122656 464596
rect 122708 464584 122714 464636
rect 194502 464584 194508 464636
rect 194560 464624 194566 464636
rect 214466 464624 214472 464636
rect 194560 464596 214472 464624
rect 194560 464584 194566 464596
rect 214466 464584 214472 464596
rect 214524 464584 214530 464636
rect 54570 464516 54576 464568
rect 54628 464556 54634 464568
rect 121822 464556 121828 464568
rect 54628 464528 121828 464556
rect 54628 464516 54634 464528
rect 121822 464516 121828 464528
rect 121880 464516 121886 464568
rect 180794 464516 180800 464568
rect 180852 464556 180858 464568
rect 210878 464556 210884 464568
rect 180852 464528 210884 464556
rect 180852 464516 180858 464528
rect 210878 464516 210884 464528
rect 210936 464516 210942 464568
rect 57054 464448 57060 464500
rect 57112 464488 57118 464500
rect 134978 464488 134984 464500
rect 57112 464460 134984 464488
rect 57112 464448 57118 464460
rect 134978 464448 134984 464460
rect 135036 464448 135042 464500
rect 142890 464448 142896 464500
rect 142948 464488 142954 464500
rect 197814 464488 197820 464500
rect 142948 464460 197820 464488
rect 142948 464448 142954 464460
rect 197814 464448 197820 464460
rect 197872 464448 197878 464500
rect 207382 464488 207388 464500
rect 200086 464460 207388 464488
rect 52178 464380 52184 464432
rect 52236 464420 52242 464432
rect 134150 464420 134156 464432
rect 52236 464392 134156 464420
rect 52236 464380 52242 464392
rect 134150 464380 134156 464392
rect 134208 464380 134214 464432
rect 137186 464380 137192 464432
rect 137244 464420 137250 464432
rect 199010 464420 199016 464432
rect 137244 464392 199016 464420
rect 137244 464380 137250 464392
rect 199010 464380 199016 464392
rect 199068 464380 199074 464432
rect 47578 464312 47584 464364
rect 47636 464352 47642 464364
rect 200086 464352 200114 464460
rect 207382 464448 207388 464460
rect 207440 464488 207446 464500
rect 208210 464488 208216 464500
rect 207440 464460 208216 464488
rect 207440 464448 207446 464460
rect 208210 464448 208216 464460
rect 208268 464448 208274 464500
rect 294414 464448 294420 464500
rect 294472 464488 294478 464500
rect 370222 464488 370228 464500
rect 294472 464460 370228 464488
rect 294472 464448 294478 464460
rect 370222 464448 370228 464460
rect 370280 464448 370286 464500
rect 288710 464380 288716 464432
rect 288768 464420 288774 464432
rect 367462 464420 367468 464432
rect 288768 464392 367468 464420
rect 288768 464380 288774 464392
rect 367462 464380 367468 464392
rect 367520 464380 367526 464432
rect 47636 464324 200114 464352
rect 47636 464312 47642 464324
rect 207474 464312 207480 464364
rect 207532 464352 207538 464364
rect 208118 464352 208124 464364
rect 207532 464324 208124 464352
rect 207532 464312 207538 464324
rect 208118 464312 208124 464324
rect 208176 464312 208182 464364
rect 276842 464312 276848 464364
rect 276900 464352 276906 464364
rect 357894 464352 357900 464364
rect 276900 464324 357900 464352
rect 276900 464312 276906 464324
rect 357894 464312 357900 464324
rect 357952 464312 357958 464364
rect 46014 464244 46020 464296
rect 46072 464284 46078 464296
rect 207492 464284 207520 464312
rect 46072 464256 207520 464284
rect 46072 464244 46078 464256
rect 208210 418752 208216 418804
rect 208268 418792 208274 418804
rect 216858 418792 216864 418804
rect 208268 418764 216864 418792
rect 208268 418752 208274 418764
rect 216858 418752 216864 418764
rect 216916 418752 216922 418804
rect 46014 418072 46020 418124
rect 46072 418112 46078 418124
rect 57790 418112 57796 418124
rect 46072 418084 57796 418112
rect 46072 418072 46078 418084
rect 57790 418072 57796 418084
rect 57848 418072 57854 418124
rect 47578 418004 47584 418056
rect 47636 418044 47642 418056
rect 57238 418044 57244 418056
rect 47636 418016 57244 418044
rect 47636 418004 47642 418016
rect 57238 418004 57244 418016
rect 57296 418004 57302 418056
rect 203058 418004 203064 418056
rect 203116 418044 203122 418056
rect 208210 418044 208216 418056
rect 203116 418016 208216 418044
rect 203116 418004 203122 418016
rect 208210 418004 208216 418016
rect 208268 418004 208274 418056
rect 208118 417392 208124 417444
rect 208176 417432 208182 417444
rect 216766 417432 216772 417444
rect 208176 417404 216772 417432
rect 208176 417392 208182 417404
rect 216766 417392 216772 417404
rect 216824 417392 216830 417444
rect 358078 417392 358084 417444
rect 358136 417432 358142 417444
rect 377030 417432 377036 417444
rect 358136 417404 377036 417432
rect 358136 417392 358142 417404
rect 377030 417392 377036 417404
rect 377088 417432 377094 417444
rect 377582 417432 377588 417444
rect 377088 417404 377588 417432
rect 377088 417392 377094 417404
rect 377582 417392 377588 417404
rect 377640 417392 377646 417444
rect 206830 416712 206836 416764
rect 206888 416752 206894 416764
rect 207198 416752 207204 416764
rect 206888 416724 207204 416752
rect 206888 416712 206894 416724
rect 207198 416712 207204 416724
rect 207256 416712 207262 416764
rect 198182 416032 198188 416084
rect 198240 416072 198246 416084
rect 203058 416072 203064 416084
rect 198240 416044 203064 416072
rect 198240 416032 198246 416044
rect 203058 416032 203064 416044
rect 203116 416032 203122 416084
rect 207198 414808 207204 414860
rect 207256 414848 207262 414860
rect 216858 414848 216864 414860
rect 207256 414820 216864 414848
rect 207256 414808 207262 414820
rect 216858 414808 216864 414820
rect 216916 414808 216922 414860
rect 206186 414672 206192 414724
rect 206244 414712 206250 414724
rect 216950 414712 216956 414724
rect 206244 414684 216956 414712
rect 206244 414672 206250 414684
rect 216950 414672 216956 414684
rect 217008 414672 217014 414724
rect 47486 413992 47492 414044
rect 47544 414032 47550 414044
rect 57790 414032 57796 414044
rect 47544 414004 57796 414032
rect 47544 413992 47550 414004
rect 57790 413992 57796 414004
rect 57848 413992 57854 414044
rect 206002 413244 206008 413296
rect 206060 413284 206066 413296
rect 216674 413284 216680 413296
rect 206060 413256 216680 413284
rect 206060 413244 206066 413256
rect 216674 413244 216680 413256
rect 216732 413244 216738 413296
rect 359826 413244 359832 413296
rect 359884 413284 359890 413296
rect 377674 413284 377680 413296
rect 359884 413256 377680 413284
rect 359884 413244 359890 413256
rect 377674 413244 377680 413256
rect 377732 413244 377738 413296
rect 47394 412632 47400 412684
rect 47452 412672 47458 412684
rect 57790 412672 57796 412684
rect 47452 412644 57796 412672
rect 47452 412632 47458 412644
rect 57790 412632 57796 412644
rect 57848 412632 57854 412684
rect 359734 411884 359740 411936
rect 359792 411924 359798 411936
rect 377030 411924 377036 411936
rect 359792 411896 377036 411924
rect 359792 411884 359798 411896
rect 377030 411884 377036 411896
rect 377088 411884 377094 411936
rect 204438 411476 204444 411528
rect 204496 411516 204502 411528
rect 206830 411516 206836 411528
rect 204496 411488 206836 411516
rect 204496 411476 204502 411488
rect 206830 411476 206836 411488
rect 206888 411476 206894 411528
rect 47578 411272 47584 411324
rect 47636 411312 47642 411324
rect 57790 411312 57796 411324
rect 47636 411284 57796 411312
rect 47636 411272 47642 411284
rect 57790 411272 57796 411284
rect 57848 411272 57854 411324
rect 2958 411204 2964 411256
rect 3016 411244 3022 411256
rect 15838 411244 15844 411256
rect 3016 411216 15844 411244
rect 3016 411204 3022 411216
rect 15838 411204 15844 411216
rect 15896 411204 15902 411256
rect 51626 410592 51632 410644
rect 51684 410632 51690 410644
rect 52914 410632 52920 410644
rect 51684 410604 52920 410632
rect 51684 410592 51690 410604
rect 52914 410592 52920 410604
rect 52972 410592 52978 410644
rect 198090 410524 198096 410576
rect 198148 410564 198154 410576
rect 204438 410564 204444 410576
rect 198148 410536 204444 410564
rect 198148 410524 198154 410536
rect 204438 410524 204444 410536
rect 204496 410524 204502 410576
rect 360010 410524 360016 410576
rect 360068 410564 360074 410576
rect 377398 410564 377404 410576
rect 360068 410536 377404 410564
rect 360068 410524 360074 410536
rect 377398 410524 377404 410536
rect 377456 410564 377462 410576
rect 377858 410564 377864 410576
rect 377456 410536 377864 410564
rect 377456 410524 377462 410536
rect 377858 410524 377864 410536
rect 377916 410524 377922 410576
rect 51626 409844 51632 409896
rect 51684 409884 51690 409896
rect 57790 409884 57796 409896
rect 51684 409856 57796 409884
rect 51684 409844 51690 409856
rect 57790 409844 57796 409856
rect 57848 409844 57854 409896
rect 217962 409844 217968 409896
rect 218020 409884 218026 409896
rect 218606 409884 218612 409896
rect 218020 409856 218612 409884
rect 218020 409844 218026 409856
rect 218606 409844 218612 409856
rect 218664 409844 218670 409896
rect 206830 409096 206836 409148
rect 206888 409136 206894 409148
rect 216766 409136 216772 409148
rect 206888 409108 216772 409136
rect 206888 409096 206894 409108
rect 216766 409096 216772 409108
rect 216824 409136 216830 409148
rect 216950 409136 216956 409148
rect 216824 409108 216956 409136
rect 216824 409096 216830 409108
rect 216950 409096 216956 409108
rect 217008 409096 217014 409148
rect 359918 409096 359924 409148
rect 359976 409136 359982 409148
rect 377398 409136 377404 409148
rect 359976 409108 377404 409136
rect 359976 409096 359982 409108
rect 377398 409096 377404 409108
rect 377456 409096 377462 409148
rect 52362 408484 52368 408536
rect 52420 408524 52426 408536
rect 57790 408524 57796 408536
rect 52420 408496 57796 408524
rect 52420 408484 52426 408496
rect 57790 408484 57796 408496
rect 57848 408484 57854 408536
rect 216674 407600 216680 407652
rect 216732 407640 216738 407652
rect 216732 407612 216812 407640
rect 216732 407600 216738 407612
rect 216784 407448 216812 407612
rect 216766 407396 216772 407448
rect 216824 407396 216830 407448
rect 520918 405628 520924 405680
rect 520976 405668 520982 405680
rect 580166 405668 580172 405680
rect 520976 405640 580172 405668
rect 520976 405628 520982 405640
rect 580166 405628 580172 405640
rect 580224 405628 580230 405680
rect 199010 400528 199016 400580
rect 199068 400528 199074 400580
rect 199102 400528 199108 400580
rect 199160 400568 199166 400580
rect 199838 400568 199844 400580
rect 199160 400540 199844 400568
rect 199160 400528 199166 400540
rect 199838 400528 199844 400540
rect 199896 400528 199902 400580
rect 199028 400376 199056 400528
rect 199010 400324 199016 400376
rect 199068 400324 199074 400376
rect 198918 400188 198924 400240
rect 198976 400228 198982 400240
rect 208486 400228 208492 400240
rect 198976 400200 208492 400228
rect 198976 400188 198982 400200
rect 208486 400188 208492 400200
rect 208544 400188 208550 400240
rect 378134 398080 378140 398132
rect 378192 398120 378198 398132
rect 378318 398120 378324 398132
rect 378192 398092 378324 398120
rect 378192 398080 378198 398092
rect 378318 398080 378324 398092
rect 378376 398080 378382 398132
rect 198090 397400 198096 397452
rect 198148 397440 198154 397452
rect 199102 397440 199108 397452
rect 198148 397412 199108 397440
rect 198148 397400 198154 397412
rect 199102 397400 199108 397412
rect 199160 397400 199166 397452
rect 56502 391960 56508 392012
rect 56560 392000 56566 392012
rect 57054 392000 57060 392012
rect 56560 391972 57060 392000
rect 56560 391960 56566 391972
rect 57054 391960 57060 391972
rect 57112 391960 57118 392012
rect 43254 391892 43260 391944
rect 43312 391932 43318 391944
rect 57698 391932 57704 391944
rect 43312 391904 57704 391932
rect 43312 391892 43318 391904
rect 57698 391892 57704 391904
rect 57756 391892 57762 391944
rect 208210 391892 208216 391944
rect 208268 391932 208274 391944
rect 216950 391932 216956 391944
rect 208268 391904 216956 391932
rect 208268 391892 208274 391904
rect 216950 391892 216956 391904
rect 217008 391892 217014 391944
rect 359642 391892 359648 391944
rect 359700 391932 359706 391944
rect 376846 391932 376852 391944
rect 359700 391904 376852 391932
rect 359700 391892 359706 391904
rect 376846 391892 376852 391904
rect 376904 391892 376910 391944
rect 57146 390532 57152 390584
rect 57204 390572 57210 390584
rect 58434 390572 58440 390584
rect 57204 390544 58440 390572
rect 57204 390532 57210 390544
rect 58434 390532 58440 390544
rect 58492 390532 58498 390584
rect 358814 390464 358820 390516
rect 358872 390504 358878 390516
rect 376938 390504 376944 390516
rect 358872 390476 376944 390504
rect 358872 390464 358878 390476
rect 376938 390464 376944 390476
rect 376996 390464 377002 390516
rect 210418 389308 210424 389360
rect 210476 389348 210482 389360
rect 216674 389348 216680 389360
rect 210476 389320 216680 389348
rect 210476 389308 210482 389320
rect 216674 389308 216680 389320
rect 216732 389308 216738 389360
rect 52454 389172 52460 389224
rect 52512 389212 52518 389224
rect 53742 389212 53748 389224
rect 52512 389184 53748 389212
rect 52512 389172 52518 389184
rect 53742 389172 53748 389184
rect 53800 389212 53806 389224
rect 57422 389212 57428 389224
rect 53800 389184 57428 389212
rect 53800 389172 53806 389184
rect 57422 389172 57428 389184
rect 57480 389172 57486 389224
rect 358078 389172 358084 389224
rect 358136 389212 358142 389224
rect 358814 389212 358820 389224
rect 358136 389184 358820 389212
rect 358136 389172 358142 389184
rect 358814 389172 358820 389184
rect 358872 389172 358878 389224
rect 47762 389104 47768 389156
rect 47820 389144 47826 389156
rect 57238 389144 57244 389156
rect 47820 389116 57244 389144
rect 47820 389104 47826 389116
rect 57238 389104 57244 389116
rect 57296 389104 57302 389156
rect 202138 389104 202144 389156
rect 202196 389144 202202 389156
rect 216950 389144 216956 389156
rect 202196 389116 216956 389144
rect 202196 389104 202202 389116
rect 216950 389104 216956 389116
rect 217008 389104 217014 389156
rect 359550 389104 359556 389156
rect 359608 389144 359614 389156
rect 376938 389144 376944 389156
rect 359608 389116 376944 389144
rect 359608 389104 359614 389116
rect 376938 389104 376944 389116
rect 376996 389104 377002 389156
rect 56778 388492 56784 388544
rect 56836 388532 56842 388544
rect 58526 388532 58532 388544
rect 56836 388504 58532 388532
rect 56836 388492 56842 388504
rect 58526 388492 58532 388504
rect 58584 388492 58590 388544
rect 45462 388424 45468 388476
rect 45520 388464 45526 388476
rect 52454 388464 52460 388476
rect 45520 388436 52460 388464
rect 45520 388424 45526 388436
rect 52454 388424 52460 388436
rect 52512 388424 52518 388476
rect 57054 388424 57060 388476
rect 57112 388464 57118 388476
rect 58434 388464 58440 388476
rect 57112 388436 58440 388464
rect 57112 388424 57118 388436
rect 58434 388424 58440 388436
rect 58492 388424 58498 388476
rect 57146 387948 57152 388000
rect 57204 387988 57210 388000
rect 57790 387988 57796 388000
rect 57204 387960 57796 387988
rect 57204 387948 57210 387960
rect 57790 387948 57796 387960
rect 57848 387948 57854 388000
rect 378134 383936 378140 383988
rect 378192 383976 378198 383988
rect 378318 383976 378324 383988
rect 378192 383948 378324 383976
rect 378192 383936 378198 383948
rect 378318 383936 378324 383948
rect 378376 383936 378382 383988
rect 199286 382916 199292 382968
rect 199344 382956 199350 382968
rect 219802 382956 219808 382968
rect 199344 382928 219808 382956
rect 199344 382916 199350 382928
rect 219802 382916 219808 382928
rect 219860 382916 219866 382968
rect 57790 382032 57796 382084
rect 57848 382072 57854 382084
rect 59354 382072 59360 382084
rect 57848 382044 59360 382072
rect 57848 382032 57854 382044
rect 59354 382032 59360 382044
rect 59412 382032 59418 382084
rect 195054 380944 195060 380996
rect 195112 380984 195118 380996
rect 200574 380984 200580 380996
rect 195112 380956 200580 380984
rect 195112 380944 195118 380956
rect 200574 380944 200580 380956
rect 200632 380944 200638 380996
rect 55766 380876 55772 380928
rect 55824 380916 55830 380928
rect 57054 380916 57060 380928
rect 55824 380888 57060 380916
rect 55824 380876 55830 380888
rect 57054 380876 57060 380888
rect 57112 380876 57118 380928
rect 58342 380876 58348 380928
rect 58400 380916 58406 380928
rect 60734 380916 60740 380928
rect 58400 380888 60740 380916
rect 58400 380876 58406 380888
rect 60734 380876 60740 380888
rect 60792 380876 60798 380928
rect 194594 380876 194600 380928
rect 194652 380916 194658 380928
rect 197722 380916 197728 380928
rect 194652 380888 197728 380916
rect 194652 380876 194658 380888
rect 197722 380876 197728 380888
rect 197780 380876 197786 380928
rect 217594 380876 217600 380928
rect 217652 380916 217658 380928
rect 248230 380916 248236 380928
rect 217652 380888 248236 380916
rect 217652 380876 217658 380888
rect 248230 380876 248236 380888
rect 248288 380876 248294 380928
rect 358722 380876 358728 380928
rect 358780 380916 358786 380928
rect 421098 380916 421104 380928
rect 358780 380888 421104 380916
rect 358780 380876 358786 380888
rect 421098 380876 421104 380888
rect 421156 380876 421162 380928
rect 47394 380808 47400 380860
rect 47452 380848 47458 380860
rect 216766 380848 216772 380860
rect 47452 380820 216772 380848
rect 47452 380808 47458 380820
rect 216766 380808 216772 380820
rect 216824 380808 216830 380860
rect 47486 380740 47492 380792
rect 47544 380780 47550 380792
rect 216674 380780 216680 380792
rect 47544 380752 216680 380780
rect 47544 380740 47550 380752
rect 216674 380740 216680 380752
rect 216732 380740 216738 380792
rect 356974 380740 356980 380792
rect 357032 380780 357038 380792
rect 380986 380780 380992 380792
rect 357032 380752 380992 380780
rect 357032 380740 357038 380752
rect 380986 380740 380992 380752
rect 381044 380740 381050 380792
rect 51626 380672 51632 380724
rect 51684 380712 51690 380724
rect 217134 380712 217140 380724
rect 51684 380684 217140 380712
rect 51684 380672 51690 380684
rect 217134 380672 217140 380684
rect 217192 380672 217198 380724
rect 377306 380672 377312 380724
rect 377364 380712 377370 380724
rect 413554 380712 413560 380724
rect 377364 380684 413560 380712
rect 377364 380672 377370 380684
rect 413554 380672 413560 380684
rect 413612 380672 413618 380724
rect 52362 380604 52368 380656
rect 52420 380644 52426 380656
rect 216858 380644 216864 380656
rect 52420 380616 216864 380644
rect 52420 380604 52426 380616
rect 216858 380604 216864 380616
rect 216916 380604 216922 380656
rect 357986 380604 357992 380656
rect 358044 380644 358050 380656
rect 376478 380644 376484 380656
rect 358044 380616 376484 380644
rect 358044 380604 358050 380616
rect 376478 380604 376484 380616
rect 376536 380604 376542 380656
rect 377122 380604 377128 380656
rect 377180 380644 377186 380656
rect 425974 380644 425980 380656
rect 377180 380616 425980 380644
rect 377180 380604 377186 380616
rect 425974 380604 425980 380616
rect 426032 380604 426038 380656
rect 155954 380536 155960 380588
rect 156012 380576 156018 380588
rect 204622 380576 204628 380588
rect 156012 380548 204628 380576
rect 156012 380536 156018 380548
rect 204622 380536 204628 380548
rect 204680 380536 204686 380588
rect 360562 380536 360568 380588
rect 360620 380576 360626 380588
rect 369578 380576 369584 380588
rect 360620 380548 369584 380576
rect 360620 380536 360626 380548
rect 369578 380536 369584 380548
rect 369636 380536 369642 380588
rect 372246 380536 372252 380588
rect 372304 380576 372310 380588
rect 433610 380576 433616 380588
rect 372304 380548 433616 380576
rect 372304 380536 372310 380548
rect 433610 380536 433616 380548
rect 433668 380536 433674 380588
rect 143626 380468 143632 380520
rect 143684 380508 143690 380520
rect 205726 380508 205732 380520
rect 143684 380480 205732 380508
rect 143684 380468 143690 380480
rect 205726 380468 205732 380480
rect 205784 380468 205790 380520
rect 368842 380468 368848 380520
rect 368900 380508 368906 380520
rect 436002 380508 436008 380520
rect 368900 380480 436008 380508
rect 368900 380468 368906 380480
rect 436002 380468 436008 380480
rect 436060 380468 436066 380520
rect 56502 380400 56508 380452
rect 56560 380440 56566 380452
rect 118326 380440 118332 380452
rect 56560 380412 118332 380440
rect 56560 380400 56566 380412
rect 118326 380400 118332 380412
rect 118384 380400 118390 380452
rect 120994 380400 121000 380452
rect 121052 380440 121058 380452
rect 203058 380440 203064 380452
rect 121052 380412 203064 380440
rect 121052 380400 121058 380412
rect 203058 380400 203064 380412
rect 203116 380400 203122 380452
rect 366266 380400 366272 380452
rect 366324 380440 366330 380452
rect 438486 380440 438492 380452
rect 366324 380412 438492 380440
rect 366324 380400 366330 380412
rect 438486 380400 438492 380412
rect 438544 380400 438550 380452
rect 52178 380332 52184 380384
rect 52236 380372 52242 380384
rect 113542 380372 113548 380384
rect 52236 380344 113548 380372
rect 52236 380332 52242 380344
rect 113542 380332 113548 380344
rect 113600 380332 113606 380384
rect 163498 380332 163504 380384
rect 163556 380372 163562 380384
rect 197814 380372 197820 380384
rect 163556 380344 197820 380372
rect 163556 380332 163562 380344
rect 197814 380332 197820 380344
rect 197872 380332 197878 380384
rect 201586 380332 201592 380384
rect 201644 380372 201650 380384
rect 291838 380372 291844 380384
rect 201644 380344 291844 380372
rect 201644 380332 201650 380344
rect 291838 380332 291844 380344
rect 291896 380332 291902 380384
rect 364242 380332 364248 380384
rect 364300 380372 364306 380384
rect 440878 380372 440884 380384
rect 364300 380344 440884 380372
rect 364300 380332 364306 380344
rect 440878 380332 440884 380344
rect 440936 380332 440942 380384
rect 48774 380264 48780 380316
rect 48832 380304 48838 380316
rect 110966 380304 110972 380316
rect 48832 380276 110972 380304
rect 48832 380264 48838 380276
rect 110966 380264 110972 380276
rect 111024 380264 111030 380316
rect 148594 380264 148600 380316
rect 148652 380304 148658 380316
rect 196894 380304 196900 380316
rect 148652 380276 196900 380304
rect 148652 380264 148658 380276
rect 196894 380264 196900 380276
rect 196952 380264 196958 380316
rect 199746 380264 199752 380316
rect 199804 380304 199810 380316
rect 298002 380304 298008 380316
rect 199804 380276 298008 380304
rect 199804 380264 199810 380276
rect 298002 380264 298008 380276
rect 298060 380264 298066 380316
rect 364886 380264 364892 380316
rect 364944 380304 364950 380316
rect 448238 380304 448244 380316
rect 364944 380276 448244 380304
rect 364944 380264 364950 380276
rect 448238 380264 448244 380276
rect 448296 380264 448302 380316
rect 57882 380196 57888 380248
rect 57940 380236 57946 380248
rect 123478 380236 123484 380248
rect 57940 380208 123484 380236
rect 57940 380196 57946 380208
rect 123478 380196 123484 380208
rect 123536 380196 123542 380248
rect 135898 380196 135904 380248
rect 135956 380236 135962 380248
rect 200298 380236 200304 380248
rect 135956 380208 200304 380236
rect 135956 380196 135962 380208
rect 200298 380196 200304 380208
rect 200356 380196 200362 380248
rect 201034 380196 201040 380248
rect 201092 380236 201098 380248
rect 313458 380236 313464 380248
rect 201092 380208 313464 380236
rect 201092 380196 201098 380208
rect 313458 380196 313464 380208
rect 313516 380196 313522 380248
rect 360654 380196 360660 380248
rect 360712 380236 360718 380248
rect 443454 380236 443460 380248
rect 360712 380208 443460 380236
rect 360712 380196 360718 380208
rect 443454 380196 443460 380208
rect 443512 380196 443518 380248
rect 48866 380128 48872 380180
rect 48924 380168 48930 380180
rect 115934 380168 115940 380180
rect 48924 380140 115940 380168
rect 48924 380128 48930 380140
rect 115934 380128 115940 380140
rect 115992 380128 115998 380180
rect 128354 380128 128360 380180
rect 128412 380168 128418 380180
rect 197630 380168 197636 380180
rect 128412 380140 197636 380168
rect 128412 380128 128418 380140
rect 197630 380128 197636 380140
rect 197688 380128 197694 380180
rect 201494 380128 201500 380180
rect 201552 380168 201558 380180
rect 315850 380168 315856 380180
rect 201552 380140 315856 380168
rect 201552 380128 201558 380140
rect 315850 380128 315856 380140
rect 315908 380128 315914 380180
rect 362126 380128 362132 380180
rect 362184 380168 362190 380180
rect 445938 380168 445944 380180
rect 362184 380140 445944 380168
rect 362184 380128 362190 380140
rect 445938 380128 445944 380140
rect 445996 380128 446002 380180
rect 158530 380060 158536 380112
rect 158588 380100 158594 380112
rect 205818 380100 205824 380112
rect 158588 380072 205824 380100
rect 158588 380060 158594 380072
rect 205818 380060 205824 380072
rect 205876 380060 205882 380112
rect 160922 379992 160928 380044
rect 160980 380032 160986 380044
rect 207106 380032 207112 380044
rect 160980 380004 207112 380032
rect 160980 379992 160986 380004
rect 207106 379992 207112 380004
rect 207164 379992 207170 380044
rect 213730 379992 213736 380044
rect 213788 380032 213794 380044
rect 235994 380032 236000 380044
rect 213788 380004 236000 380032
rect 213788 379992 213794 380004
rect 235994 379992 236000 380004
rect 236052 379992 236058 380044
rect 166074 379924 166080 379976
rect 166132 379964 166138 379976
rect 200482 379964 200488 379976
rect 166132 379936 200488 379964
rect 166132 379924 166138 379936
rect 200482 379924 200488 379936
rect 200540 379924 200546 379976
rect 215294 379924 215300 379976
rect 215352 379964 215358 379976
rect 216398 379964 216404 379976
rect 215352 379936 216404 379964
rect 215352 379924 215358 379936
rect 216398 379924 216404 379936
rect 216456 379964 216462 379976
rect 243078 379964 243084 379976
rect 216456 379936 243084 379964
rect 216456 379924 216462 379936
rect 243078 379924 243084 379936
rect 243136 379924 243142 379976
rect 208302 379856 208308 379908
rect 208360 379896 208366 379908
rect 237098 379896 237104 379908
rect 208360 379868 237104 379896
rect 208360 379856 208366 379868
rect 237098 379856 237104 379868
rect 237156 379856 237162 379908
rect 239766 379856 239772 379908
rect 239824 379896 239830 379908
rect 261754 379896 261760 379908
rect 239824 379868 261760 379896
rect 239824 379856 239830 379868
rect 261754 379856 261760 379868
rect 261812 379856 261818 379908
rect 213638 379788 213644 379840
rect 213696 379828 213702 379840
rect 214098 379828 214104 379840
rect 213696 379800 214104 379828
rect 213696 379788 213702 379800
rect 214098 379788 214104 379800
rect 214156 379828 214162 379840
rect 244274 379828 244280 379840
rect 214156 379800 244280 379828
rect 214156 379788 214162 379800
rect 244274 379788 244280 379800
rect 244332 379788 244338 379840
rect 375282 379788 375288 379840
rect 375340 379828 375346 379840
rect 405458 379828 405464 379840
rect 375340 379800 405464 379828
rect 375340 379788 375346 379800
rect 405458 379788 405464 379800
rect 405516 379788 405522 379840
rect 212626 379720 212632 379772
rect 212684 379760 212690 379772
rect 219710 379760 219716 379772
rect 212684 379732 219716 379760
rect 212684 379720 212690 379732
rect 219710 379720 219716 379732
rect 219768 379760 219774 379772
rect 254486 379760 254492 379772
rect 219768 379732 254492 379760
rect 219768 379720 219774 379732
rect 254486 379720 254492 379732
rect 254544 379720 254550 379772
rect 380986 379720 380992 379772
rect 381044 379760 381050 379772
rect 413462 379760 413468 379772
rect 381044 379732 413468 379760
rect 381044 379720 381050 379732
rect 413462 379720 413468 379732
rect 413520 379720 413526 379772
rect 215662 379652 215668 379704
rect 215720 379692 215726 379704
rect 216030 379692 216036 379704
rect 215720 379664 216036 379692
rect 215720 379652 215726 379664
rect 216030 379652 216036 379664
rect 216088 379692 216094 379704
rect 217318 379692 217324 379704
rect 216088 379664 217324 379692
rect 216088 379652 216094 379664
rect 217318 379652 217324 379664
rect 217376 379692 217382 379704
rect 217376 379664 217732 379692
rect 217376 379652 217382 379664
rect 216674 379584 216680 379636
rect 216732 379624 216738 379636
rect 217594 379624 217600 379636
rect 216732 379596 217600 379624
rect 216732 379584 216738 379596
rect 217594 379584 217600 379596
rect 217652 379584 217658 379636
rect 204162 379516 204168 379568
rect 204220 379556 204226 379568
rect 213730 379556 213736 379568
rect 204220 379528 213736 379556
rect 204220 379516 204226 379528
rect 213730 379516 213736 379528
rect 213788 379516 213794 379568
rect 216858 379516 216864 379568
rect 216916 379556 216922 379568
rect 217318 379556 217324 379568
rect 216916 379528 217324 379556
rect 216916 379516 216922 379528
rect 217318 379516 217324 379528
rect 217376 379516 217382 379568
rect 217704 379556 217732 379664
rect 217962 379652 217968 379704
rect 218020 379692 218026 379704
rect 255866 379692 255872 379704
rect 218020 379664 255872 379692
rect 218020 379652 218026 379664
rect 255866 379652 255872 379664
rect 255924 379652 255930 379704
rect 369762 379652 369768 379704
rect 369820 379692 369826 379704
rect 371142 379692 371148 379704
rect 369820 379664 371148 379692
rect 369820 379652 369826 379664
rect 371142 379652 371148 379664
rect 371200 379692 371206 379704
rect 404170 379692 404176 379704
rect 371200 379664 404176 379692
rect 371200 379652 371206 379664
rect 404170 379652 404176 379664
rect 404228 379652 404234 379704
rect 219250 379584 219256 379636
rect 219308 379624 219314 379636
rect 219434 379624 219440 379636
rect 219308 379596 219440 379624
rect 219308 379584 219314 379596
rect 219434 379584 219440 379596
rect 219492 379624 219498 379636
rect 258074 379624 258080 379636
rect 219492 379596 258080 379624
rect 219492 379584 219498 379596
rect 258074 379584 258080 379596
rect 258132 379584 258138 379636
rect 369578 379584 369584 379636
rect 369636 379624 369642 379636
rect 369636 379596 373994 379624
rect 369636 379584 369642 379596
rect 263870 379556 263876 379568
rect 217704 379528 263876 379556
rect 263870 379516 263876 379528
rect 263928 379516 263934 379568
rect 54478 379448 54484 379500
rect 54536 379488 54542 379500
rect 88334 379488 88340 379500
rect 54536 379460 88340 379488
rect 54536 379448 54542 379460
rect 88334 379448 88340 379460
rect 88392 379448 88398 379500
rect 92382 379448 92388 379500
rect 92440 379488 92446 379500
rect 219526 379488 219532 379500
rect 92440 379460 213684 379488
rect 92440 379448 92446 379460
rect 86586 379380 86592 379432
rect 86644 379420 86650 379432
rect 210050 379420 210056 379432
rect 86644 379392 210056 379420
rect 86644 379380 86650 379392
rect 210050 379380 210056 379392
rect 210108 379420 210114 379432
rect 211522 379420 211528 379432
rect 210108 379392 211528 379420
rect 210108 379380 210114 379392
rect 211522 379380 211528 379392
rect 211580 379380 211586 379432
rect 85482 379312 85488 379364
rect 85540 379352 85546 379364
rect 208762 379352 208768 379364
rect 85540 379324 208768 379352
rect 85540 379312 85546 379324
rect 208762 379312 208768 379324
rect 208820 379312 208826 379364
rect 88794 379244 88800 379296
rect 88852 379284 88858 379296
rect 210326 379284 210332 379296
rect 88852 379256 210332 379284
rect 88852 379244 88858 379256
rect 210326 379244 210332 379256
rect 210384 379284 210390 379296
rect 210970 379284 210976 379296
rect 210384 379256 210976 379284
rect 210384 379244 210390 379256
rect 210970 379244 210976 379256
rect 211028 379244 211034 379296
rect 213656 379284 213684 379460
rect 215864 379460 219532 379488
rect 213730 379380 213736 379432
rect 213788 379420 213794 379432
rect 215864 379420 215892 379460
rect 219526 379448 219532 379460
rect 219584 379488 219590 379500
rect 273254 379488 273260 379500
rect 219584 379460 273260 379488
rect 219584 379448 219590 379460
rect 273254 379448 273260 379460
rect 273312 379448 273318 379500
rect 291838 379448 291844 379500
rect 291896 379488 291902 379500
rect 320910 379488 320916 379500
rect 291896 379460 320916 379488
rect 291896 379448 291902 379460
rect 320910 379448 320916 379460
rect 320968 379448 320974 379500
rect 369596 379488 369624 379584
rect 369670 379516 369676 379568
rect 369728 379556 369734 379568
rect 371234 379556 371240 379568
rect 369728 379528 371240 379556
rect 369728 379516 369734 379528
rect 371234 379516 371240 379528
rect 371292 379556 371298 379568
rect 373966 379556 373994 379596
rect 376478 379584 376484 379636
rect 376536 379624 376542 379636
rect 376662 379624 376668 379636
rect 376536 379596 376668 379624
rect 376536 379584 376542 379596
rect 376662 379584 376668 379596
rect 376720 379624 376726 379636
rect 420638 379624 420644 379636
rect 376720 379596 420644 379624
rect 376720 379584 376726 379596
rect 420638 379584 420644 379596
rect 420696 379584 420702 379636
rect 431126 379556 431132 379568
rect 371292 379528 371648 379556
rect 373966 379528 431132 379556
rect 371292 379516 371298 379528
rect 369762 379488 369768 379500
rect 369596 379460 369768 379488
rect 369762 379448 369768 379460
rect 369820 379448 369826 379500
rect 371620 379488 371648 379528
rect 431126 379516 431132 379528
rect 431184 379516 431190 379568
rect 437934 379488 437940 379500
rect 371620 379460 437940 379488
rect 437934 379448 437940 379460
rect 437992 379448 437998 379500
rect 213788 379392 215892 379420
rect 213788 379380 213794 379392
rect 218238 379380 218244 379432
rect 218296 379420 218302 379432
rect 269758 379420 269764 379432
rect 218296 379392 269764 379420
rect 218296 379380 218302 379392
rect 269758 379380 269764 379392
rect 269816 379380 269822 379432
rect 298002 379380 298008 379432
rect 298060 379420 298066 379432
rect 305822 379420 305828 379432
rect 298060 379392 305828 379420
rect 298060 379380 298066 379392
rect 305822 379380 305828 379392
rect 305880 379380 305886 379432
rect 378226 379380 378232 379432
rect 378284 379420 378290 379432
rect 434254 379420 434260 379432
rect 378284 379392 434260 379420
rect 378284 379380 378290 379392
rect 434254 379380 434260 379392
rect 434312 379380 434318 379432
rect 220446 379312 220452 379364
rect 220504 379352 220510 379364
rect 271046 379352 271052 379364
rect 220504 379324 271052 379352
rect 220504 379312 220510 379324
rect 271046 379312 271052 379324
rect 271104 379312 271110 379364
rect 375190 379312 375196 379364
rect 375248 379352 375254 379364
rect 408310 379352 408316 379364
rect 375248 379324 408316 379352
rect 375248 379312 375254 379324
rect 408310 379312 408316 379324
rect 408368 379312 408374 379364
rect 218146 379284 218152 379296
rect 213656 379256 218152 379284
rect 218146 379244 218152 379256
rect 218204 379284 218210 379296
rect 220998 379284 221004 379296
rect 218204 379256 221004 379284
rect 218204 379244 218210 379256
rect 220998 379244 221004 379256
rect 221056 379284 221062 379296
rect 222010 379284 222016 379296
rect 221056 379256 222016 379284
rect 221056 379244 221062 379256
rect 222010 379244 222016 379256
rect 222068 379244 222074 379296
rect 91370 379176 91376 379228
rect 91428 379216 91434 379228
rect 91428 379188 200114 379216
rect 91428 379176 91434 379188
rect 44634 379108 44640 379160
rect 44692 379148 44698 379160
rect 90726 379148 90732 379160
rect 44692 379120 90732 379148
rect 44692 379108 44698 379120
rect 90726 379108 90732 379120
rect 90784 379108 90790 379160
rect 90818 379108 90824 379160
rect 90876 379148 90882 379160
rect 195974 379148 195980 379160
rect 90876 379120 195980 379148
rect 90876 379108 90882 379120
rect 195974 379108 195980 379120
rect 196032 379108 196038 379160
rect 200086 379148 200114 379188
rect 211154 379148 211160 379160
rect 200086 379120 211160 379148
rect 211154 379108 211160 379120
rect 211212 379148 211218 379160
rect 221458 379148 221464 379160
rect 211212 379120 221464 379148
rect 211212 379108 211218 379120
rect 221458 379108 221464 379120
rect 221516 379108 221522 379160
rect 44818 379040 44824 379092
rect 44876 379080 44882 379092
rect 93486 379080 93492 379092
rect 44876 379052 93492 379080
rect 44876 379040 44882 379052
rect 93486 379040 93492 379052
rect 93544 379040 93550 379092
rect 93578 379040 93584 379092
rect 93636 379080 93642 379092
rect 198642 379080 198648 379092
rect 93636 379052 198648 379080
rect 93636 379040 93642 379052
rect 198642 379040 198648 379052
rect 198700 379080 198706 379092
rect 220814 379080 220820 379092
rect 198700 379052 220820 379080
rect 198700 379040 198706 379052
rect 220814 379040 220820 379052
rect 220872 379080 220878 379092
rect 222102 379080 222108 379092
rect 220872 379052 222108 379080
rect 220872 379040 220878 379052
rect 222102 379040 222108 379052
rect 222160 379040 222166 379092
rect 46198 378972 46204 379024
rect 46256 379012 46262 379024
rect 108206 379012 108212 379024
rect 46256 378984 108212 379012
rect 46256 378972 46262 378984
rect 108206 378972 108212 378984
rect 108264 378972 108270 379024
rect 115842 378972 115848 379024
rect 115900 379012 115906 379024
rect 219894 379012 219900 379024
rect 115900 378984 219900 379012
rect 115900 378972 115906 378984
rect 219894 378972 219900 378984
rect 219952 379012 219958 379024
rect 220722 379012 220728 379024
rect 219952 378984 220728 379012
rect 219952 378972 219958 378984
rect 220722 378972 220728 378984
rect 220780 378972 220786 379024
rect 58618 378904 58624 378956
rect 58676 378944 58682 378956
rect 105354 378944 105360 378956
rect 58676 378916 105360 378944
rect 58676 378904 58682 378916
rect 105354 378904 105360 378916
rect 105412 378904 105418 378956
rect 112346 378904 112352 378956
rect 112404 378944 112410 378956
rect 204070 378944 204076 378956
rect 112404 378916 204076 378944
rect 112404 378904 112410 378916
rect 204070 378904 204076 378916
rect 204128 378944 204134 378956
rect 211706 378944 211712 378956
rect 204128 378916 211712 378944
rect 204128 378904 204134 378916
rect 211706 378904 211712 378916
rect 211764 378904 211770 378956
rect 368382 378904 368388 378956
rect 368440 378944 368446 378956
rect 379606 378944 379612 378956
rect 368440 378916 379612 378944
rect 368440 378904 368446 378916
rect 379606 378904 379612 378916
rect 379664 378904 379670 378956
rect 379974 378904 379980 378956
rect 380032 378944 380038 378956
rect 396074 378944 396080 378956
rect 380032 378916 396080 378944
rect 380032 378904 380038 378916
rect 396074 378904 396080 378916
rect 396132 378904 396138 378956
rect 58434 378836 58440 378888
rect 58492 378876 58498 378888
rect 103514 378876 103520 378888
rect 58492 378848 103520 378876
rect 58492 378836 58498 378848
rect 103514 378836 103520 378848
rect 103572 378836 103578 378888
rect 117130 378836 117136 378888
rect 117188 378876 117194 378888
rect 205542 378876 205548 378888
rect 117188 378848 205548 378876
rect 117188 378836 117194 378848
rect 205542 378836 205548 378848
rect 205600 378836 205606 378888
rect 213822 378836 213828 378888
rect 213880 378876 213886 378888
rect 214098 378876 214104 378888
rect 213880 378848 214104 378876
rect 213880 378836 213886 378848
rect 214098 378836 214104 378848
rect 214156 378836 214162 378888
rect 266446 378836 266452 378888
rect 266504 378876 266510 378888
rect 268286 378876 268292 378888
rect 266504 378848 268292 378876
rect 266504 378836 266510 378848
rect 268286 378836 268292 378848
rect 268344 378836 268350 378888
rect 360746 378836 360752 378888
rect 360804 378876 360810 378888
rect 379514 378876 379520 378888
rect 360804 378848 379520 378876
rect 360804 378836 360810 378848
rect 379514 378836 379520 378848
rect 379572 378836 379578 378888
rect 56410 378768 56416 378820
rect 56468 378808 56474 378820
rect 101030 378808 101036 378820
rect 56468 378780 101036 378808
rect 56468 378768 56474 378780
rect 101030 378768 101036 378780
rect 101088 378768 101094 378820
rect 195974 378768 195980 378820
rect 196032 378808 196038 378820
rect 197262 378808 197268 378820
rect 196032 378780 197268 378808
rect 196032 378768 196038 378780
rect 197262 378768 197268 378780
rect 197320 378808 197326 378820
rect 197320 378780 219434 378808
rect 197320 378768 197326 378780
rect 77202 378700 77208 378752
rect 77260 378740 77266 378752
rect 99374 378740 99380 378752
rect 77260 378712 99380 378740
rect 77260 378700 77266 378712
rect 99374 378700 99380 378712
rect 99432 378700 99438 378752
rect 211522 378700 211528 378752
rect 211580 378740 211586 378752
rect 218330 378740 218336 378752
rect 211580 378712 218336 378740
rect 211580 378700 211586 378712
rect 218330 378700 218336 378712
rect 218388 378700 218394 378752
rect 219406 378740 219434 378780
rect 220630 378768 220636 378820
rect 220688 378808 220694 378820
rect 248598 378808 248604 378820
rect 220688 378780 248604 378808
rect 220688 378768 220694 378780
rect 248598 378768 248604 378780
rect 248656 378768 248662 378820
rect 374546 378768 374552 378820
rect 374604 378808 374610 378820
rect 396350 378808 396356 378820
rect 374604 378780 396356 378808
rect 374604 378768 374610 378780
rect 396350 378768 396356 378780
rect 396408 378768 396414 378820
rect 219526 378740 219532 378752
rect 219406 378712 219532 378740
rect 219526 378700 219532 378712
rect 219584 378740 219590 378752
rect 250070 378740 250076 378752
rect 219584 378712 250076 378740
rect 219584 378700 219590 378712
rect 250070 378700 250076 378712
rect 250128 378700 250134 378752
rect 343542 378700 343548 378752
rect 343600 378740 343606 378752
rect 503622 378740 503628 378752
rect 343600 378712 503628 378740
rect 343600 378700 343606 378712
rect 503622 378700 503628 378712
rect 503680 378700 503686 378752
rect 50154 378632 50160 378684
rect 50212 378672 50218 378684
rect 98454 378672 98460 378684
rect 50212 378644 98460 378672
rect 50212 378632 50218 378644
rect 98454 378632 98460 378644
rect 98512 378632 98518 378684
rect 210970 378632 210976 378684
rect 211028 378672 211034 378684
rect 219986 378672 219992 378684
rect 211028 378644 219992 378672
rect 211028 378632 211034 378644
rect 219986 378632 219992 378644
rect 220044 378672 220050 378684
rect 220630 378672 220636 378684
rect 220044 378644 220636 378672
rect 220044 378632 220050 378644
rect 220630 378632 220636 378644
rect 220688 378632 220694 378684
rect 221090 378632 221096 378684
rect 221148 378672 221154 378684
rect 221458 378672 221464 378684
rect 221148 378644 221464 378672
rect 221148 378632 221154 378644
rect 221458 378632 221464 378644
rect 221516 378672 221522 378684
rect 251174 378672 251180 378684
rect 221516 378644 251180 378672
rect 221516 378632 221522 378644
rect 251174 378632 251180 378644
rect 251232 378632 251238 378684
rect 369578 378632 369584 378684
rect 369636 378672 369642 378684
rect 398190 378672 398196 378684
rect 369636 378644 398196 378672
rect 369636 378632 369642 378644
rect 398190 378632 398196 378644
rect 398248 378632 398254 378684
rect 47854 378564 47860 378616
rect 47912 378604 47918 378616
rect 96062 378604 96068 378616
rect 47912 378576 96068 378604
rect 47912 378564 47918 378576
rect 96062 378564 96068 378576
rect 96120 378564 96126 378616
rect 205634 378564 205640 378616
rect 205692 378604 205698 378616
rect 206830 378604 206836 378616
rect 205692 378576 206836 378604
rect 205692 378564 205698 378576
rect 206830 378564 206836 378576
rect 206888 378604 206894 378616
rect 219618 378604 219624 378616
rect 206888 378576 219624 378604
rect 206888 378564 206894 378576
rect 219618 378564 219624 378576
rect 219676 378604 219682 378616
rect 220446 378604 220452 378616
rect 219676 378576 220452 378604
rect 219676 378564 219682 378576
rect 220446 378564 220452 378576
rect 220504 378564 220510 378616
rect 222010 378564 222016 378616
rect 222068 378604 222074 378616
rect 252278 378604 252284 378616
rect 222068 378576 252284 378604
rect 222068 378564 222074 378576
rect 252278 378564 252284 378576
rect 252336 378564 252342 378616
rect 342898 378564 342904 378616
rect 342956 378604 342962 378616
rect 343450 378604 343456 378616
rect 342956 378576 343456 378604
rect 342956 378564 342962 378576
rect 343450 378564 343456 378576
rect 343508 378604 343514 378616
rect 358814 378604 358820 378616
rect 343508 378576 358820 378604
rect 343508 378564 343514 378576
rect 358814 378564 358820 378576
rect 358872 378604 358878 378616
rect 359274 378604 359280 378616
rect 358872 378576 359280 378604
rect 358872 378564 358878 378576
rect 359274 378564 359280 378576
rect 359332 378564 359338 378616
rect 370406 378564 370412 378616
rect 370464 378604 370470 378616
rect 376478 378604 376484 378616
rect 370464 378576 376484 378604
rect 370464 378564 370470 378576
rect 376478 378564 376484 378576
rect 376536 378604 376542 378616
rect 405826 378604 405832 378616
rect 376536 378576 405832 378604
rect 376536 378564 376542 378576
rect 405826 378564 405832 378576
rect 405884 378564 405890 378616
rect 113450 378496 113456 378548
rect 113508 378536 113514 378548
rect 212994 378536 213000 378548
rect 113508 378508 213000 378536
rect 113508 378496 113514 378508
rect 212994 378496 213000 378508
rect 213052 378536 213058 378548
rect 213730 378536 213736 378548
rect 213052 378508 213736 378536
rect 213052 378496 213058 378508
rect 213730 378496 213736 378508
rect 213788 378496 213794 378548
rect 222102 378496 222108 378548
rect 222160 378536 222166 378548
rect 253382 378536 253388 378548
rect 222160 378508 253388 378536
rect 222160 378496 222166 378508
rect 253382 378496 253388 378508
rect 253440 378496 253446 378548
rect 262214 378496 262220 378548
rect 262272 378536 262278 378548
rect 266354 378536 266360 378548
rect 262272 378508 266360 378536
rect 262272 378496 262278 378508
rect 266354 378496 266360 378508
rect 266412 378496 266418 378548
rect 280062 378496 280068 378548
rect 280120 378536 280126 378548
rect 360010 378536 360016 378548
rect 280120 378508 360016 378536
rect 280120 378496 280126 378508
rect 360010 378496 360016 378508
rect 360068 378496 360074 378548
rect 368290 378536 368296 378548
rect 364306 378508 368296 378536
rect 208762 378428 208768 378480
rect 208820 378468 208826 378480
rect 212350 378468 212356 378480
rect 208820 378440 212356 378468
rect 208820 378428 208826 378440
rect 212350 378428 212356 378440
rect 212408 378468 212414 378480
rect 244918 378468 244924 378480
rect 212408 378440 244924 378468
rect 212408 378428 212414 378440
rect 244918 378428 244924 378440
rect 244976 378428 244982 378480
rect 276014 378428 276020 378480
rect 276072 378468 276078 378480
rect 277026 378468 277032 378480
rect 276072 378440 277032 378468
rect 276072 378428 276078 378440
rect 277026 378428 277032 378440
rect 277084 378468 277090 378480
rect 356974 378468 356980 378480
rect 277084 378440 356980 378468
rect 277084 378428 277090 378440
rect 356974 378428 356980 378440
rect 357032 378428 357038 378480
rect 114462 378360 114468 378412
rect 114520 378400 114526 378412
rect 207014 378400 207020 378412
rect 114520 378372 207020 378400
rect 114520 378360 114526 378372
rect 207014 378360 207020 378372
rect 207072 378400 207078 378412
rect 207566 378400 207572 378412
rect 207072 378372 207572 378400
rect 207072 378360 207078 378372
rect 207566 378360 207572 378372
rect 207624 378360 207630 378412
rect 210326 378360 210332 378412
rect 210384 378400 210390 378412
rect 239582 378400 239588 378412
rect 210384 378372 239588 378400
rect 210384 378360 210390 378372
rect 239582 378360 239588 378372
rect 239640 378400 239646 378412
rect 364306 378400 364334 378508
rect 368290 378496 368296 378508
rect 368348 378536 368354 378548
rect 399478 378536 399484 378548
rect 368348 378508 399484 378536
rect 368348 378496 368354 378508
rect 399478 378496 399484 378508
rect 399536 378496 399542 378548
rect 379606 378428 379612 378480
rect 379664 378468 379670 378480
rect 412358 378468 412364 378480
rect 379664 378440 412364 378468
rect 379664 378428 379670 378440
rect 412358 378428 412364 378440
rect 412416 378428 412422 378480
rect 239640 378372 364334 378400
rect 239640 378360 239646 378372
rect 369026 378360 369032 378412
rect 369084 378400 369090 378412
rect 373810 378400 373816 378412
rect 369084 378372 373816 378400
rect 369084 378360 369090 378372
rect 373810 378360 373816 378372
rect 373868 378400 373874 378412
rect 373868 378372 373994 378400
rect 373868 378360 373874 378372
rect 111242 378292 111248 378344
rect 111300 378332 111306 378344
rect 205634 378332 205640 378344
rect 111300 378304 205640 378332
rect 111300 378292 111306 378304
rect 205634 378292 205640 378304
rect 205692 378292 205698 378344
rect 205726 378292 205732 378344
rect 205784 378332 205790 378344
rect 206922 378332 206928 378344
rect 205784 378304 206928 378332
rect 205784 378292 205790 378304
rect 206922 378292 206928 378304
rect 206980 378332 206986 378344
rect 238202 378332 238208 378344
rect 206980 378304 238208 378332
rect 206980 378292 206986 378304
rect 238202 378292 238208 378304
rect 238260 378332 238266 378344
rect 369578 378332 369584 378344
rect 238260 378304 369584 378332
rect 238260 378292 238266 378304
rect 369578 378292 369584 378304
rect 369636 378292 369642 378344
rect 373966 378332 373994 378372
rect 379514 378360 379520 378412
rect 379572 378400 379578 378412
rect 411254 378400 411260 378412
rect 379572 378372 411260 378400
rect 379572 378360 379578 378372
rect 411254 378360 411260 378372
rect 411312 378360 411318 378412
rect 511902 378360 511908 378412
rect 511960 378400 511966 378412
rect 517514 378400 517520 378412
rect 511960 378372 517520 378400
rect 511960 378360 511966 378372
rect 517514 378360 517520 378372
rect 517572 378360 517578 378412
rect 407574 378332 407580 378344
rect 373966 378304 407580 378332
rect 407574 378292 407580 378304
rect 407632 378292 407638 378344
rect 204806 378224 204812 378276
rect 204864 378264 204870 378276
rect 210970 378264 210976 378276
rect 204864 378236 210976 378264
rect 204864 378224 204870 378236
rect 210970 378224 210976 378236
rect 211028 378224 211034 378276
rect 218238 378264 218244 378276
rect 211632 378236 218244 378264
rect 44726 378156 44732 378208
rect 44784 378196 44790 378208
rect 47762 378196 47768 378208
rect 44784 378168 47768 378196
rect 44784 378156 44790 378168
rect 47762 378156 47768 378168
rect 47820 378196 47826 378208
rect 80422 378196 80428 378208
rect 47820 378168 80428 378196
rect 47820 378156 47826 378168
rect 80422 378156 80428 378168
rect 80480 378156 80486 378208
rect 109770 378156 109776 378208
rect 109828 378196 109834 378208
rect 211632 378196 211660 378236
rect 218238 378224 218244 378236
rect 218296 378224 218302 378276
rect 218330 378224 218336 378276
rect 218388 378264 218394 378276
rect 246206 378264 246212 378276
rect 218388 378236 246212 378264
rect 218388 378224 218394 378236
rect 246206 378224 246212 378236
rect 246264 378224 246270 378276
rect 263870 378224 263876 378276
rect 263928 378264 263934 378276
rect 267550 378264 267556 378276
rect 263928 378236 267556 378264
rect 263928 378224 263934 378236
rect 267550 378224 267556 378236
rect 267608 378224 267614 378276
rect 274634 378224 274640 378276
rect 274692 378264 274698 378276
rect 275738 378264 275744 378276
rect 274692 378236 275744 378264
rect 274692 378224 274698 378236
rect 275738 378224 275744 378236
rect 275796 378264 275802 378276
rect 356606 378264 356612 378276
rect 275796 378236 356612 378264
rect 275796 378224 275802 378236
rect 356606 378224 356612 378236
rect 356664 378224 356670 378276
rect 359274 378224 359280 378276
rect 359332 378264 359338 378276
rect 359332 378236 489914 378264
rect 359332 378224 359338 378236
rect 109828 378168 211660 378196
rect 109828 378156 109834 378168
rect 198918 378128 198924 378140
rect 180766 378100 198924 378128
rect 40862 378020 40868 378072
rect 40920 378060 40926 378072
rect 180766 378060 180794 378100
rect 198918 378088 198924 378100
rect 198976 378128 198982 378140
rect 199654 378128 199660 378140
rect 198976 378100 199660 378128
rect 198976 378088 198982 378100
rect 199654 378088 199660 378100
rect 199712 378088 199718 378140
rect 210988 378072 211016 378168
rect 211706 378156 211712 378208
rect 211764 378196 211770 378208
rect 272150 378196 272156 378208
rect 211764 378168 272156 378196
rect 211764 378156 211770 378168
rect 272150 378156 272156 378168
rect 272208 378156 272214 378208
rect 273254 378156 273260 378208
rect 273312 378196 273318 378208
rect 285950 378196 285956 378208
rect 273312 378168 285956 378196
rect 273312 378156 273318 378168
rect 285950 378156 285956 378168
rect 286008 378156 286014 378208
rect 489886 378196 489914 378236
rect 503622 378224 503628 378276
rect 503680 378264 503686 378276
rect 517606 378264 517612 378276
rect 503680 378236 517612 378264
rect 503680 378224 503686 378236
rect 517606 378224 517612 378236
rect 517664 378264 517670 378276
rect 580258 378264 580264 378276
rect 517664 378236 580264 378264
rect 517664 378224 517670 378236
rect 580258 378224 580264 378236
rect 580316 378224 580322 378276
rect 503346 378196 503352 378208
rect 489886 378168 503352 378196
rect 503346 378156 503352 378168
rect 503404 378196 503410 378208
rect 517698 378196 517704 378208
rect 503404 378168 517704 378196
rect 503404 378156 503410 378168
rect 517698 378156 517704 378168
rect 517756 378196 517762 378208
rect 580166 378196 580172 378208
rect 517756 378168 580172 378196
rect 517756 378156 517762 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 217410 378088 217416 378140
rect 217468 378128 217474 378140
rect 310974 378128 310980 378140
rect 217468 378100 310980 378128
rect 217468 378088 217474 378100
rect 310974 378088 310980 378100
rect 311032 378088 311038 378140
rect 360838 378088 360844 378140
rect 360896 378128 360902 378140
rect 473446 378128 473452 378140
rect 360896 378100 473452 378128
rect 360896 378088 360902 378100
rect 473446 378088 473452 378100
rect 473504 378088 473510 378140
rect 40920 378032 180794 378060
rect 40920 378020 40926 378032
rect 205358 378020 205364 378072
rect 205416 378060 205422 378072
rect 206186 378060 206192 378072
rect 205416 378032 206192 378060
rect 205416 378020 205422 378032
rect 206186 378020 206192 378032
rect 206244 378020 206250 378072
rect 210970 378020 210976 378072
rect 211028 378020 211034 378072
rect 212258 378020 212264 378072
rect 212316 378060 212322 378072
rect 325878 378060 325884 378072
rect 212316 378032 325884 378060
rect 212316 378020 212322 378032
rect 325878 378020 325884 378032
rect 325936 378020 325942 378072
rect 368934 378020 368940 378072
rect 368992 378060 368998 378072
rect 480622 378060 480628 378072
rect 368992 378032 480628 378060
rect 368992 378020 368998 378032
rect 480622 378020 480628 378032
rect 480680 378020 480686 378072
rect 54294 377952 54300 378004
rect 54352 377992 54358 378004
rect 182358 377992 182364 378004
rect 54352 377964 182364 377992
rect 54352 377952 54358 377964
rect 182358 377952 182364 377964
rect 182416 377992 182422 378004
rect 182910 377992 182916 378004
rect 182416 377964 182916 377992
rect 182416 377952 182422 377964
rect 182910 377952 182916 377964
rect 182968 377952 182974 378004
rect 205450 377952 205456 378004
rect 205508 377992 205514 378004
rect 206554 377992 206560 378004
rect 205508 377964 206560 377992
rect 205508 377952 205514 377964
rect 206554 377952 206560 377964
rect 206612 377952 206618 378004
rect 206646 377952 206652 378004
rect 206704 377992 206710 378004
rect 317782 377992 317788 378004
rect 206704 377964 317788 377992
rect 206704 377952 206710 377964
rect 317782 377952 317788 377964
rect 317840 377952 317846 378004
rect 376570 377952 376576 378004
rect 376628 377992 376634 378004
rect 485958 377992 485964 378004
rect 376628 377964 485964 377992
rect 376628 377952 376634 377964
rect 485958 377952 485964 377964
rect 486016 377952 486022 378004
rect 54386 377884 54392 377936
rect 54444 377924 54450 377936
rect 182266 377924 182272 377936
rect 54444 377896 182272 377924
rect 54444 377884 54450 377896
rect 182266 377884 182272 377896
rect 182324 377884 182330 377936
rect 200206 377884 200212 377936
rect 200264 377924 200270 377936
rect 307846 377924 307852 377936
rect 200264 377896 307852 377924
rect 200264 377884 200270 377896
rect 307846 377884 307852 377896
rect 307904 377884 307910 377936
rect 357894 377884 357900 377936
rect 357952 377924 357958 377936
rect 460934 377924 460940 377936
rect 357952 377896 460940 377924
rect 357952 377884 357958 377896
rect 460934 377884 460940 377896
rect 460992 377884 460998 377936
rect 196618 377816 196624 377868
rect 196676 377856 196682 377868
rect 273254 377856 273260 377868
rect 196676 377828 273260 377856
rect 196676 377816 196682 377828
rect 273254 377816 273260 377828
rect 273312 377816 273318 377868
rect 367554 377816 367560 377868
rect 367612 377856 367618 377868
rect 463510 377856 463516 377868
rect 367612 377828 463516 377856
rect 367612 377816 367618 377828
rect 463510 377816 463516 377828
rect 463568 377816 463574 377868
rect 150986 377748 150992 377800
rect 151044 377788 151050 377800
rect 198090 377788 198096 377800
rect 151044 377760 198096 377788
rect 151044 377748 151050 377760
rect 198090 377748 198096 377760
rect 198148 377748 198154 377800
rect 198458 377748 198464 377800
rect 198516 377788 198522 377800
rect 298094 377788 298100 377800
rect 198516 377760 298100 377788
rect 198516 377748 198522 377760
rect 298094 377748 298100 377760
rect 298152 377748 298158 377800
rect 372982 377748 372988 377800
rect 373040 377788 373046 377800
rect 455598 377788 455604 377800
rect 373040 377760 455604 377788
rect 373040 377748 373046 377760
rect 455598 377748 455604 377760
rect 455656 377748 455662 377800
rect 197998 377680 198004 377732
rect 198056 377720 198062 377732
rect 295886 377720 295892 377732
rect 198056 377692 295892 377720
rect 198056 377680 198062 377692
rect 295886 377680 295892 377692
rect 295944 377680 295950 377732
rect 370314 377680 370320 377732
rect 370372 377720 370378 377732
rect 453022 377720 453028 377732
rect 370372 377692 453028 377720
rect 370372 377680 370378 377692
rect 453022 377680 453028 377692
rect 453080 377680 453086 377732
rect 197538 377612 197544 377664
rect 197596 377652 197602 377664
rect 293310 377652 293316 377664
rect 197596 377624 293316 377652
rect 197596 377612 197602 377624
rect 293310 377612 293316 377624
rect 293368 377612 293374 377664
rect 367646 377612 367652 377664
rect 367704 377652 367710 377664
rect 450998 377652 451004 377664
rect 367704 377624 451004 377652
rect 367704 377612 367710 377624
rect 450998 377612 451004 377624
rect 451056 377612 451062 377664
rect 197078 377544 197084 377596
rect 197136 377584 197142 377596
rect 290182 377584 290188 377596
rect 197136 377556 290188 377584
rect 197136 377544 197142 377556
rect 290182 377544 290188 377556
rect 290240 377544 290246 377596
rect 373166 377544 373172 377596
rect 373224 377584 373230 377596
rect 428182 377584 428188 377596
rect 373224 377556 428188 377584
rect 373224 377544 373230 377556
rect 428182 377544 428188 377556
rect 428240 377544 428246 377596
rect 196710 377476 196716 377528
rect 196768 377516 196774 377528
rect 287698 377516 287704 377528
rect 196768 377488 287704 377516
rect 196768 377476 196774 377488
rect 287698 377476 287704 377488
rect 287756 377476 287762 377528
rect 377214 377476 377220 377528
rect 377272 377516 377278 377528
rect 410334 377516 410340 377528
rect 377272 377488 410340 377516
rect 377272 377476 377278 377488
rect 410334 377476 410340 377488
rect 410392 377476 410398 377528
rect 199378 377408 199384 377460
rect 199436 377448 199442 377460
rect 280798 377448 280804 377460
rect 199436 377420 280804 377448
rect 199436 377408 199442 377420
rect 280798 377408 280804 377420
rect 280856 377408 280862 377460
rect 363506 377408 363512 377460
rect 363564 377448 363570 377460
rect 379882 377448 379888 377460
rect 363564 377420 379888 377448
rect 363564 377408 363570 377420
rect 379882 377408 379888 377420
rect 379940 377448 379946 377460
rect 414566 377448 414572 377460
rect 379940 377420 414572 377448
rect 379940 377408 379946 377420
rect 414566 377408 414572 377420
rect 414624 377408 414630 377460
rect 196802 377340 196808 377392
rect 196860 377380 196866 377392
rect 278406 377380 278412 377392
rect 196860 377352 278412 377380
rect 196860 377340 196866 377352
rect 278406 377340 278412 377352
rect 278464 377340 278470 377392
rect 366174 377340 366180 377392
rect 366232 377380 366238 377392
rect 372246 377380 372252 377392
rect 366232 377352 372252 377380
rect 366232 377340 366238 377352
rect 372246 377340 372252 377352
rect 372304 377380 372310 377392
rect 402974 377380 402980 377392
rect 372304 377352 402980 377380
rect 372304 377340 372310 377352
rect 402974 377340 402980 377352
rect 403032 377340 403038 377392
rect 146018 377272 146024 377324
rect 146076 377312 146082 377324
rect 207290 377312 207296 377324
rect 146076 377284 207296 377312
rect 146076 377272 146082 377284
rect 207290 377272 207296 377284
rect 207348 377272 207354 377324
rect 213086 377272 213092 377324
rect 213144 377312 213150 377324
rect 270954 377312 270960 377324
rect 213144 377284 270960 377312
rect 213144 377272 213150 377284
rect 270954 377272 270960 377284
rect 271012 377272 271018 377324
rect 104250 377204 104256 377256
rect 104308 377244 104314 377256
rect 215662 377244 215668 377256
rect 104308 377216 215668 377244
rect 104308 377204 104314 377216
rect 215662 377204 215668 377216
rect 215720 377204 215726 377256
rect 217042 377204 217048 377256
rect 217100 377244 217106 377256
rect 217686 377244 217692 377256
rect 217100 377216 217692 377244
rect 217100 377204 217106 377216
rect 217686 377204 217692 377216
rect 217744 377204 217750 377256
rect 264974 377244 264980 377256
rect 219406 377216 264980 377244
rect 141050 377136 141056 377188
rect 141108 377176 141114 377188
rect 201862 377176 201868 377188
rect 141108 377148 201868 377176
rect 141108 377136 141114 377148
rect 201862 377136 201868 377148
rect 201920 377136 201926 377188
rect 219250 377136 219256 377188
rect 219308 377176 219314 377188
rect 219406 377176 219434 377216
rect 264974 377204 264980 377216
rect 265032 377204 265038 377256
rect 219308 377148 219434 377176
rect 219308 377136 219314 377148
rect 153562 377068 153568 377120
rect 153620 377108 153626 377120
rect 200390 377108 200396 377120
rect 153620 377080 200396 377108
rect 153620 377068 153626 377080
rect 200390 377068 200396 377080
rect 200448 377068 200454 377120
rect 42518 377000 42524 377052
rect 42576 377040 42582 377052
rect 199746 377040 199752 377052
rect 42576 377012 199752 377040
rect 42576 377000 42582 377012
rect 199746 377000 199752 377012
rect 199804 377000 199810 377052
rect 369762 377000 369768 377052
rect 369820 377000 369826 377052
rect 47578 376932 47584 376984
rect 47636 376972 47642 376984
rect 217042 376972 217048 376984
rect 47636 376944 217048 376972
rect 47636 376932 47642 376944
rect 217042 376932 217048 376944
rect 217100 376932 217106 376984
rect 369578 376796 369584 376848
rect 369636 376836 369642 376848
rect 369780 376836 369808 377000
rect 369636 376808 369808 376836
rect 369636 376796 369642 376808
rect 368382 376728 368388 376780
rect 368440 376768 368446 376780
rect 378134 376768 378140 376780
rect 368440 376740 378140 376768
rect 368440 376728 368446 376740
rect 378134 376728 378140 376740
rect 378192 376768 378198 376780
rect 378594 376768 378600 376780
rect 378192 376740 378600 376768
rect 378192 376728 378198 376740
rect 378594 376728 378600 376740
rect 378652 376728 378658 376780
rect 198826 376660 198832 376712
rect 198884 376700 198890 376712
rect 300854 376700 300860 376712
rect 198884 376672 300860 376700
rect 198884 376660 198890 376672
rect 300854 376660 300860 376672
rect 300912 376660 300918 376712
rect 357158 376660 357164 376712
rect 357216 376700 357222 376712
rect 470870 376700 470876 376712
rect 357216 376672 470876 376700
rect 357216 376660 357222 376672
rect 470870 376660 470876 376672
rect 470928 376660 470934 376712
rect 99466 376592 99472 376644
rect 99524 376632 99530 376644
rect 214374 376632 214380 376644
rect 99524 376604 214380 376632
rect 99524 376592 99530 376604
rect 214374 376592 214380 376604
rect 214432 376592 214438 376644
rect 219802 376592 219808 376644
rect 219860 376632 219866 376644
rect 302510 376632 302516 376644
rect 219860 376604 302516 376632
rect 219860 376592 219866 376604
rect 302510 376592 302516 376604
rect 302568 376592 302574 376644
rect 364150 376592 364156 376644
rect 364208 376632 364214 376644
rect 474734 376632 474740 376644
rect 364208 376604 474740 376632
rect 364208 376592 364214 376604
rect 474734 376592 474740 376604
rect 474792 376592 474798 376644
rect 101858 376524 101864 376576
rect 101916 376564 101922 376576
rect 214006 376564 214012 376576
rect 101916 376536 214012 376564
rect 101916 376524 101922 376536
rect 214006 376524 214012 376536
rect 214064 376524 214070 376576
rect 214466 376524 214472 376576
rect 214524 376564 214530 376576
rect 276106 376564 276112 376576
rect 214524 376536 276112 376564
rect 214524 376524 214530 376536
rect 276106 376524 276112 376536
rect 276164 376524 276170 376576
rect 367002 376524 367008 376576
rect 367060 376564 367066 376576
rect 477494 376564 477500 376576
rect 367060 376536 477500 376564
rect 367060 376524 367066 376536
rect 477494 376524 477500 376536
rect 477552 376524 477558 376576
rect 97074 376456 97080 376508
rect 97132 376496 97138 376508
rect 205910 376496 205916 376508
rect 97132 376468 205916 376496
rect 97132 376456 97138 376468
rect 205910 376456 205916 376468
rect 205968 376456 205974 376508
rect 206738 376456 206744 376508
rect 206796 376496 206802 376508
rect 283098 376496 283104 376508
rect 206796 376468 283104 376496
rect 206796 376456 206802 376468
rect 283098 376456 283104 376468
rect 283156 376456 283162 376508
rect 374454 376456 374460 376508
rect 374512 376496 374518 376508
rect 483382 376496 483388 376508
rect 374512 376468 483388 376496
rect 374512 376456 374518 376468
rect 483382 376456 483388 376468
rect 483440 376456 483446 376508
rect 107562 376388 107568 376440
rect 107620 376428 107626 376440
rect 207290 376428 207296 376440
rect 107620 376400 207296 376428
rect 107620 376388 107626 376400
rect 207290 376388 207296 376400
rect 207348 376428 207354 376440
rect 207934 376428 207940 376440
rect 207348 376400 207940 376428
rect 207348 376388 207354 376400
rect 207934 376388 207940 376400
rect 207992 376388 207998 376440
rect 212902 376388 212908 376440
rect 212960 376428 212966 376440
rect 273438 376428 273444 376440
rect 212960 376400 273444 376428
rect 212960 376388 212966 376400
rect 273438 376388 273444 376400
rect 273496 376388 273502 376440
rect 362770 376388 362776 376440
rect 362828 376428 362834 376440
rect 467926 376428 467932 376440
rect 362828 376400 467932 376428
rect 362828 376388 362834 376400
rect 467926 376388 467932 376400
rect 467984 376388 467990 376440
rect 125962 376320 125968 376372
rect 126020 376360 126026 376372
rect 204438 376360 204444 376372
rect 126020 376332 204444 376360
rect 126020 376320 126026 376332
rect 204438 376320 204444 376332
rect 204496 376320 204502 376372
rect 208946 376320 208952 376372
rect 209004 376360 209010 376372
rect 263594 376360 263600 376372
rect 209004 376332 263600 376360
rect 209004 376320 209010 376332
rect 263594 376320 263600 376332
rect 263652 376320 263658 376372
rect 364794 376320 364800 376372
rect 364852 376360 364858 376372
rect 465074 376360 465080 376372
rect 364852 376332 465080 376360
rect 364852 376320 364858 376332
rect 465074 376320 465080 376332
rect 465132 376320 465138 376372
rect 131022 376252 131028 376304
rect 131080 376292 131086 376304
rect 199010 376292 199016 376304
rect 131080 376264 199016 376292
rect 131080 376252 131086 376264
rect 199010 376252 199016 376264
rect 199068 376252 199074 376304
rect 214926 376252 214932 376304
rect 214984 376292 214990 376304
rect 268010 376292 268016 376304
rect 214984 376264 268016 376292
rect 214984 376252 214990 376264
rect 268010 376252 268016 376264
rect 268068 376252 268074 376304
rect 357066 376252 357072 376304
rect 357124 376292 357130 376304
rect 422846 376292 422852 376304
rect 357124 376264 422852 376292
rect 357124 376252 357130 376264
rect 422846 376252 422852 376264
rect 422904 376252 422910 376304
rect 133506 376184 133512 376236
rect 133564 376224 133570 376236
rect 194594 376224 194600 376236
rect 133564 376196 194600 376224
rect 133564 376184 133570 376196
rect 194594 376184 194600 376196
rect 194652 376184 194658 376236
rect 211614 376184 211620 376236
rect 211672 376224 211678 376236
rect 260926 376224 260932 376236
rect 211672 376196 260932 376224
rect 211672 376184 211678 376196
rect 260926 376184 260932 376196
rect 260984 376184 260990 376236
rect 371786 376184 371792 376236
rect 371844 376224 371850 376236
rect 430666 376224 430672 376236
rect 371844 376196 430672 376224
rect 371844 376184 371850 376196
rect 430666 376184 430672 376196
rect 430724 376184 430730 376236
rect 138474 376116 138480 376168
rect 138532 376156 138538 376168
rect 195054 376156 195060 376168
rect 138532 376128 195060 376156
rect 138532 376116 138538 376128
rect 195054 376116 195060 376128
rect 195112 376116 195118 376168
rect 210234 376116 210240 376168
rect 210292 376156 210298 376168
rect 258350 376156 258356 376168
rect 210292 376128 258356 376156
rect 210292 376116 210298 376128
rect 258350 376116 258356 376128
rect 258408 376116 258414 376168
rect 359458 376116 359464 376168
rect 359516 376156 359522 376168
rect 418430 376156 418436 376168
rect 359516 376128 418436 376156
rect 359516 376116 359522 376128
rect 418430 376116 418436 376128
rect 418488 376116 418494 376168
rect 77110 376048 77116 376100
rect 77168 376088 77174 376100
rect 204162 376088 204168 376100
rect 77168 376060 204168 376088
rect 77168 376048 77174 376060
rect 204162 376048 204168 376060
rect 204220 376048 204226 376100
rect 218606 376048 218612 376100
rect 218664 376088 218670 376100
rect 265894 376088 265900 376100
rect 218664 376060 265900 376088
rect 218664 376048 218670 376060
rect 265894 376048 265900 376060
rect 265952 376048 265958 376100
rect 378594 376048 378600 376100
rect 378652 376088 378658 376100
rect 436186 376088 436192 376100
rect 378652 376060 436192 376088
rect 378652 376048 378658 376060
rect 436186 376048 436192 376060
rect 436244 376048 436250 376100
rect 98546 375980 98552 376032
rect 98604 376020 98610 376032
rect 213086 376020 213092 376032
rect 98604 375992 213092 376020
rect 98604 375980 98610 375992
rect 213086 375980 213092 375992
rect 213144 376020 213150 376032
rect 219434 376020 219440 376032
rect 213144 375992 219440 376020
rect 213144 375980 213150 375992
rect 219434 375980 219440 375992
rect 219492 375980 219498 376032
rect 359918 375980 359924 376032
rect 359976 376020 359982 376032
rect 519078 376020 519084 376032
rect 359976 375992 519084 376020
rect 359976 375980 359982 375992
rect 519078 375980 519084 375992
rect 519136 375980 519142 376032
rect 208026 375912 208032 375964
rect 208084 375952 208090 375964
rect 250622 375952 250628 375964
rect 208084 375924 250628 375952
rect 208084 375912 208090 375924
rect 250622 375912 250628 375924
rect 250680 375912 250686 375964
rect 370958 375912 370964 375964
rect 371016 375952 371022 375964
rect 416038 375952 416044 375964
rect 371016 375924 416044 375952
rect 371016 375912 371022 375924
rect 416038 375912 416044 375924
rect 416096 375912 416102 375964
rect 217502 375844 217508 375896
rect 217560 375884 217566 375896
rect 253382 375884 253388 375896
rect 217560 375856 253388 375884
rect 217560 375844 217566 375856
rect 253382 375844 253388 375856
rect 253440 375844 253446 375896
rect 375834 375844 375840 375896
rect 375892 375884 375898 375896
rect 379330 375884 379336 375896
rect 375892 375856 379336 375884
rect 375892 375844 375898 375856
rect 379330 375844 379336 375856
rect 379388 375884 379394 375896
rect 408678 375884 408684 375896
rect 379388 375856 408684 375884
rect 379388 375844 379394 375856
rect 408678 375844 408684 375856
rect 408736 375844 408742 375896
rect 214006 375776 214012 375828
rect 214064 375816 214070 375828
rect 217410 375816 217416 375828
rect 214064 375788 217416 375816
rect 214064 375776 214070 375788
rect 217410 375776 217416 375788
rect 217468 375816 217474 375828
rect 239766 375816 239772 375828
rect 217468 375788 239772 375816
rect 217468 375776 217474 375788
rect 239766 375776 239772 375788
rect 239824 375776 239830 375828
rect 215846 375708 215852 375760
rect 215904 375748 215910 375760
rect 255958 375748 255964 375760
rect 215904 375720 255964 375748
rect 215904 375708 215910 375720
rect 255958 375708 255964 375720
rect 256016 375708 256022 375760
rect 219434 375640 219440 375692
rect 219492 375680 219498 375692
rect 220078 375680 220084 375692
rect 219492 375652 220084 375680
rect 219492 375640 219498 375652
rect 220078 375640 220084 375652
rect 220136 375640 220142 375692
rect 100754 375300 100760 375352
rect 100812 375340 100818 375352
rect 213914 375340 213920 375352
rect 100812 375312 213920 375340
rect 100812 375300 100818 375312
rect 213914 375300 213920 375312
rect 213972 375300 213978 375352
rect 214926 375300 214932 375352
rect 214984 375340 214990 375352
rect 215570 375340 215576 375352
rect 214984 375312 215576 375340
rect 214984 375300 214990 375312
rect 215570 375300 215576 375312
rect 215628 375340 215634 375352
rect 262766 375340 262772 375352
rect 215628 375312 262772 375340
rect 215628 375300 215634 375312
rect 262766 375300 262772 375312
rect 262824 375300 262830 375352
rect 375926 375300 375932 375352
rect 375984 375340 375990 375352
rect 376754 375340 376760 375352
rect 375984 375312 376760 375340
rect 375984 375300 375990 375312
rect 376754 375300 376760 375312
rect 376812 375340 376818 375352
rect 422570 375340 422576 375352
rect 376812 375312 422576 375340
rect 376812 375300 376818 375312
rect 422570 375300 422576 375312
rect 422628 375300 422634 375352
rect 199378 375232 199384 375284
rect 199436 375272 199442 375284
rect 199562 375272 199568 375284
rect 199436 375244 199568 375272
rect 199436 375232 199442 375244
rect 199562 375232 199568 375244
rect 199620 375232 199626 375284
rect 216674 375232 216680 375284
rect 216732 375272 216738 375284
rect 263870 375272 263876 375284
rect 216732 375244 263876 375272
rect 216732 375232 216738 375244
rect 263870 375232 263876 375244
rect 263928 375232 263934 375284
rect 372430 375232 372436 375284
rect 372488 375272 372494 375284
rect 378134 375272 378140 375284
rect 372488 375244 378140 375272
rect 372488 375232 372494 375244
rect 378134 375232 378140 375244
rect 378192 375232 378198 375284
rect 379238 375232 379244 375284
rect 379296 375272 379302 375284
rect 423950 375272 423956 375284
rect 379296 375244 423956 375272
rect 379296 375232 379302 375244
rect 423950 375232 423956 375244
rect 424008 375232 424014 375284
rect 367462 375164 367468 375216
rect 367520 375204 367526 375216
rect 377214 375204 377220 375216
rect 367520 375176 377220 375204
rect 367520 375164 367526 375176
rect 377214 375164 377220 375176
rect 377272 375204 377278 375216
rect 409966 375204 409972 375216
rect 377272 375176 409972 375204
rect 377272 375164 377278 375176
rect 409966 375164 409972 375176
rect 410024 375164 410030 375216
rect 370222 375096 370228 375148
rect 370280 375136 370286 375148
rect 377030 375136 377036 375148
rect 370280 375108 377036 375136
rect 370280 375096 370286 375108
rect 377030 375096 377036 375108
rect 377088 375096 377094 375148
rect 377122 375096 377128 375148
rect 377180 375136 377186 375148
rect 415854 375136 415860 375148
rect 377180 375108 415860 375136
rect 377180 375096 377186 375108
rect 415854 375096 415860 375108
rect 415912 375096 415918 375148
rect 368198 375028 368204 375080
rect 368256 375068 368262 375080
rect 378686 375068 378692 375080
rect 368256 375040 378692 375068
rect 368256 375028 368262 375040
rect 378686 375028 378692 375040
rect 378744 375068 378750 375080
rect 419350 375068 419356 375080
rect 378744 375040 419356 375068
rect 378744 375028 378750 375040
rect 419350 375028 419356 375040
rect 419408 375028 419414 375080
rect 365622 374960 365628 375012
rect 365680 375000 365686 375012
rect 376570 375000 376576 375012
rect 365680 374972 376576 375000
rect 365680 374960 365686 374972
rect 376570 374960 376576 374972
rect 376628 375000 376634 375012
rect 418154 375000 418160 375012
rect 376628 374972 418160 375000
rect 376628 374960 376634 374972
rect 418154 374960 418160 374972
rect 418212 374960 418218 375012
rect 206554 374892 206560 374944
rect 206612 374932 206618 374944
rect 219802 374932 219808 374944
rect 206612 374904 219808 374932
rect 206612 374892 206618 374904
rect 219802 374892 219808 374904
rect 219860 374932 219866 374944
rect 220630 374932 220636 374944
rect 219860 374904 220636 374932
rect 219860 374892 219866 374904
rect 220630 374892 220636 374904
rect 220688 374892 220694 374944
rect 374454 374932 374460 374944
rect 373966 374904 374460 374932
rect 215846 374824 215852 374876
rect 215904 374864 215910 374876
rect 260558 374864 260564 374876
rect 215904 374836 260564 374864
rect 215904 374824 215910 374836
rect 260558 374824 260564 374836
rect 260616 374824 260622 374876
rect 362678 374824 362684 374876
rect 362736 374864 362742 374876
rect 373966 374864 373994 374904
rect 374454 374892 374460 374904
rect 374512 374932 374518 374944
rect 416958 374932 416964 374944
rect 374512 374904 416964 374932
rect 374512 374892 374518 374904
rect 416958 374892 416964 374904
rect 417016 374892 417022 374944
rect 362736 374836 373994 374864
rect 362736 374824 362742 374836
rect 377030 374824 377036 374876
rect 377088 374864 377094 374876
rect 425146 374864 425152 374876
rect 377088 374836 425152 374864
rect 377088 374824 377094 374836
rect 425146 374824 425152 374836
rect 425204 374824 425210 374876
rect 206186 374756 206192 374808
rect 206244 374796 206250 374808
rect 216030 374796 216036 374808
rect 206244 374768 216036 374796
rect 206244 374756 206250 374768
rect 216030 374756 216036 374768
rect 216088 374796 216094 374808
rect 262214 374796 262220 374808
rect 216088 374768 262220 374796
rect 216088 374756 216094 374768
rect 262214 374756 262220 374768
rect 262272 374756 262278 374808
rect 357250 374756 357256 374808
rect 357308 374796 357314 374808
rect 357308 374768 359780 374796
rect 357308 374756 357314 374768
rect 102962 374688 102968 374740
rect 103020 374728 103026 374740
rect 214926 374728 214932 374740
rect 103020 374700 214932 374728
rect 103020 374688 103026 374700
rect 214926 374688 214932 374700
rect 214984 374688 214990 374740
rect 220630 374688 220636 374740
rect 220688 374728 220694 374740
rect 266446 374728 266452 374740
rect 220688 374700 266452 374728
rect 220688 374688 220694 374700
rect 266446 374688 266452 374700
rect 266504 374688 266510 374740
rect 358998 374728 359004 374740
rect 354646 374700 359004 374728
rect 199378 374620 199384 374672
rect 199436 374660 199442 374672
rect 354646 374660 354674 374700
rect 358998 374688 359004 374700
rect 359056 374728 359062 374740
rect 359642 374728 359648 374740
rect 359056 374700 359648 374728
rect 359056 374688 359062 374700
rect 359642 374688 359648 374700
rect 359700 374688 359706 374740
rect 359752 374728 359780 374768
rect 361390 374756 361396 374808
rect 361448 374796 361454 374808
rect 377122 374796 377128 374808
rect 361448 374768 377128 374796
rect 361448 374756 361454 374768
rect 377122 374756 377128 374768
rect 377180 374756 377186 374808
rect 378134 374756 378140 374808
rect 378192 374796 378198 374808
rect 426434 374796 426440 374808
rect 378192 374768 426440 374796
rect 378192 374756 378198 374768
rect 426434 374756 426440 374768
rect 426492 374756 426498 374808
rect 367002 374728 367008 374740
rect 359752 374700 367008 374728
rect 367002 374688 367008 374700
rect 367060 374728 367066 374740
rect 428274 374728 428280 374740
rect 367060 374700 428280 374728
rect 367060 374688 367066 374700
rect 428274 374688 428280 374700
rect 428332 374688 428338 374740
rect 199436 374632 354674 374660
rect 199436 374620 199442 374632
rect 362862 374620 362868 374672
rect 362920 374660 362926 374672
rect 370958 374660 370964 374672
rect 362920 374632 370964 374660
rect 362920 374620 362926 374632
rect 370958 374620 370964 374632
rect 371016 374660 371022 374672
rect 432230 374660 432236 374672
rect 371016 374632 432236 374660
rect 371016 374620 371022 374632
rect 432230 374620 432236 374632
rect 432288 374620 432294 374672
rect 213914 374280 213920 374332
rect 213972 374320 213978 374332
rect 215846 374320 215852 374332
rect 213972 374292 215852 374320
rect 213972 374280 213978 374292
rect 215846 374280 215852 374292
rect 215904 374280 215910 374332
rect 359826 373260 359832 373312
rect 359884 373300 359890 373312
rect 519262 373300 519268 373312
rect 359884 373272 519268 373300
rect 359884 373260 359890 373272
rect 519262 373260 519268 373272
rect 519320 373260 519326 373312
rect 359458 372580 359464 372632
rect 359516 372620 359522 372632
rect 359826 372620 359832 372632
rect 359516 372592 359832 372620
rect 359516 372580 359522 372592
rect 359826 372580 359832 372592
rect 359884 372580 359890 372632
rect 519262 372580 519268 372632
rect 519320 372620 519326 372632
rect 519630 372620 519636 372632
rect 519320 372592 519636 372620
rect 519320 372580 519326 372592
rect 519630 372580 519636 372592
rect 519688 372580 519694 372632
rect 199562 371152 199568 371204
rect 199620 371192 199626 371204
rect 199746 371192 199752 371204
rect 199620 371164 199752 371192
rect 199620 371152 199626 371164
rect 199746 371152 199752 371164
rect 199804 371192 199810 371204
rect 208486 371192 208492 371204
rect 199804 371164 208492 371192
rect 199804 371152 199810 371164
rect 208486 371152 208492 371164
rect 208544 371192 208550 371204
rect 359090 371192 359096 371204
rect 208544 371164 359096 371192
rect 208544 371152 208550 371164
rect 359090 371152 359096 371164
rect 359148 371152 359154 371204
rect 359734 370472 359740 370524
rect 359792 370512 359798 370524
rect 519170 370512 519176 370524
rect 359792 370484 519176 370512
rect 359792 370472 359798 370484
rect 519170 370472 519176 370484
rect 519228 370512 519234 370524
rect 519538 370512 519544 370524
rect 519228 370484 519544 370512
rect 519228 370472 519234 370484
rect 519538 370472 519544 370484
rect 519596 370472 519602 370524
rect 359090 369180 359096 369232
rect 359148 369220 359154 369232
rect 359550 369220 359556 369232
rect 359148 369192 359556 369220
rect 359148 369180 359154 369192
rect 359550 369180 359556 369192
rect 359608 369220 359614 369232
rect 519354 369220 519360 369232
rect 359608 369192 519360 369220
rect 359608 369180 359614 369192
rect 519354 369180 519360 369192
rect 519412 369180 519418 369232
rect 199470 369112 199476 369164
rect 199528 369152 199534 369164
rect 358906 369152 358912 369164
rect 199528 369124 358912 369152
rect 199528 369112 199534 369124
rect 358906 369112 358912 369124
rect 358964 369152 358970 369164
rect 359734 369152 359740 369164
rect 358964 369124 359740 369152
rect 358964 369112 358970 369124
rect 359734 369112 359740 369124
rect 359792 369112 359798 369164
rect 182910 367752 182916 367804
rect 182968 367792 182974 367804
rect 201586 367792 201592 367804
rect 182968 367764 201592 367792
rect 182968 367752 182974 367764
rect 201586 367752 201592 367764
rect 201644 367792 201650 367804
rect 342898 367792 342904 367804
rect 201644 367764 342904 367792
rect 201644 367752 201650 367764
rect 342898 367752 342904 367764
rect 342956 367752 342962 367804
rect 379238 365032 379244 365084
rect 379296 365072 379302 365084
rect 379422 365072 379428 365084
rect 379296 365044 379428 365072
rect 379296 365032 379302 365044
rect 379422 365032 379428 365044
rect 379480 365032 379486 365084
rect 359642 364964 359648 365016
rect 359700 365004 359706 365016
rect 518986 365004 518992 365016
rect 359700 364976 518992 365004
rect 359700 364964 359706 364976
rect 518986 364964 518992 364976
rect 519044 364964 519050 365016
rect 199654 363604 199660 363656
rect 199712 363644 199718 363656
rect 199712 363616 354674 363644
rect 199712 363604 199718 363616
rect 354646 363508 354674 363616
rect 359182 363508 359188 363520
rect 354646 363480 359188 363508
rect 359182 363468 359188 363480
rect 359240 363508 359246 363520
rect 359918 363508 359924 363520
rect 359240 363480 359924 363508
rect 359240 363468 359246 363480
rect 359918 363468 359924 363480
rect 359976 363468 359982 363520
rect 199746 362176 199752 362228
rect 199804 362216 199810 362228
rect 359458 362216 359464 362228
rect 199804 362188 359464 362216
rect 199804 362176 199810 362188
rect 359458 362176 359464 362188
rect 359516 362176 359522 362228
rect 359274 361564 359280 361616
rect 359332 361604 359338 361616
rect 359458 361604 359464 361616
rect 359332 361576 359464 361604
rect 359332 361564 359338 361576
rect 359458 361564 359464 361576
rect 359516 361564 359522 361616
rect 202782 360816 202788 360868
rect 202840 360856 202846 360868
rect 210418 360856 210424 360868
rect 202840 360828 210424 360856
rect 202840 360816 202846 360828
rect 210418 360816 210424 360828
rect 210476 360816 210482 360868
rect 197538 360136 197544 360188
rect 197596 360176 197602 360188
rect 201770 360176 201776 360188
rect 197596 360148 201776 360176
rect 197596 360136 197602 360148
rect 201770 360136 201776 360148
rect 201828 360136 201834 360188
rect 500770 359660 500776 359712
rect 500828 359700 500834 359712
rect 518066 359700 518072 359712
rect 500828 359672 518072 359700
rect 500828 359660 500834 359672
rect 518066 359660 518072 359672
rect 518124 359660 518130 359712
rect 498838 359592 498844 359644
rect 498896 359632 498902 359644
rect 517974 359632 517980 359644
rect 498896 359604 517980 359632
rect 498896 359592 498902 359604
rect 517974 359592 517980 359604
rect 518032 359592 518038 359644
rect 197722 359524 197728 359576
rect 197780 359564 197786 359576
rect 204530 359564 204536 359576
rect 197780 359536 204536 359564
rect 197780 359524 197786 359536
rect 204530 359524 204536 359536
rect 204588 359524 204594 359576
rect 277302 359524 277308 359576
rect 277360 359564 277366 359576
rect 357434 359564 357440 359576
rect 277360 359536 357440 359564
rect 277360 359524 277366 359536
rect 357434 359524 357440 359536
rect 357492 359524 357498 359576
rect 438118 359524 438124 359576
rect 438176 359564 438182 359576
rect 516594 359564 516600 359576
rect 438176 359536 516600 359564
rect 438176 359524 438182 359536
rect 516594 359524 516600 359536
rect 516652 359524 516658 359576
rect 190914 359456 190920 359508
rect 190972 359496 190978 359508
rect 201494 359496 201500 359508
rect 190972 359468 201500 359496
rect 190972 359456 190978 359468
rect 201494 359456 201500 359468
rect 201552 359496 201558 359508
rect 202782 359496 202788 359508
rect 201552 359468 202788 359496
rect 201552 359456 201558 359468
rect 202782 359456 202788 359468
rect 202840 359456 202846 359508
rect 351730 359456 351736 359508
rect 351788 359496 351794 359508
rect 358078 359496 358084 359508
rect 351788 359468 358084 359496
rect 351788 359456 351794 359468
rect 358078 359456 358084 359468
rect 358136 359456 358142 359508
rect 360286 359252 360292 359304
rect 360344 359292 360350 359304
rect 361574 359292 361580 359304
rect 360344 359264 361580 359292
rect 360344 359252 360350 359264
rect 361574 359252 361580 359264
rect 361632 359252 361638 359304
rect 342254 358912 342260 358964
rect 342312 358952 342318 358964
rect 343542 358952 343548 358964
rect 342312 358924 343548 358952
rect 342312 358912 342318 358924
rect 343542 358912 343548 358924
rect 343600 358952 343606 358964
rect 359090 358952 359096 358964
rect 343600 358924 359096 358952
rect 343600 358912 343606 358924
rect 359090 358912 359096 358924
rect 359148 358912 359154 358964
rect 179690 358844 179696 358896
rect 179748 358884 179754 358896
rect 197538 358884 197544 358896
rect 179748 358856 197544 358884
rect 179748 358844 179754 358856
rect 197538 358844 197544 358856
rect 197596 358844 197602 358896
rect 339770 358844 339776 358896
rect 339828 358884 339834 358896
rect 357342 358884 357348 358896
rect 339828 358856 357348 358884
rect 339828 358844 339834 358856
rect 357342 358844 357348 358856
rect 357400 358884 357406 358896
rect 362954 358884 362960 358896
rect 357400 358856 362960 358884
rect 357400 358844 357406 358856
rect 362954 358844 362960 358856
rect 363012 358844 363018 358896
rect 178586 358776 178592 358828
rect 178644 358816 178650 358828
rect 197722 358816 197728 358828
rect 178644 358788 197728 358816
rect 178644 358776 178650 358788
rect 197722 358776 197728 358788
rect 197780 358776 197786 358828
rect 338482 358776 338488 358828
rect 338540 358816 338546 358828
rect 360286 358816 360292 358828
rect 338540 358788 360292 358816
rect 338540 358776 338546 358788
rect 360286 358776 360292 358788
rect 360344 358776 360350 358828
rect 510890 358776 510896 358828
rect 510948 358816 510954 358828
rect 511902 358816 511908 358828
rect 510948 358788 511908 358816
rect 510948 358776 510954 358788
rect 511902 358776 511908 358788
rect 511960 358816 511966 358828
rect 517514 358816 517520 358828
rect 511960 358788 517520 358816
rect 511960 358776 511966 358788
rect 517514 358776 517520 358788
rect 517572 358776 517578 358828
rect 3326 358708 3332 358760
rect 3384 358748 3390 358760
rect 18598 358748 18604 358760
rect 3384 358720 18604 358748
rect 3384 358708 3390 358720
rect 18598 358708 18604 358720
rect 18656 358708 18662 358760
rect 218514 358708 218520 358760
rect 218572 358748 218578 358760
rect 220814 358748 220820 358760
rect 218572 358720 220820 358748
rect 218572 358708 218578 358720
rect 220814 358708 220820 358720
rect 220872 358708 220878 358760
rect 379422 358708 379428 358760
rect 379480 358748 379486 358760
rect 380894 358748 380900 358760
rect 379480 358720 380900 358748
rect 379480 358708 379486 358720
rect 380894 358708 380900 358720
rect 380952 358708 380958 358760
rect 218606 358436 218612 358488
rect 218664 358476 218670 358488
rect 221090 358476 221096 358488
rect 218664 358448 221096 358476
rect 218664 358436 218670 358448
rect 221090 358436 221096 358448
rect 221148 358436 221154 358488
rect 375926 358368 375932 358420
rect 375984 358408 375990 358420
rect 381262 358408 381268 358420
rect 375984 358380 381268 358408
rect 375984 358368 375990 358380
rect 381262 358368 381268 358380
rect 381320 358368 381326 358420
rect 217226 358232 217232 358284
rect 217284 358272 217290 358284
rect 220998 358272 221004 358284
rect 217284 358244 221004 358272
rect 217284 358232 217290 358244
rect 220998 358232 221004 358244
rect 221056 358232 221062 358284
rect 373166 358096 373172 358148
rect 373224 358136 373230 358148
rect 381170 358136 381176 358148
rect 373224 358108 381176 358136
rect 373224 358096 373230 358108
rect 381170 358096 381176 358108
rect 381228 358096 381234 358148
rect 182818 358028 182824 358080
rect 182876 358068 182882 358080
rect 197722 358068 197728 358080
rect 182876 358040 197728 358068
rect 182876 358028 182882 358040
rect 197722 358028 197728 358040
rect 197780 358068 197786 358080
rect 342254 358068 342260 358080
rect 197780 358040 342260 358068
rect 197780 358028 197786 358040
rect 342254 358028 342260 358040
rect 342312 358028 342318 358080
rect 372430 358028 372436 358080
rect 372488 358068 372494 358080
rect 381078 358068 381084 358080
rect 372488 358040 381084 358068
rect 372488 358028 372494 358040
rect 381078 358028 381084 358040
rect 381136 358028 381142 358080
rect 214466 357620 214472 357672
rect 214524 357660 214530 357672
rect 220906 357660 220912 357672
rect 214524 357632 220912 357660
rect 214524 357620 214530 357632
rect 220906 357620 220912 357632
rect 220964 357620 220970 357672
rect 379330 357484 379336 357536
rect 379388 357524 379394 357536
rect 380986 357524 380992 357536
rect 379388 357496 380992 357524
rect 379388 357484 379394 357496
rect 380986 357484 380992 357496
rect 381044 357484 381050 357536
rect 55766 357348 55772 357400
rect 55824 357388 55830 357400
rect 60734 357388 60740 357400
rect 55824 357360 60740 357388
rect 55824 357348 55830 357360
rect 60734 357348 60740 357360
rect 60792 357348 60798 357400
rect 58618 355988 58624 356040
rect 58676 356028 58682 356040
rect 59630 356028 59636 356040
rect 58676 356000 59636 356028
rect 58676 355988 58682 356000
rect 59630 355988 59636 356000
rect 59688 355988 59694 356040
rect 518158 353200 518164 353252
rect 518216 353240 518222 353252
rect 580166 353240 580172 353252
rect 518216 353212 580172 353240
rect 518216 353200 518222 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 46290 300772 46296 300824
rect 46348 300812 46354 300824
rect 56962 300812 56968 300824
rect 46348 300784 56968 300812
rect 46348 300772 46354 300784
rect 56962 300772 56968 300784
rect 57020 300772 57026 300824
rect 57054 300772 57060 300824
rect 57112 300812 57118 300824
rect 58526 300812 58532 300824
rect 57112 300784 58532 300812
rect 57112 300772 57118 300784
rect 58526 300772 58532 300784
rect 58584 300772 58590 300824
rect 520182 288396 520188 288448
rect 520240 288436 520246 288448
rect 580258 288436 580264 288448
rect 520240 288408 580264 288436
rect 520240 288396 520246 288408
rect 580258 288396 580264 288408
rect 580316 288396 580322 288448
rect 519170 287036 519176 287088
rect 519228 287076 519234 287088
rect 519630 287076 519636 287088
rect 519228 287048 519636 287076
rect 519228 287036 519234 287048
rect 519630 287036 519636 287048
rect 519688 287076 519694 287088
rect 580350 287076 580356 287088
rect 519688 287048 580356 287076
rect 519688 287036 519694 287048
rect 580350 287036 580356 287048
rect 580408 287036 580414 287088
rect 200758 284248 200764 284300
rect 200816 284288 200822 284300
rect 216674 284288 216680 284300
rect 200816 284260 216680 284288
rect 200816 284248 200822 284260
rect 216674 284248 216680 284260
rect 216732 284248 216738 284300
rect 358630 284248 358636 284300
rect 358688 284288 358694 284300
rect 376938 284288 376944 284300
rect 358688 284260 376944 284288
rect 358688 284248 358694 284260
rect 376938 284248 376944 284260
rect 376996 284248 377002 284300
rect 201494 282820 201500 282872
rect 201552 282860 201558 282872
rect 216674 282860 216680 282872
rect 201552 282832 216680 282860
rect 201552 282820 201558 282832
rect 216674 282820 216680 282832
rect 216732 282820 216738 282872
rect 361298 282820 361304 282872
rect 361356 282860 361362 282872
rect 376754 282860 376760 282872
rect 361356 282832 376760 282860
rect 361356 282820 361362 282832
rect 376754 282820 376760 282832
rect 376812 282820 376818 282872
rect 203886 282752 203892 282804
rect 203944 282792 203950 282804
rect 216766 282792 216772 282804
rect 203944 282764 216772 282792
rect 203944 282752 203950 282764
rect 216766 282752 216772 282764
rect 216824 282752 216830 282804
rect 200758 282412 200764 282464
rect 200816 282452 200822 282464
rect 201494 282452 201500 282464
rect 200816 282424 201500 282452
rect 200816 282412 200822 282424
rect 201494 282412 201500 282424
rect 201552 282412 201558 282464
rect 54478 282140 54484 282192
rect 54536 282180 54542 282192
rect 57974 282180 57980 282192
rect 54536 282152 57980 282180
rect 54536 282140 54542 282152
rect 57974 282140 57980 282152
rect 58032 282140 58038 282192
rect 376938 281568 376944 281580
rect 360212 281540 376944 281568
rect 360212 281512 360240 281540
rect 376938 281528 376944 281540
rect 376996 281528 377002 281580
rect 45462 281460 45468 281512
rect 45520 281500 45526 281512
rect 57238 281500 57244 281512
rect 45520 281472 57244 281500
rect 45520 281460 45526 281472
rect 57238 281460 57244 281472
rect 57296 281500 57302 281512
rect 57514 281500 57520 281512
rect 57296 281472 57520 281500
rect 57296 281460 57302 281472
rect 57514 281460 57520 281472
rect 57572 281460 57578 281512
rect 358078 281460 358084 281512
rect 358136 281500 358142 281512
rect 360194 281500 360200 281512
rect 358136 281472 360200 281500
rect 358136 281460 358142 281472
rect 360194 281460 360200 281472
rect 360252 281460 360258 281512
rect 45278 273640 45284 273692
rect 45336 273680 45342 273692
rect 145926 273680 145932 273692
rect 45336 273652 145932 273680
rect 45336 273640 45342 273652
rect 145926 273640 145932 273652
rect 145984 273640 145990 273692
rect 42610 273572 42616 273624
rect 42668 273612 42674 273624
rect 131022 273612 131028 273624
rect 42668 273584 131028 273612
rect 42668 273572 42674 273584
rect 131022 273572 131028 273584
rect 131080 273572 131086 273624
rect 372522 273572 372528 273624
rect 372580 273612 372586 273624
rect 379238 273612 379244 273624
rect 372580 273584 379244 273612
rect 372580 273572 372586 273584
rect 379238 273572 379244 273584
rect 379296 273572 379302 273624
rect 43346 273504 43352 273556
rect 43404 273544 43410 273556
rect 133414 273544 133420 273556
rect 43404 273516 133420 273544
rect 43404 273504 43410 273516
rect 133414 273504 133420 273516
rect 133472 273504 133478 273556
rect 369026 273504 369032 273556
rect 369084 273544 369090 273556
rect 378134 273544 378140 273556
rect 369084 273516 378140 273544
rect 369084 273504 369090 273516
rect 378134 273504 378140 273516
rect 378192 273544 378198 273556
rect 378594 273544 378600 273556
rect 378192 273516 378600 273544
rect 378192 273504 378198 273516
rect 378594 273504 378600 273516
rect 378652 273504 378658 273556
rect 379422 273504 379428 273556
rect 379480 273544 379486 273556
rect 379790 273544 379796 273556
rect 379480 273516 379796 273544
rect 379480 273504 379486 273516
rect 379790 273504 379796 273516
rect 379848 273544 379854 273556
rect 427630 273544 427636 273556
rect 379848 273516 427636 273544
rect 379848 273504 379854 273516
rect 427630 273504 427636 273516
rect 427688 273504 427694 273556
rect 45186 273436 45192 273488
rect 45244 273476 45250 273488
rect 135898 273476 135904 273488
rect 45244 273448 135904 273476
rect 45244 273436 45250 273448
rect 135898 273436 135904 273448
rect 135956 273436 135962 273488
rect 212074 273436 212080 273488
rect 212132 273476 212138 273488
rect 250714 273476 250720 273488
rect 212132 273448 250720 273476
rect 212132 273436 212138 273448
rect 250714 273436 250720 273448
rect 250772 273436 250778 273488
rect 361206 273436 361212 273488
rect 361264 273476 361270 273488
rect 416038 273476 416044 273488
rect 361264 273448 416044 273476
rect 361264 273436 361270 273448
rect 416038 273436 416044 273448
rect 416096 273436 416102 273488
rect 45002 273368 45008 273420
rect 45060 273408 45066 273420
rect 138474 273408 138480 273420
rect 45060 273380 138480 273408
rect 45060 273368 45066 273380
rect 138474 273368 138480 273380
rect 138532 273368 138538 273420
rect 211706 273368 211712 273420
rect 211764 273408 211770 273420
rect 272242 273408 272248 273420
rect 211764 273380 272248 273408
rect 211764 273368 211770 273380
rect 272242 273368 272248 273380
rect 272300 273368 272306 273420
rect 373166 273368 373172 273420
rect 373224 273408 373230 273420
rect 433334 273408 433340 273420
rect 373224 273380 433340 273408
rect 373224 273368 373230 273380
rect 433334 273368 433340 273380
rect 433392 273368 433398 273420
rect 45094 273300 45100 273352
rect 45152 273340 45158 273352
rect 140866 273340 140872 273352
rect 45152 273312 140872 273340
rect 45152 273300 45158 273312
rect 140866 273300 140872 273312
rect 140924 273300 140930 273352
rect 212810 273300 212816 273352
rect 212868 273340 212874 273352
rect 273254 273340 273260 273352
rect 212868 273312 273260 273340
rect 212868 273300 212874 273312
rect 273254 273300 273260 273312
rect 273312 273300 273318 273352
rect 368106 273300 368112 273352
rect 368164 273340 368170 273352
rect 440878 273340 440884 273352
rect 368164 273312 440884 273340
rect 368164 273300 368170 273312
rect 440878 273300 440884 273312
rect 440936 273300 440942 273352
rect 52362 273232 52368 273284
rect 52420 273272 52426 273284
rect 57974 273272 57980 273284
rect 52420 273244 57980 273272
rect 52420 273232 52426 273244
rect 57974 273232 57980 273244
rect 58032 273272 58038 273284
rect 58802 273272 58808 273284
rect 58032 273244 58808 273272
rect 58032 273232 58038 273244
rect 58802 273232 58808 273244
rect 58860 273232 58866 273284
rect 64846 273244 77248 273272
rect 50522 272960 50528 273012
rect 50580 273000 50586 273012
rect 53834 273000 53840 273012
rect 50580 272972 53840 273000
rect 50580 272960 50586 272972
rect 53834 272960 53840 272972
rect 53892 272960 53898 273012
rect 46474 272892 46480 272944
rect 46532 272932 46538 272944
rect 50982 272932 50988 272944
rect 46532 272904 50988 272932
rect 46532 272892 46538 272904
rect 50982 272892 50988 272904
rect 51040 272932 51046 272944
rect 64846 272932 64874 273244
rect 77220 273204 77248 273244
rect 207842 273232 207848 273284
rect 207900 273272 207906 273284
rect 280890 273272 280896 273284
rect 207900 273244 280896 273272
rect 207900 273232 207906 273244
rect 280890 273232 280896 273244
rect 280948 273232 280954 273284
rect 358446 273232 358452 273284
rect 358504 273272 358510 273284
rect 430942 273272 430948 273284
rect 358504 273244 430948 273272
rect 358504 273232 358510 273244
rect 430942 273232 430948 273244
rect 431000 273232 431006 273284
rect 77220 273176 84194 273204
rect 51040 272904 64874 272932
rect 84166 272932 84194 273176
rect 374454 273164 374460 273216
rect 374512 273204 374518 273216
rect 396718 273204 396724 273216
rect 374512 273176 396724 273204
rect 374512 273164 374518 273176
rect 396718 273164 396724 273176
rect 396776 273164 396782 273216
rect 379238 273096 379244 273148
rect 379296 273136 379302 273148
rect 423766 273136 423772 273148
rect 379296 273108 423772 273136
rect 379296 273096 379302 273108
rect 423766 273096 423772 273108
rect 423824 273096 423830 273148
rect 378594 273028 378600 273080
rect 378652 273068 378658 273080
rect 426434 273068 426440 273080
rect 378652 273040 426440 273068
rect 378652 273028 378658 273040
rect 426434 273028 426440 273040
rect 426492 273028 426498 273080
rect 366818 272960 366824 273012
rect 366876 273000 366882 273012
rect 423398 273000 423404 273012
rect 366876 272972 423404 273000
rect 366876 272960 366882 272972
rect 423398 272960 423404 272972
rect 423456 272960 423462 273012
rect 98086 272932 98092 272944
rect 84166 272904 98092 272932
rect 51040 272892 51046 272904
rect 98086 272892 98092 272904
rect 98144 272892 98150 272944
rect 356882 272892 356888 272944
rect 356940 272932 356946 272944
rect 428182 272932 428188 272944
rect 356940 272904 428188 272932
rect 356940 272892 356946 272904
rect 428182 272892 428188 272904
rect 428240 272892 428246 272944
rect 54846 272824 54852 272876
rect 54904 272864 54910 272876
rect 88334 272864 88340 272876
rect 54904 272836 88340 272864
rect 54904 272824 54910 272836
rect 88334 272824 88340 272836
rect 88392 272824 88398 272876
rect 210878 272824 210884 272876
rect 210936 272864 210942 272876
rect 283374 272864 283380 272876
rect 210936 272836 283380 272864
rect 210936 272824 210942 272836
rect 283374 272824 283380 272836
rect 283432 272824 283438 272876
rect 369486 272824 369492 272876
rect 369544 272864 369550 272876
rect 468478 272864 468484 272876
rect 369544 272836 468484 272864
rect 369544 272824 369550 272836
rect 468478 272824 468484 272836
rect 468536 272824 468542 272876
rect 58802 272756 58808 272808
rect 58860 272796 58866 272808
rect 99374 272796 99380 272808
rect 58860 272768 99380 272796
rect 58860 272756 58866 272768
rect 99374 272756 99380 272768
rect 99432 272756 99438 272808
rect 216122 272756 216128 272808
rect 216180 272796 216186 272808
rect 295886 272796 295892 272808
rect 216180 272768 295892 272796
rect 216180 272756 216186 272768
rect 295886 272756 295892 272768
rect 295944 272756 295950 272808
rect 372154 272756 372160 272808
rect 372212 272796 372218 272808
rect 470870 272796 470876 272808
rect 372212 272768 470876 272796
rect 372212 272756 372218 272768
rect 470870 272756 470876 272768
rect 470928 272756 470934 272808
rect 49050 272688 49056 272740
rect 49108 272728 49114 272740
rect 90726 272728 90732 272740
rect 49108 272700 90732 272728
rect 49108 272688 49114 272700
rect 90726 272688 90732 272700
rect 90784 272688 90790 272740
rect 209590 272688 209596 272740
rect 209648 272728 209654 272740
rect 290918 272728 290924 272740
rect 209648 272700 290924 272728
rect 209648 272688 209654 272700
rect 290918 272688 290924 272700
rect 290976 272688 290982 272740
rect 373718 272688 373724 272740
rect 373776 272728 373782 272740
rect 478414 272728 478420 272740
rect 373776 272700 478420 272728
rect 373776 272688 373782 272700
rect 478414 272688 478420 272700
rect 478472 272688 478478 272740
rect 50430 272620 50436 272672
rect 50488 272660 50494 272672
rect 93670 272660 93676 272672
rect 50488 272632 93676 272660
rect 50488 272620 50494 272632
rect 93670 272620 93676 272632
rect 93728 272620 93734 272672
rect 203794 272620 203800 272672
rect 203852 272660 203858 272672
rect 288158 272660 288164 272672
rect 203852 272632 288164 272660
rect 203852 272620 203858 272632
rect 288158 272620 288164 272632
rect 288216 272620 288222 272672
rect 376294 272620 376300 272672
rect 376352 272660 376358 272672
rect 480806 272660 480812 272672
rect 376352 272632 480812 272660
rect 376352 272620 376358 272632
rect 480806 272620 480812 272632
rect 480864 272620 480870 272672
rect 51810 272552 51816 272604
rect 51868 272592 51874 272604
rect 98454 272592 98460 272604
rect 51868 272564 98460 272592
rect 51868 272552 51874 272564
rect 98454 272552 98460 272564
rect 98512 272552 98518 272604
rect 205174 272552 205180 272604
rect 205232 272592 205238 272604
rect 298462 272592 298468 272604
rect 205232 272564 298468 272592
rect 205232 272552 205238 272564
rect 298462 272552 298468 272564
rect 298520 272552 298526 272604
rect 363966 272552 363972 272604
rect 364024 272592 364030 272604
rect 475838 272592 475844 272604
rect 364024 272564 475844 272592
rect 364024 272552 364030 272564
rect 475838 272552 475844 272564
rect 475896 272552 475902 272604
rect 47946 272484 47952 272536
rect 48004 272524 48010 272536
rect 95878 272524 95884 272536
rect 48004 272496 95884 272524
rect 48004 272484 48010 272496
rect 95878 272484 95884 272496
rect 95936 272484 95942 272536
rect 200942 272484 200948 272536
rect 201000 272524 201006 272536
rect 300854 272524 300860 272536
rect 201000 272496 300860 272524
rect 201000 272484 201006 272496
rect 300854 272484 300860 272496
rect 300912 272484 300918 272536
rect 362586 272484 362592 272536
rect 362644 272524 362650 272536
rect 473446 272524 473452 272536
rect 362644 272496 473452 272524
rect 362644 272484 362650 272496
rect 473446 272484 473452 272496
rect 473504 272484 473510 272536
rect 55766 272416 55772 272468
rect 55824 272456 55830 272468
rect 59630 272456 59636 272468
rect 55824 272428 59636 272456
rect 55824 272416 55830 272428
rect 59630 272416 59636 272428
rect 59688 272416 59694 272468
rect 59722 272416 59728 272468
rect 59780 272456 59786 272468
rect 60826 272456 60832 272468
rect 59780 272428 60832 272456
rect 59780 272416 59786 272428
rect 60826 272416 60832 272428
rect 60884 272416 60890 272468
rect 48038 272348 48044 272400
rect 48096 272388 48102 272400
rect 77110 272388 77116 272400
rect 48096 272360 77116 272388
rect 48096 272348 48102 272360
rect 77110 272348 77116 272360
rect 77168 272348 77174 272400
rect 377030 272348 377036 272400
rect 377088 272388 377094 272400
rect 379698 272388 379704 272400
rect 377088 272360 379704 272388
rect 377088 272348 377094 272360
rect 379698 272348 379704 272360
rect 379756 272348 379762 272400
rect 48958 272280 48964 272332
rect 49016 272320 49022 272332
rect 54294 272320 54300 272332
rect 49016 272292 54300 272320
rect 49016 272280 49022 272292
rect 54294 272280 54300 272292
rect 54352 272320 54358 272332
rect 82998 272320 83004 272332
rect 54352 272292 83004 272320
rect 54352 272280 54358 272292
rect 82998 272280 83004 272292
rect 83056 272280 83062 272332
rect 374454 272280 374460 272332
rect 374512 272320 374518 272332
rect 375190 272320 375196 272332
rect 374512 272292 375196 272320
rect 374512 272280 374518 272292
rect 375190 272280 375196 272292
rect 375248 272280 375254 272332
rect 67542 272212 67548 272264
rect 67600 272252 67606 272264
rect 95970 272252 95976 272264
rect 67600 272224 95976 272252
rect 67600 272212 67606 272224
rect 95970 272212 95976 272224
rect 96028 272212 96034 272264
rect 53834 272144 53840 272196
rect 53892 272184 53898 272196
rect 54110 272184 54116 272196
rect 53892 272156 54116 272184
rect 53892 272144 53898 272156
rect 54110 272144 54116 272156
rect 54168 272184 54174 272196
rect 85390 272184 85396 272196
rect 54168 272156 85396 272184
rect 54168 272144 54174 272156
rect 85390 272144 85396 272156
rect 85448 272144 85454 272196
rect 46382 272076 46388 272128
rect 46440 272116 46446 272128
rect 75914 272116 75920 272128
rect 46440 272088 75920 272116
rect 46440 272076 46446 272088
rect 75914 272076 75920 272088
rect 75972 272076 75978 272128
rect 60826 272008 60832 272060
rect 60884 272048 60890 272060
rect 94222 272048 94228 272060
rect 60884 272020 94228 272048
rect 60884 272008 60890 272020
rect 94222 272008 94228 272020
rect 94280 272008 94286 272060
rect 379606 272008 379612 272060
rect 379664 272048 379670 272060
rect 380066 272048 380072 272060
rect 379664 272020 380072 272048
rect 379664 272008 379670 272020
rect 380066 272008 380072 272020
rect 380124 272008 380130 272060
rect 54202 271940 54208 271992
rect 54260 271980 54266 271992
rect 54754 271980 54760 271992
rect 54260 271952 54760 271980
rect 54260 271940 54266 271952
rect 54754 271940 54760 271952
rect 54812 271980 54818 271992
rect 88334 271980 88340 271992
rect 54812 271952 88340 271980
rect 54812 271940 54818 271952
rect 88334 271940 88340 271952
rect 88392 271940 88398 271992
rect 379698 271940 379704 271992
rect 379756 271980 379762 271992
rect 425054 271980 425060 271992
rect 379756 271952 425060 271980
rect 379756 271940 379762 271952
rect 425054 271940 425060 271952
rect 425112 271940 425118 271992
rect 58526 271872 58532 271924
rect 58584 271912 58590 271924
rect 102134 271912 102140 271924
rect 58584 271884 102140 271912
rect 58584 271872 58590 271884
rect 102134 271872 102140 271884
rect 102192 271872 102198 271924
rect 213638 271872 213644 271924
rect 213696 271912 213702 271924
rect 215662 271912 215668 271924
rect 213696 271884 215668 271912
rect 213696 271872 213702 271884
rect 215662 271872 215668 271884
rect 215720 271912 215726 271924
rect 235994 271912 236000 271924
rect 215720 271884 236000 271912
rect 215720 271872 215726 271884
rect 235994 271872 236000 271884
rect 236052 271872 236058 271924
rect 359090 271912 359096 271924
rect 356900 271884 359096 271912
rect 45370 271804 45376 271856
rect 45428 271844 45434 271856
rect 143534 271844 143540 271856
rect 45428 271816 143540 271844
rect 45428 271804 45434 271816
rect 143534 271804 143540 271816
rect 143592 271804 143598 271856
rect 154482 271804 154488 271856
rect 154540 271844 154546 271856
rect 200114 271844 200120 271856
rect 154540 271816 200120 271844
rect 154540 271804 154546 271816
rect 200114 271804 200120 271816
rect 200172 271804 200178 271856
rect 212166 271804 212172 271856
rect 212224 271844 212230 271856
rect 307754 271844 307760 271856
rect 212224 271816 307760 271844
rect 212224 271804 212230 271816
rect 307754 271804 307760 271816
rect 307812 271804 307818 271856
rect 125594 271776 125600 271788
rect 45526 271748 125600 271776
rect 43438 271668 43444 271720
rect 43496 271708 43502 271720
rect 45526 271708 45554 271748
rect 125594 271736 125600 271748
rect 125652 271736 125658 271788
rect 157242 271736 157248 271788
rect 157300 271776 157306 271788
rect 201678 271776 201684 271788
rect 157300 271748 201684 271776
rect 157300 271736 157306 271748
rect 201678 271736 201684 271748
rect 201736 271736 201742 271788
rect 219526 271736 219532 271788
rect 219584 271776 219590 271788
rect 219802 271776 219808 271788
rect 219584 271748 219808 271776
rect 219584 271736 219590 271748
rect 219802 271736 219808 271748
rect 219860 271736 219866 271788
rect 223574 271736 223580 271788
rect 223632 271776 223638 271788
rect 302234 271776 302240 271788
rect 223632 271748 302240 271776
rect 223632 271736 223638 271748
rect 302234 271736 302240 271748
rect 302292 271736 302298 271788
rect 43496 271680 45554 271708
rect 43496 271668 43502 271680
rect 47670 271668 47676 271720
rect 47728 271708 47734 271720
rect 47946 271708 47952 271720
rect 47728 271680 47952 271708
rect 47728 271668 47734 271680
rect 47946 271668 47952 271680
rect 48004 271668 48010 271720
rect 107654 271708 107660 271720
rect 50356 271680 107660 271708
rect 41046 271600 41052 271652
rect 41104 271640 41110 271652
rect 50356 271640 50384 271680
rect 107654 271668 107660 271680
rect 107712 271668 107718 271720
rect 158622 271668 158628 271720
rect 158680 271708 158686 271720
rect 197354 271708 197360 271720
rect 158680 271680 197360 271708
rect 158680 271668 158686 271680
rect 197354 271668 197360 271680
rect 197412 271668 197418 271720
rect 200850 271668 200856 271720
rect 200908 271708 200914 271720
rect 270494 271708 270500 271720
rect 200908 271680 270500 271708
rect 200908 271668 200914 271680
rect 270494 271668 270500 271680
rect 270552 271668 270558 271720
rect 41104 271612 50384 271640
rect 41104 271600 41110 271612
rect 54662 271600 54668 271652
rect 54720 271640 54726 271652
rect 120074 271640 120080 271652
rect 54720 271612 120080 271640
rect 54720 271600 54726 271612
rect 120074 271600 120080 271612
rect 120132 271600 120138 271652
rect 202322 271600 202328 271652
rect 202380 271640 202386 271652
rect 264974 271640 264980 271652
rect 202380 271612 264980 271640
rect 202380 271600 202386 271612
rect 264974 271600 264980 271612
rect 265032 271600 265038 271652
rect 46658 271532 46664 271584
rect 46716 271572 46722 271584
rect 52454 271572 52460 271584
rect 46716 271544 52460 271572
rect 46716 271532 46722 271544
rect 52454 271532 52460 271544
rect 52512 271532 52518 271584
rect 56870 271532 56876 271584
rect 56928 271572 56934 271584
rect 123110 271572 123116 271584
rect 56928 271544 123116 271572
rect 56928 271532 56934 271544
rect 123110 271532 123116 271544
rect 123168 271532 123174 271584
rect 164142 271532 164148 271584
rect 164200 271572 164206 271584
rect 197446 271572 197452 271584
rect 164200 271544 197452 271572
rect 164200 271532 164206 271544
rect 197446 271532 197452 271544
rect 197504 271532 197510 271584
rect 203702 271532 203708 271584
rect 203760 271572 203766 271584
rect 263594 271572 263600 271584
rect 203760 271544 263600 271572
rect 203760 271532 203766 271544
rect 263594 271532 263600 271544
rect 263652 271532 263658 271584
rect 343542 271532 343548 271584
rect 343600 271572 343606 271584
rect 356900 271572 356928 271884
rect 359090 271872 359096 271884
rect 359148 271872 359154 271924
rect 370406 271872 370412 271924
rect 370464 271912 370470 271924
rect 427998 271912 428004 271924
rect 370464 271884 428004 271912
rect 370464 271872 370470 271884
rect 427998 271872 428004 271884
rect 428056 271872 428062 271924
rect 440142 271872 440148 271924
rect 440200 271912 440206 271924
rect 516594 271912 516600 271924
rect 440200 271884 516600 271912
rect 440200 271872 440206 271884
rect 516594 271872 516600 271884
rect 516652 271872 516658 271924
rect 368014 271804 368020 271856
rect 368072 271844 368078 271856
rect 458174 271844 458180 271856
rect 368072 271816 458180 271844
rect 368072 271804 368078 271816
rect 458174 271804 458180 271816
rect 458232 271804 458238 271856
rect 366726 271736 366732 271788
rect 366784 271776 366790 271788
rect 455782 271776 455788 271788
rect 366784 271748 455788 271776
rect 366784 271736 366790 271748
rect 455782 271736 455788 271748
rect 455840 271736 455846 271788
rect 362494 271668 362500 271720
rect 362552 271708 362558 271720
rect 449894 271708 449900 271720
rect 362552 271680 449900 271708
rect 362552 271668 362558 271680
rect 449894 271668 449900 271680
rect 449952 271668 449958 271720
rect 367002 271600 367008 271652
rect 367060 271640 367066 271652
rect 370406 271640 370412 271652
rect 367060 271612 370412 271640
rect 367060 271600 367066 271612
rect 370406 271600 370412 271612
rect 370464 271600 370470 271652
rect 376386 271600 376392 271652
rect 376444 271640 376450 271652
rect 460934 271640 460940 271652
rect 376444 271612 460940 271640
rect 376444 271600 376450 271612
rect 460934 271600 460940 271612
rect 460992 271600 460998 271652
rect 357066 271572 357072 271584
rect 343600 271544 357072 271572
rect 343600 271532 343606 271544
rect 357066 271532 357072 271544
rect 357124 271532 357130 271584
rect 369394 271532 369400 271584
rect 369452 271572 369458 271584
rect 452654 271572 452660 271584
rect 369452 271544 452660 271572
rect 369452 271532 369458 271544
rect 452654 271532 452660 271544
rect 452712 271532 452718 271584
rect 53006 271464 53012 271516
rect 53064 271504 53070 271516
rect 117314 271504 117320 271516
rect 53064 271476 117320 271504
rect 53064 271464 53070 271476
rect 117314 271464 117320 271476
rect 117372 271464 117378 271516
rect 161382 271464 161388 271516
rect 161440 271504 161446 271516
rect 202966 271504 202972 271516
rect 161440 271476 202972 271504
rect 161440 271464 161446 271476
rect 202966 271464 202972 271476
rect 203024 271464 203030 271516
rect 216306 271464 216312 271516
rect 216364 271504 216370 271516
rect 276106 271504 276112 271516
rect 216364 271476 276112 271504
rect 216364 271464 216370 271476
rect 276106 271464 276112 271476
rect 276164 271464 276170 271516
rect 365438 271464 365444 271516
rect 365496 271504 365502 271516
rect 442994 271504 443000 271516
rect 365496 271476 443000 271504
rect 365496 271464 365502 271476
rect 442994 271464 443000 271476
rect 443052 271464 443058 271516
rect 46106 271396 46112 271448
rect 46164 271436 46170 271448
rect 46658 271436 46664 271448
rect 46164 271408 46664 271436
rect 46164 271396 46170 271408
rect 46658 271396 46664 271408
rect 46716 271396 46722 271448
rect 52822 271396 52828 271448
rect 52880 271436 52886 271448
rect 115934 271436 115940 271448
rect 52880 271408 115940 271436
rect 52880 271396 52886 271408
rect 115934 271396 115940 271408
rect 115992 271396 115998 271448
rect 197354 271396 197360 271448
rect 197412 271436 197418 271448
rect 197722 271436 197728 271448
rect 197412 271408 197728 271436
rect 197412 271396 197418 271408
rect 197722 271396 197728 271408
rect 197780 271396 197786 271448
rect 216490 271396 216496 271448
rect 216548 271436 216554 271448
rect 273254 271436 273260 271448
rect 216548 271408 273260 271436
rect 216548 271396 216554 271408
rect 273254 271396 273260 271408
rect 273312 271396 273318 271448
rect 343450 271396 343456 271448
rect 343508 271436 343514 271448
rect 358814 271436 358820 271448
rect 343508 271408 358820 271436
rect 343508 271396 343514 271408
rect 358814 271396 358820 271408
rect 358872 271396 358878 271448
rect 370866 271396 370872 271448
rect 370924 271436 370930 271448
rect 447134 271436 447140 271448
rect 370924 271408 447140 271436
rect 370924 271396 370930 271408
rect 447134 271396 447140 271408
rect 447192 271396 447198 271448
rect 53190 271328 53196 271380
rect 53248 271368 53254 271380
rect 113542 271368 113548 271380
rect 53248 271340 113548 271368
rect 53248 271328 53254 271340
rect 113542 271328 113548 271340
rect 113600 271328 113606 271380
rect 214834 271328 214840 271380
rect 214892 271368 214898 271380
rect 223574 271368 223580 271380
rect 214892 271340 223580 271368
rect 214892 271328 214898 271340
rect 223574 271328 223580 271340
rect 223632 271328 223638 271380
rect 224218 271328 224224 271380
rect 224276 271368 224282 271380
rect 268010 271368 268016 271380
rect 224276 271340 268016 271368
rect 224276 271328 224282 271340
rect 268010 271328 268016 271340
rect 268068 271328 268074 271380
rect 278682 271328 278688 271380
rect 278740 271368 278746 271380
rect 357434 271368 357440 271380
rect 278740 271340 357440 271368
rect 278740 271328 278746 271340
rect 357434 271328 357440 271340
rect 357492 271328 357498 271380
rect 372062 271328 372068 271380
rect 372120 271368 372126 271380
rect 445754 271368 445760 271380
rect 372120 271340 445760 271368
rect 372120 271328 372126 271340
rect 445754 271328 445760 271340
rect 445812 271328 445818 271380
rect 52914 271260 52920 271312
rect 52972 271300 52978 271312
rect 110414 271300 110420 271312
rect 52972 271272 110420 271300
rect 52972 271260 52978 271272
rect 110414 271260 110420 271272
rect 110472 271260 110478 271312
rect 183462 271260 183468 271312
rect 183520 271300 183526 271312
rect 197354 271300 197360 271312
rect 183520 271272 197360 271300
rect 183520 271260 183526 271272
rect 197354 271260 197360 271272
rect 197412 271260 197418 271312
rect 205082 271260 205088 271312
rect 205140 271300 205146 271312
rect 255314 271300 255320 271312
rect 205140 271272 255320 271300
rect 205140 271260 205146 271272
rect 255314 271260 255320 271272
rect 255372 271260 255378 271312
rect 277210 271260 277216 271312
rect 277268 271300 277274 271312
rect 357158 271300 357164 271312
rect 277268 271272 357164 271300
rect 277268 271260 277274 271272
rect 357158 271260 357164 271272
rect 357216 271260 357222 271312
rect 358814 271260 358820 271312
rect 358872 271300 358878 271312
rect 360010 271300 360016 271312
rect 358872 271272 360016 271300
rect 358872 271260 358878 271272
rect 360010 271260 360016 271272
rect 360068 271260 360074 271312
rect 366910 271260 366916 271312
rect 366968 271300 366974 271312
rect 434714 271300 434720 271312
rect 366968 271272 434720 271300
rect 366968 271260 366974 271272
rect 434714 271260 434720 271272
rect 434772 271260 434778 271312
rect 503622 271260 503628 271312
rect 503680 271300 503686 271312
rect 517698 271300 517704 271312
rect 503680 271272 517704 271300
rect 503680 271260 503686 271272
rect 517698 271260 517704 271272
rect 517756 271260 517762 271312
rect 51718 271192 51724 271244
rect 51776 271232 51782 271244
rect 104894 271232 104900 271244
rect 51776 271204 104900 271232
rect 51776 271192 51782 271204
rect 104894 271192 104900 271204
rect 104952 271192 104958 271244
rect 210694 271192 210700 271244
rect 210752 271232 210758 271244
rect 260834 271232 260840 271244
rect 210752 271204 260840 271232
rect 210752 271192 210758 271204
rect 260834 271192 260840 271204
rect 260892 271192 260898 271244
rect 280062 271192 280068 271244
rect 280120 271232 280126 271244
rect 358832 271232 358860 271260
rect 280120 271204 358860 271232
rect 280120 271192 280126 271204
rect 367922 271192 367928 271244
rect 367980 271232 367986 271244
rect 367980 271204 423076 271232
rect 367980 271192 367986 271204
rect 51902 271124 51908 271176
rect 51960 271164 51966 271176
rect 103514 271164 103520 271176
rect 51960 271136 103520 271164
rect 51960 271124 51966 271136
rect 103514 271124 103520 271136
rect 103572 271124 103578 271176
rect 183462 271124 183468 271176
rect 183520 271164 183526 271176
rect 201586 271164 201592 271176
rect 183520 271136 201592 271164
rect 183520 271124 183526 271136
rect 201586 271124 201592 271136
rect 201644 271124 201650 271176
rect 209498 271124 209504 271176
rect 209556 271164 209562 271176
rect 258258 271164 258264 271176
rect 209556 271136 258264 271164
rect 209556 271124 209562 271136
rect 258258 271124 258264 271136
rect 258316 271124 258322 271176
rect 275922 271124 275928 271176
rect 275980 271164 275986 271176
rect 356606 271164 356612 271176
rect 275980 271136 356612 271164
rect 275980 271124 275986 271136
rect 356606 271124 356612 271136
rect 356664 271164 356670 271176
rect 356882 271164 356888 271176
rect 356664 271136 356888 271164
rect 356664 271124 356670 271136
rect 356882 271124 356888 271136
rect 356940 271124 356946 271176
rect 373534 271124 373540 271176
rect 373592 271164 373598 271176
rect 373592 271136 422892 271164
rect 373592 271124 373598 271136
rect 50246 271056 50252 271108
rect 50304 271096 50310 271108
rect 100754 271096 100760 271108
rect 50304 271068 100760 271096
rect 50304 271056 50310 271068
rect 100754 271056 100760 271068
rect 100812 271056 100818 271108
rect 219526 271056 219532 271108
rect 219584 271096 219590 271108
rect 268102 271096 268108 271108
rect 219584 271068 268108 271096
rect 219584 271056 219590 271068
rect 268102 271056 268108 271068
rect 268160 271056 268166 271108
rect 375098 271056 375104 271108
rect 375156 271096 375162 271108
rect 420914 271096 420920 271108
rect 375156 271068 420920 271096
rect 375156 271056 375162 271068
rect 420914 271056 420920 271068
rect 420972 271056 420978 271108
rect 46658 270988 46664 271040
rect 46716 271028 46722 271040
rect 77294 271028 77300 271040
rect 46716 271000 77300 271028
rect 46716 270988 46722 271000
rect 77294 270988 77300 271000
rect 77352 270988 77358 271040
rect 210786 270988 210792 271040
rect 210844 271028 210850 271040
rect 252554 271028 252560 271040
rect 210844 271000 252560 271028
rect 210844 270988 210850 271000
rect 252554 270988 252560 271000
rect 252612 270988 252618 271040
rect 373626 270988 373632 271040
rect 373684 271028 373690 271040
rect 418338 271028 418344 271040
rect 373684 271000 418344 271028
rect 373684 270988 373690 271000
rect 418338 270988 418344 271000
rect 418396 270988 418402 271040
rect 422864 271028 422892 271136
rect 423048 271096 423076 271204
rect 437474 271164 437480 271176
rect 437446 271124 437480 271164
rect 437532 271124 437538 271176
rect 503530 271124 503536 271176
rect 503588 271164 503594 271176
rect 517606 271164 517612 271176
rect 503588 271136 517612 271164
rect 503588 271124 503594 271136
rect 517606 271124 517612 271136
rect 517664 271124 517670 271176
rect 433334 271096 433340 271108
rect 423048 271068 433340 271096
rect 433334 271056 433340 271068
rect 433392 271056 433398 271108
rect 437446 271028 437474 271124
rect 422864 271000 437474 271028
rect 47946 270920 47952 270972
rect 48004 270960 48010 270972
rect 78674 270960 78680 270972
rect 48004 270932 78680 270960
rect 48004 270920 48010 270932
rect 78674 270920 78680 270932
rect 78732 270920 78738 270972
rect 219158 270920 219164 270972
rect 219216 270960 219222 270972
rect 247034 270960 247040 270972
rect 219216 270932 247040 270960
rect 219216 270920 219222 270932
rect 247034 270920 247040 270932
rect 247092 270920 247098 270972
rect 375006 270920 375012 270972
rect 375064 270960 375070 270972
rect 409874 270960 409880 270972
rect 375064 270932 409880 270960
rect 375064 270920 375070 270932
rect 409874 270920 409880 270932
rect 409932 270920 409938 270972
rect 215202 270852 215208 270904
rect 215260 270892 215266 270904
rect 224218 270892 224224 270904
rect 215260 270864 224224 270892
rect 215260 270852 215266 270864
rect 224218 270852 224224 270864
rect 224276 270852 224282 270904
rect 264238 270852 264244 270904
rect 264296 270892 264302 270904
rect 266354 270892 266360 270904
rect 264296 270864 266360 270892
rect 264296 270852 264302 270864
rect 266354 270852 266360 270864
rect 266412 270852 266418 270904
rect 425698 270852 425704 270904
rect 425756 270892 425762 270904
rect 429194 270892 429200 270904
rect 425756 270864 429200 270892
rect 425756 270852 425762 270864
rect 429194 270852 429200 270864
rect 429252 270852 429258 270904
rect 517606 270784 517612 270836
rect 517664 270824 517670 270836
rect 517882 270824 517888 270836
rect 517664 270796 517888 270824
rect 517664 270784 517670 270796
rect 517882 270784 517888 270796
rect 517940 270784 517946 270836
rect 422938 270580 422944 270632
rect 422996 270620 423002 270632
rect 437474 270620 437480 270632
rect 422996 270592 437480 270620
rect 422996 270580 423002 270592
rect 437474 270580 437480 270592
rect 437532 270580 437538 270632
rect 102778 270512 102784 270564
rect 102836 270552 102842 270564
rect 113174 270552 113180 270564
rect 102836 270524 113180 270552
rect 102836 270512 102842 270524
rect 113174 270512 113180 270524
rect 113232 270512 113238 270564
rect 268838 270512 268844 270564
rect 268896 270552 268902 270564
rect 273254 270552 273260 270564
rect 268896 270524 273260 270552
rect 268896 270512 268902 270524
rect 273254 270512 273260 270524
rect 273312 270512 273318 270564
rect 421558 270512 421564 270564
rect 421616 270552 421622 270564
rect 436094 270552 436100 270564
rect 421616 270524 436100 270552
rect 421616 270512 421622 270524
rect 436094 270512 436100 270524
rect 436152 270512 436158 270564
rect 44910 270444 44916 270496
rect 44968 270484 44974 270496
rect 147674 270484 147680 270496
rect 44968 270456 147680 270484
rect 44968 270444 44974 270456
rect 147674 270444 147680 270456
rect 147732 270444 147738 270496
rect 210326 270444 210332 270496
rect 210384 270484 210390 270496
rect 210878 270484 210884 270496
rect 210384 270456 210884 270484
rect 210384 270444 210390 270456
rect 210878 270444 210884 270456
rect 210936 270444 210942 270496
rect 211522 270444 211528 270496
rect 211580 270484 211586 270496
rect 216950 270484 216956 270496
rect 211580 270456 216956 270484
rect 211580 270444 211586 270456
rect 216950 270444 216956 270456
rect 217008 270444 217014 270496
rect 224218 270444 224224 270496
rect 224276 270484 224282 270496
rect 262214 270484 262220 270496
rect 224276 270456 262220 270484
rect 224276 270444 224282 270456
rect 262214 270444 262220 270456
rect 262272 270444 262278 270496
rect 369762 270444 369768 270496
rect 369820 270484 369826 270496
rect 371694 270484 371700 270496
rect 369820 270456 371700 270484
rect 369820 270444 369826 270456
rect 371694 270444 371700 270456
rect 371752 270444 371758 270496
rect 379330 270444 379336 270496
rect 379388 270484 379394 270496
rect 379514 270484 379520 270496
rect 379388 270456 379520 270484
rect 379388 270444 379394 270456
rect 379514 270444 379520 270456
rect 379572 270444 379578 270496
rect 379974 270444 379980 270496
rect 380032 270484 380038 270496
rect 396074 270484 396080 270496
rect 380032 270456 396080 270484
rect 380032 270444 380038 270456
rect 396074 270444 396080 270456
rect 396132 270444 396138 270496
rect 58710 270376 58716 270428
rect 58768 270416 58774 270428
rect 115934 270416 115940 270428
rect 58768 270388 115940 270416
rect 58768 270376 58774 270388
rect 115934 270376 115940 270388
rect 115992 270376 115998 270428
rect 212350 270376 212356 270428
rect 212408 270416 212414 270428
rect 244274 270416 244280 270428
rect 212408 270388 244280 270416
rect 212408 270376 212414 270388
rect 244274 270376 244280 270388
rect 244332 270376 244338 270428
rect 378594 270376 378600 270428
rect 378652 270416 378658 270428
rect 379606 270416 379612 270428
rect 378652 270388 379612 270416
rect 378652 270376 378658 270388
rect 379606 270376 379612 270388
rect 379664 270376 379670 270428
rect 380066 270376 380072 270428
rect 380124 270416 380130 270428
rect 411254 270416 411260 270428
rect 380124 270388 411260 270416
rect 380124 270376 380130 270388
rect 411254 270376 411260 270388
rect 411312 270376 411318 270428
rect 60734 270308 60740 270360
rect 60792 270348 60798 270360
rect 91094 270348 91100 270360
rect 60792 270320 91100 270348
rect 60792 270308 60798 270320
rect 91094 270308 91100 270320
rect 91152 270308 91158 270360
rect 210970 270308 210976 270360
rect 211028 270348 211034 270360
rect 214834 270348 214840 270360
rect 211028 270320 214840 270348
rect 211028 270308 211034 270320
rect 214834 270308 214840 270320
rect 214892 270308 214898 270360
rect 219618 270308 219624 270360
rect 219676 270348 219682 270360
rect 220446 270348 220452 270360
rect 219676 270320 220452 270348
rect 219676 270308 219682 270320
rect 220446 270308 220452 270320
rect 220504 270348 220510 270360
rect 249794 270348 249800 270360
rect 220504 270320 249800 270348
rect 220504 270308 220510 270320
rect 249794 270308 249800 270320
rect 249852 270308 249858 270360
rect 368290 270308 368296 270360
rect 368348 270348 368354 270360
rect 398834 270348 398840 270360
rect 368348 270320 398840 270348
rect 368348 270308 368354 270320
rect 398834 270308 398840 270320
rect 398892 270308 398898 270360
rect 79042 270240 79048 270292
rect 79100 270280 79106 270292
rect 110414 270280 110420 270292
rect 79100 270252 110420 270280
rect 79100 270240 79106 270252
rect 110414 270240 110420 270252
rect 110472 270240 110478 270292
rect 220170 270240 220176 270292
rect 220228 270280 220234 270292
rect 248506 270280 248512 270292
rect 220228 270252 248512 270280
rect 220228 270240 220234 270252
rect 248506 270240 248512 270252
rect 248564 270240 248570 270292
rect 377030 270240 377036 270292
rect 377088 270280 377094 270292
rect 380066 270280 380072 270292
rect 377088 270252 380072 270280
rect 377088 270240 377094 270252
rect 380066 270240 380072 270252
rect 380124 270240 380130 270292
rect 405734 270280 405740 270292
rect 380176 270252 405740 270280
rect 58618 270172 58624 270224
rect 58676 270212 58682 270224
rect 89714 270212 89720 270224
rect 58676 270184 89720 270212
rect 58676 270172 58682 270184
rect 89714 270172 89720 270184
rect 89772 270172 89778 270224
rect 217226 270172 217232 270224
rect 217284 270212 217290 270224
rect 219894 270212 219900 270224
rect 217284 270184 219900 270212
rect 217284 270172 217290 270184
rect 219894 270172 219900 270184
rect 219952 270212 219958 270224
rect 251266 270212 251272 270224
rect 219952 270184 251272 270212
rect 219952 270172 219958 270184
rect 251266 270172 251272 270184
rect 251324 270172 251330 270224
rect 376478 270172 376484 270224
rect 376536 270212 376542 270224
rect 380176 270212 380204 270252
rect 405734 270240 405740 270252
rect 405792 270240 405798 270292
rect 376536 270184 380204 270212
rect 376536 270172 376542 270184
rect 380250 270172 380256 270224
rect 380308 270212 380314 270224
rect 404354 270212 404360 270224
rect 380308 270184 404360 270212
rect 380308 270172 380314 270184
rect 404354 270172 404360 270184
rect 404412 270172 404418 270224
rect 56502 270104 56508 270156
rect 56560 270144 56566 270156
rect 86954 270144 86960 270156
rect 56560 270116 86960 270144
rect 56560 270104 56566 270116
rect 86954 270104 86960 270116
rect 87012 270104 87018 270156
rect 210878 270104 210884 270156
rect 210936 270144 210942 270156
rect 239122 270144 239128 270156
rect 210936 270116 239128 270144
rect 210936 270104 210942 270116
rect 239122 270104 239128 270116
rect 239180 270104 239186 270156
rect 371694 270104 371700 270156
rect 371752 270144 371758 270156
rect 397454 270144 397460 270156
rect 371752 270116 397460 270144
rect 371752 270104 371758 270116
rect 397454 270104 397460 270116
rect 397512 270104 397518 270156
rect 59354 270036 59360 270088
rect 59412 270076 59418 270088
rect 92474 270076 92480 270088
rect 59412 270048 92480 270076
rect 59412 270036 59418 270048
rect 92474 270036 92480 270048
rect 92532 270036 92538 270088
rect 215202 270036 215208 270088
rect 215260 270076 215266 270088
rect 219434 270076 219440 270088
rect 215260 270048 219440 270076
rect 215260 270036 215266 270048
rect 219434 270036 219440 270048
rect 219492 270076 219498 270088
rect 220538 270076 220544 270088
rect 219492 270048 220544 270076
rect 219492 270036 219498 270048
rect 220538 270036 220544 270048
rect 220596 270036 220602 270088
rect 220630 270036 220636 270088
rect 220688 270076 220694 270088
rect 251174 270076 251180 270088
rect 220688 270048 251180 270076
rect 220688 270036 220694 270048
rect 251174 270036 251180 270048
rect 251232 270036 251238 270088
rect 371142 270036 371148 270088
rect 371200 270076 371206 270088
rect 375742 270076 375748 270088
rect 371200 270048 375748 270076
rect 371200 270036 371206 270048
rect 375742 270036 375748 270048
rect 375800 270076 375806 270088
rect 403526 270076 403532 270088
rect 375800 270048 403532 270076
rect 375800 270036 375806 270048
rect 403526 270036 403532 270048
rect 403584 270036 403590 270088
rect 51718 269968 51724 270020
rect 51776 270008 51782 270020
rect 84194 270008 84200 270020
rect 51776 269980 84200 270008
rect 51776 269968 51782 269980
rect 84194 269968 84200 269980
rect 84252 269968 84258 270020
rect 217134 269968 217140 270020
rect 217192 270008 217198 270020
rect 217318 270008 217324 270020
rect 217192 269980 217324 270008
rect 217192 269968 217198 269980
rect 217318 269968 217324 269980
rect 217376 270008 217382 270020
rect 217376 269980 219434 270008
rect 217376 269968 217382 269980
rect 53098 269900 53104 269952
rect 53156 269940 53162 269952
rect 85574 269940 85580 269952
rect 53156 269912 85580 269940
rect 53156 269900 53162 269912
rect 85574 269900 85580 269912
rect 85632 269900 85638 269952
rect 88242 269900 88248 269952
rect 88300 269940 88306 269952
rect 106274 269940 106280 269952
rect 88300 269912 106280 269940
rect 88300 269900 88306 269912
rect 106274 269900 106280 269912
rect 106332 269900 106338 269952
rect 214282 269900 214288 269952
rect 214340 269940 214346 269952
rect 214926 269940 214932 269952
rect 214340 269912 214932 269940
rect 214340 269900 214346 269912
rect 214926 269900 214932 269912
rect 214984 269900 214990 269952
rect 219406 269940 219434 269980
rect 220722 269968 220728 270020
rect 220780 270008 220786 270020
rect 252554 270008 252560 270020
rect 220780 269980 252560 270008
rect 220780 269968 220786 269980
rect 252554 269968 252560 269980
rect 252612 269968 252618 270020
rect 371050 269968 371056 270020
rect 371108 270008 371114 270020
rect 372062 270008 372068 270020
rect 371108 269980 372068 270008
rect 371108 269968 371114 269980
rect 372062 269968 372068 269980
rect 372120 270008 372126 270020
rect 400214 270008 400220 270020
rect 372120 269980 400220 270008
rect 372120 269968 372126 269980
rect 400214 269968 400220 269980
rect 400272 269968 400278 270020
rect 263594 269940 263600 269952
rect 219406 269912 263600 269940
rect 263594 269900 263600 269912
rect 263652 269900 263658 269952
rect 376662 269900 376668 269952
rect 376720 269940 376726 269952
rect 389174 269940 389180 269952
rect 376720 269912 389180 269940
rect 376720 269900 376726 269912
rect 389174 269900 389180 269912
rect 389232 269940 389238 269952
rect 419534 269940 419540 269952
rect 389232 269912 419540 269940
rect 389232 269900 389238 269912
rect 419534 269900 419540 269912
rect 419592 269900 419598 269952
rect 57974 269832 57980 269884
rect 58032 269872 58038 269884
rect 103698 269872 103704 269884
rect 58032 269844 103704 269872
rect 58032 269832 58038 269844
rect 103698 269832 103704 269844
rect 103756 269832 103762 269884
rect 115842 269832 115848 269884
rect 115900 269872 115906 269884
rect 196710 269872 196716 269884
rect 115900 269844 196716 269872
rect 115900 269832 115906 269844
rect 196710 269832 196716 269844
rect 196768 269872 196774 269884
rect 204346 269872 204352 269884
rect 196768 269844 204352 269872
rect 196768 269832 196774 269844
rect 204346 269832 204352 269844
rect 204404 269832 204410 269884
rect 214834 269832 214840 269884
rect 214892 269872 214898 269884
rect 269114 269872 269120 269884
rect 214892 269844 269120 269872
rect 214892 269832 214898 269844
rect 269114 269832 269120 269844
rect 269172 269832 269178 269884
rect 373810 269832 373816 269884
rect 373868 269872 373874 269884
rect 375834 269872 375840 269884
rect 373868 269844 375840 269872
rect 373868 269832 373874 269844
rect 375834 269832 375840 269844
rect 375892 269872 375898 269884
rect 407114 269872 407120 269884
rect 375892 269844 407120 269872
rect 375892 269832 375898 269844
rect 407114 269832 407120 269844
rect 407172 269832 407178 269884
rect 56870 269764 56876 269816
rect 56928 269804 56934 269816
rect 104894 269804 104900 269816
rect 56928 269776 104900 269804
rect 56928 269764 56934 269776
rect 104894 269764 104900 269776
rect 104952 269764 104958 269816
rect 114462 269764 114468 269816
rect 114520 269804 114526 269816
rect 196618 269804 196624 269816
rect 114520 269776 196624 269804
rect 114520 269764 114526 269776
rect 196618 269764 196624 269776
rect 196676 269804 196682 269816
rect 202874 269804 202880 269816
rect 196676 269776 202880 269804
rect 196676 269764 196682 269776
rect 202874 269764 202880 269776
rect 202932 269764 202938 269816
rect 206830 269764 206836 269816
rect 206888 269804 206894 269816
rect 212994 269804 213000 269816
rect 206888 269776 213000 269804
rect 206888 269764 206894 269776
rect 212994 269764 213000 269776
rect 213052 269804 213058 269816
rect 270494 269804 270500 269816
rect 213052 269776 270500 269804
rect 213052 269764 213058 269776
rect 270494 269764 270500 269776
rect 270552 269764 270558 269816
rect 379514 269764 379520 269816
rect 379572 269804 379578 269816
rect 413002 269804 413008 269816
rect 379572 269776 413008 269804
rect 379572 269764 379578 269776
rect 413002 269764 413008 269776
rect 413060 269764 413066 269816
rect 62114 269696 62120 269748
rect 62172 269736 62178 269748
rect 91186 269736 91192 269748
rect 62172 269708 91192 269736
rect 62172 269696 62178 269708
rect 91186 269696 91192 269708
rect 91244 269696 91250 269748
rect 216950 269696 216956 269748
rect 217008 269736 217014 269748
rect 245654 269736 245660 269748
rect 217008 269708 245660 269736
rect 217008 269696 217014 269708
rect 245654 269696 245660 269708
rect 245712 269696 245718 269748
rect 372338 269696 372344 269748
rect 372396 269736 372402 269748
rect 375282 269736 375288 269748
rect 372396 269708 375288 269736
rect 372396 269696 372402 269708
rect 375282 269696 375288 269708
rect 375340 269736 375346 269748
rect 401686 269736 401692 269748
rect 375340 269708 401692 269736
rect 375340 269696 375346 269708
rect 401686 269696 401692 269708
rect 401744 269696 401750 269748
rect 81434 269628 81440 269680
rect 81492 269668 81498 269680
rect 107654 269668 107660 269680
rect 81492 269640 107660 269668
rect 81492 269628 81498 269640
rect 107654 269628 107660 269640
rect 107712 269628 107718 269680
rect 206922 269628 206928 269680
rect 206980 269668 206986 269680
rect 210786 269668 210792 269680
rect 206980 269640 210792 269668
rect 206980 269628 206986 269640
rect 210786 269628 210792 269640
rect 210844 269668 210850 269680
rect 237374 269668 237380 269680
rect 210844 269640 237380 269668
rect 210844 269628 210850 269640
rect 237374 269628 237380 269640
rect 237432 269628 237438 269680
rect 391934 269668 391940 269680
rect 376588 269640 391940 269668
rect 376588 269612 376616 269640
rect 391934 269628 391940 269640
rect 391992 269628 391998 269680
rect 83458 269560 83464 269612
rect 83516 269600 83522 269612
rect 106366 269600 106372 269612
rect 83516 269572 106372 269600
rect 83516 269560 83522 269572
rect 106366 269560 106372 269572
rect 106424 269560 106430 269612
rect 220538 269560 220544 269612
rect 220596 269600 220602 269612
rect 247034 269600 247040 269612
rect 220596 269572 247040 269600
rect 220596 269560 220602 269572
rect 247034 269560 247040 269572
rect 247092 269560 247098 269612
rect 375098 269560 375104 269612
rect 375156 269600 375162 269612
rect 376570 269600 376576 269612
rect 375156 269572 376576 269600
rect 375156 269560 375162 269572
rect 376570 269560 376576 269572
rect 376628 269560 376634 269612
rect 379606 269560 379612 269612
rect 379664 269600 379670 269612
rect 411346 269600 411352 269612
rect 379664 269572 411352 269600
rect 379664 269560 379670 269572
rect 411346 269560 411352 269572
rect 411404 269560 411410 269612
rect 214926 269492 214932 269544
rect 214984 269532 214990 269544
rect 224218 269532 224224 269544
rect 214984 269504 224224 269532
rect 214984 269492 214990 269504
rect 224218 269492 224224 269504
rect 224276 269492 224282 269544
rect 374546 269492 374552 269544
rect 374604 269532 374610 269544
rect 379974 269532 379980 269544
rect 374604 269504 379980 269532
rect 374604 269492 374610 269504
rect 379974 269492 379980 269504
rect 380032 269492 380038 269544
rect 218514 269288 218520 269340
rect 218572 269328 218578 269340
rect 219434 269328 219440 269340
rect 218572 269300 219440 269328
rect 218572 269288 218578 269300
rect 219434 269288 219440 269300
rect 219492 269328 219498 269340
rect 220722 269328 220728 269340
rect 219492 269300 220728 269328
rect 219492 269288 219498 269300
rect 220722 269288 220728 269300
rect 220780 269288 220786 269340
rect 218606 269220 218612 269272
rect 218664 269260 218670 269272
rect 219802 269260 219808 269272
rect 218664 269232 219808 269260
rect 218664 269220 218670 269232
rect 219802 269220 219808 269232
rect 219860 269260 219866 269272
rect 220630 269260 220636 269272
rect 219860 269232 220636 269260
rect 219860 269220 219866 269232
rect 220630 269220 220636 269232
rect 220688 269220 220694 269272
rect 216490 269152 216496 269204
rect 216548 269192 216554 269204
rect 220170 269192 220176 269204
rect 216548 269164 220176 269192
rect 216548 269152 216554 269164
rect 220170 269152 220176 269164
rect 220228 269152 220234 269204
rect 373626 269152 373632 269204
rect 373684 269192 373690 269204
rect 376478 269192 376484 269204
rect 373684 269164 376484 269192
rect 373684 269152 373690 269164
rect 376478 269152 376484 269164
rect 376536 269152 376542 269204
rect 219158 269084 219164 269136
rect 219216 269124 219222 269136
rect 220446 269124 220452 269136
rect 219216 269096 220452 269124
rect 219216 269084 219222 269096
rect 220446 269084 220452 269096
rect 220504 269084 220510 269136
rect 373718 269084 373724 269136
rect 373776 269124 373782 269136
rect 375190 269124 375196 269136
rect 373776 269096 375196 269124
rect 373776 269084 373782 269096
rect 375190 269084 375196 269096
rect 375248 269124 375254 269136
rect 380250 269124 380256 269136
rect 375248 269096 380256 269124
rect 375248 269084 375254 269096
rect 380250 269084 380256 269096
rect 380308 269084 380314 269136
rect 48130 269016 48136 269068
rect 48188 269056 48194 269068
rect 53098 269056 53104 269068
rect 48188 269028 53104 269056
rect 48188 269016 48194 269028
rect 53098 269016 53104 269028
rect 53156 269016 53162 269068
rect 205634 269016 205640 269068
rect 205692 269056 205698 269068
rect 256694 269056 256700 269068
rect 205692 269028 256700 269056
rect 205692 269016 205698 269028
rect 256694 269016 256700 269028
rect 256752 269016 256758 269068
rect 370958 269016 370964 269068
rect 371016 269056 371022 269068
rect 373534 269056 373540 269068
rect 371016 269028 373540 269056
rect 371016 269016 371022 269028
rect 373534 269016 373540 269028
rect 373592 269016 373598 269068
rect 376754 269016 376760 269068
rect 376812 269056 376818 269068
rect 377122 269056 377128 269068
rect 376812 269028 377128 269056
rect 376812 269016 376818 269028
rect 377122 269016 377128 269028
rect 377180 269016 377186 269068
rect 377214 269016 377220 269068
rect 377272 269056 377278 269068
rect 379054 269056 379060 269068
rect 377272 269028 379060 269056
rect 377272 269016 377278 269028
rect 379054 269016 379060 269028
rect 379112 269016 379118 269068
rect 379238 269016 379244 269068
rect 379296 269056 379302 269068
rect 420914 269056 420920 269068
rect 379296 269028 420920 269056
rect 379296 269016 379302 269028
rect 420914 269016 420920 269028
rect 420972 269016 420978 269068
rect 46842 268948 46848 269000
rect 46900 268988 46906 269000
rect 51718 268988 51724 269000
rect 46900 268960 51724 268988
rect 46900 268948 46906 268960
rect 51718 268948 51724 268960
rect 51776 268948 51782 269000
rect 217226 268948 217232 269000
rect 217284 268988 217290 269000
rect 217962 268988 217968 269000
rect 217284 268960 217968 268988
rect 217284 268948 217290 268960
rect 217962 268948 217968 268960
rect 218020 268988 218026 269000
rect 255314 268988 255320 269000
rect 218020 268960 255320 268988
rect 218020 268948 218026 268960
rect 255314 268948 255320 268960
rect 255372 268948 255378 269000
rect 44082 268880 44088 268932
rect 44140 268920 44146 268932
rect 59354 268920 59360 268932
rect 44140 268892 59360 268920
rect 44140 268880 44146 268892
rect 59354 268880 59360 268892
rect 59412 268880 59418 268932
rect 219710 268880 219716 268932
rect 219768 268920 219774 268932
rect 253934 268920 253940 268932
rect 219768 268892 253940 268920
rect 219768 268880 219774 268892
rect 253934 268880 253940 268892
rect 253992 268880 253998 268932
rect 377140 268920 377168 269016
rect 378686 268948 378692 269000
rect 378744 268988 378750 269000
rect 418522 268988 418528 269000
rect 378744 268960 418528 268988
rect 378744 268948 378750 268960
rect 418522 268948 418528 268960
rect 418580 268948 418586 269000
rect 415394 268920 415400 268932
rect 377140 268892 415400 268920
rect 415394 268880 415400 268892
rect 415452 268880 415458 268932
rect 43622 268812 43628 268864
rect 43680 268852 43686 268864
rect 56870 268852 56876 268864
rect 43680 268824 56876 268852
rect 43680 268812 43686 268824
rect 56870 268812 56876 268824
rect 56928 268812 56934 268864
rect 213730 268812 213736 268864
rect 213788 268852 213794 268864
rect 244366 268852 244372 268864
rect 213788 268824 244372 268852
rect 213788 268812 213794 268824
rect 244366 268812 244372 268824
rect 244424 268812 244430 268864
rect 376570 268812 376576 268864
rect 376628 268852 376634 268864
rect 378686 268852 378692 268864
rect 376628 268824 378692 268852
rect 376628 268812 376634 268824
rect 378686 268812 378692 268824
rect 378744 268812 378750 268864
rect 379238 268852 379244 268864
rect 379072 268824 379244 268852
rect 48222 268744 48228 268796
rect 48280 268784 48286 268796
rect 58618 268784 58624 268796
rect 48280 268756 58624 268784
rect 48280 268744 48286 268756
rect 58618 268744 58624 268756
rect 58676 268744 58682 268796
rect 216398 268744 216404 268796
rect 216456 268784 216462 268796
rect 242894 268784 242900 268796
rect 216456 268756 242900 268784
rect 216456 268744 216462 268756
rect 242894 268744 242900 268756
rect 242952 268744 242958 268796
rect 374454 268744 374460 268796
rect 374512 268784 374518 268796
rect 379072 268784 379100 268824
rect 379238 268812 379244 268824
rect 379296 268812 379302 268864
rect 379882 268812 379888 268864
rect 379940 268852 379946 268864
rect 414014 268852 414020 268864
rect 379940 268824 414020 268852
rect 379940 268812 379946 268824
rect 414014 268812 414020 268824
rect 414072 268812 414078 268864
rect 374512 268756 379100 268784
rect 374512 268744 374518 268756
rect 379146 268744 379152 268796
rect 379204 268784 379210 268796
rect 408494 268784 408500 268796
rect 379204 268756 408500 268784
rect 379204 268744 379210 268756
rect 408494 268744 408500 268756
rect 408552 268744 408558 268796
rect 46750 268676 46756 268728
rect 46808 268716 46814 268728
rect 55766 268716 55772 268728
rect 46808 268688 55772 268716
rect 46808 268676 46814 268688
rect 55766 268676 55772 268688
rect 55824 268716 55830 268728
rect 56502 268716 56508 268728
rect 55824 268688 56508 268716
rect 55824 268676 55830 268688
rect 56502 268676 56508 268688
rect 56560 268676 56566 268728
rect 214466 268676 214472 268728
rect 214524 268716 214530 268728
rect 235994 268716 236000 268728
rect 214524 268688 236000 268716
rect 214524 268676 214530 268688
rect 235994 268676 236000 268688
rect 236052 268676 236058 268728
rect 391934 268676 391940 268728
rect 391992 268716 391998 268728
rect 418154 268716 418160 268728
rect 391992 268688 418160 268716
rect 391992 268676 391998 268688
rect 418154 268676 418160 268688
rect 418212 268676 418218 268728
rect 43990 268608 43996 268660
rect 44048 268648 44054 268660
rect 48130 268648 48136 268660
rect 44048 268620 48136 268648
rect 44048 268608 44054 268620
rect 48130 268608 48136 268620
rect 48188 268648 48194 268660
rect 60734 268648 60740 268660
rect 48188 268620 60740 268648
rect 48188 268608 48194 268620
rect 60734 268608 60740 268620
rect 60792 268608 60798 268660
rect 213086 268608 213092 268660
rect 213144 268648 213150 268660
rect 233234 268648 233240 268660
rect 213144 268620 233240 268648
rect 213144 268608 213150 268620
rect 233234 268608 233240 268620
rect 233292 268648 233298 268660
rect 258074 268648 258080 268660
rect 233292 268620 258080 268648
rect 233292 268608 233298 268620
rect 258074 268608 258080 268620
rect 258132 268608 258138 268660
rect 46566 268540 46572 268592
rect 46624 268580 46630 268592
rect 48222 268580 48228 268592
rect 46624 268552 48228 268580
rect 46624 268540 46630 268552
rect 48222 268540 48228 268552
rect 48280 268580 48286 268592
rect 62114 268580 62120 268592
rect 48280 268552 62120 268580
rect 48280 268540 48286 268552
rect 62114 268540 62120 268552
rect 62172 268540 62178 268592
rect 214374 268540 214380 268592
rect 214432 268580 214438 268592
rect 231854 268580 231860 268592
rect 214432 268552 231860 268580
rect 214432 268540 214438 268552
rect 231854 268540 231860 268552
rect 231912 268580 231918 268592
rect 259454 268580 259460 268592
rect 231912 268552 259460 268580
rect 231912 268540 231918 268552
rect 259454 268540 259460 268552
rect 259512 268540 259518 268592
rect 43714 268472 43720 268524
rect 43772 268512 43778 268524
rect 47578 268512 47584 268524
rect 43772 268484 47584 268512
rect 43772 268472 43778 268484
rect 47578 268472 47584 268484
rect 47636 268512 47642 268524
rect 79042 268512 79048 268524
rect 47636 268484 79048 268512
rect 47636 268472 47642 268484
rect 79042 268472 79048 268484
rect 79100 268472 79106 268524
rect 215846 268472 215852 268524
rect 215904 268512 215910 268524
rect 230474 268512 230480 268524
rect 215904 268484 230480 268512
rect 215904 268472 215910 268484
rect 230474 268472 230480 268484
rect 230532 268512 230538 268524
rect 259546 268512 259552 268524
rect 230532 268484 259552 268512
rect 230532 268472 230538 268484
rect 259546 268472 259552 268484
rect 259604 268472 259610 268524
rect 372246 268472 372252 268524
rect 372304 268512 372310 268524
rect 379238 268512 379244 268524
rect 372304 268484 379244 268512
rect 372304 268472 372310 268484
rect 379238 268472 379244 268484
rect 379296 268512 379302 268524
rect 402974 268512 402980 268524
rect 379296 268484 402980 268512
rect 379296 268472 379302 268484
rect 402974 268472 402980 268484
rect 403032 268472 403038 268524
rect 43898 268404 43904 268456
rect 43956 268444 43962 268456
rect 47762 268444 47768 268456
rect 43956 268416 47768 268444
rect 43956 268404 43962 268416
rect 47762 268404 47768 268416
rect 47820 268444 47826 268456
rect 81434 268444 81440 268456
rect 47820 268416 81440 268444
rect 47820 268404 47826 268416
rect 81434 268404 81440 268416
rect 81492 268404 81498 268456
rect 208302 268404 208308 268456
rect 208360 268444 208366 268456
rect 214466 268444 214472 268456
rect 208360 268416 214472 268444
rect 208360 268404 208366 268416
rect 214466 268404 214472 268416
rect 214524 268404 214530 268456
rect 230382 268404 230388 268456
rect 230440 268444 230446 268456
rect 260834 268444 260840 268456
rect 230440 268416 260840 268444
rect 230440 268404 230446 268416
rect 260834 268404 260840 268416
rect 260892 268404 260898 268456
rect 379054 268404 379060 268456
rect 379112 268444 379118 268456
rect 409874 268444 409880 268456
rect 379112 268416 409880 268444
rect 379112 268404 379118 268416
rect 409874 268404 409880 268416
rect 409932 268404 409938 268456
rect 43806 268336 43812 268388
rect 43864 268376 43870 268388
rect 47670 268376 47676 268388
rect 43864 268348 47676 268376
rect 43864 268336 43870 268348
rect 47670 268336 47676 268348
rect 47728 268376 47734 268388
rect 88242 268376 88248 268388
rect 47728 268348 88248 268376
rect 47728 268336 47734 268348
rect 88242 268336 88248 268348
rect 88300 268336 88306 268388
rect 207566 268336 207572 268388
rect 207624 268376 207630 268388
rect 212166 268376 212172 268388
rect 207624 268348 212172 268376
rect 207624 268336 207630 268348
rect 212166 268336 212172 268348
rect 212224 268376 212230 268388
rect 268838 268376 268844 268388
rect 212224 268348 268844 268376
rect 212224 268336 212230 268348
rect 268838 268336 268844 268348
rect 268896 268336 268902 268388
rect 373534 268336 373540 268388
rect 373592 268376 373598 268388
rect 431954 268376 431960 268388
rect 373592 268348 431960 268376
rect 373592 268336 373598 268348
rect 431954 268336 431960 268348
rect 432012 268336 432018 268388
rect 43530 268268 43536 268320
rect 43588 268308 43594 268320
rect 128354 268308 128360 268320
rect 43588 268280 128360 268308
rect 43588 268268 43594 268280
rect 128354 268268 128360 268280
rect 128412 268268 128418 268320
rect 40954 268200 40960 268252
rect 41012 268240 41018 268252
rect 57974 268240 57980 268252
rect 41012 268212 57980 268240
rect 41012 268200 41018 268212
rect 57974 268200 57980 268212
rect 58032 268200 58038 268252
rect 60734 268200 60740 268252
rect 60792 268240 60798 268252
rect 60918 268240 60924 268252
rect 60792 268212 60924 268240
rect 60792 268200 60798 268212
rect 60918 268200 60924 268212
rect 60976 268200 60982 268252
rect 377950 268200 377956 268252
rect 378008 268240 378014 268252
rect 379146 268240 379152 268252
rect 378008 268212 379152 268240
rect 378008 268200 378014 268212
rect 379146 268200 379152 268212
rect 379204 268200 379210 268252
rect 357526 253988 357532 254040
rect 357584 254028 357590 254040
rect 360286 254028 360292 254040
rect 357584 254000 360292 254028
rect 357584 253988 357590 254000
rect 360286 253988 360292 254000
rect 360344 253988 360350 254040
rect 357342 253960 357348 253972
rect 356532 253932 357348 253960
rect 198642 253852 198648 253904
rect 198700 253892 198706 253904
rect 200758 253892 200764 253904
rect 198700 253864 200764 253892
rect 198700 253852 198706 253864
rect 200758 253852 200764 253864
rect 200816 253852 200822 253904
rect 340782 253852 340788 253904
rect 340840 253892 340846 253904
rect 356532 253892 356560 253932
rect 357342 253920 357348 253932
rect 357400 253960 357406 253972
rect 357618 253960 357624 253972
rect 357400 253932 357624 253960
rect 357400 253920 357406 253932
rect 357618 253920 357624 253932
rect 357676 253920 357682 253972
rect 340840 253864 356560 253892
rect 340840 253852 340846 253864
rect 180150 253308 180156 253360
rect 180208 253348 180214 253360
rect 197446 253348 197452 253360
rect 180208 253320 197452 253348
rect 180208 253308 180214 253320
rect 197446 253308 197452 253320
rect 197504 253308 197510 253360
rect 500862 253308 500868 253360
rect 500920 253348 500926 253360
rect 517698 253348 517704 253360
rect 500920 253320 517704 253348
rect 500920 253308 500926 253320
rect 517698 253308 517704 253320
rect 517756 253308 517762 253360
rect 339402 253240 339408 253292
rect 339460 253280 339466 253292
rect 357526 253280 357532 253292
rect 339460 253252 357532 253280
rect 339460 253240 339466 253252
rect 357526 253240 357532 253252
rect 357584 253280 357590 253292
rect 357710 253280 357716 253292
rect 357584 253252 357716 253280
rect 357584 253240 357590 253252
rect 357710 253240 357716 253252
rect 357768 253240 357774 253292
rect 499206 253240 499212 253292
rect 499264 253280 499270 253292
rect 517606 253280 517612 253292
rect 499264 253252 517612 253280
rect 499264 253240 499270 253252
rect 517606 253240 517612 253252
rect 517664 253280 517670 253292
rect 517974 253280 517980 253292
rect 517664 253252 517980 253280
rect 517664 253240 517670 253252
rect 517974 253240 517980 253252
rect 518032 253240 518038 253292
rect 179322 253172 179328 253224
rect 179380 253212 179386 253224
rect 197630 253212 197636 253224
rect 179380 253184 197636 253212
rect 179380 253172 179386 253184
rect 197630 253172 197636 253184
rect 197688 253172 197694 253224
rect 351822 253172 351828 253224
rect 351880 253212 351886 253224
rect 360194 253212 360200 253224
rect 351880 253184 360200 253212
rect 351880 253172 351886 253184
rect 360194 253172 360200 253184
rect 360252 253172 360258 253224
rect 517698 253172 517704 253224
rect 517756 253212 517762 253224
rect 518066 253212 518072 253224
rect 517756 253184 518072 253212
rect 517756 253172 517762 253184
rect 518066 253172 518072 253184
rect 518124 253172 518130 253224
rect 191742 252560 191748 252612
rect 191800 252600 191806 252612
rect 198642 252600 198648 252612
rect 191800 252572 198648 252600
rect 191800 252560 191806 252572
rect 198642 252560 198648 252572
rect 198700 252560 198706 252612
rect 510890 252560 510896 252612
rect 510948 252600 510954 252612
rect 517514 252600 517520 252612
rect 510948 252572 517520 252600
rect 510948 252560 510954 252572
rect 517514 252560 517520 252572
rect 517572 252560 517578 252612
rect 217962 252492 217968 252544
rect 218020 252532 218026 252544
rect 265618 252532 265624 252544
rect 218020 252504 265624 252532
rect 218020 252492 218026 252504
rect 265618 252492 265624 252504
rect 265676 252492 265682 252544
rect 218422 252424 218428 252476
rect 218480 252464 218486 252476
rect 219250 252464 219256 252476
rect 218480 252436 219256 252464
rect 218480 252424 218486 252436
rect 219250 252424 219256 252436
rect 219308 252464 219314 252476
rect 264974 252464 264980 252476
rect 219308 252436 264980 252464
rect 219308 252424 219314 252436
rect 264974 252424 264980 252436
rect 265032 252424 265038 252476
rect 58710 252016 58716 252068
rect 58768 252056 58774 252068
rect 60826 252056 60832 252068
rect 58768 252028 60832 252056
rect 58768 252016 58774 252028
rect 60826 252016 60832 252028
rect 60884 252016 60890 252068
rect 216122 252016 216128 252068
rect 216180 252056 216186 252068
rect 229094 252056 229100 252068
rect 216180 252028 229100 252056
rect 216180 252016 216186 252028
rect 229094 252016 229100 252028
rect 229152 252016 229158 252068
rect 379146 252016 379152 252068
rect 379204 252056 379210 252068
rect 396718 252056 396724 252068
rect 379204 252028 396724 252056
rect 379204 252016 379210 252028
rect 396718 252016 396724 252028
rect 396776 252016 396782 252068
rect 58526 251948 58532 252000
rect 58584 251988 58590 252000
rect 83458 251988 83464 252000
rect 58584 251960 83464 251988
rect 58584 251948 58590 251960
rect 83458 251948 83464 251960
rect 83516 251948 83522 252000
rect 216214 251948 216220 252000
rect 216272 251988 216278 252000
rect 230474 251988 230480 252000
rect 216272 251960 230480 251988
rect 216272 251948 216278 251960
rect 230474 251948 230480 251960
rect 230532 251948 230538 252000
rect 372430 251948 372436 252000
rect 372488 251988 372494 252000
rect 376386 251988 376392 252000
rect 372488 251960 376392 251988
rect 372488 251948 372494 251960
rect 376386 251948 376392 251960
rect 376444 251988 376450 252000
rect 425698 251988 425704 252000
rect 376444 251960 425704 251988
rect 376444 251948 376450 251960
rect 425698 251948 425704 251960
rect 425756 251948 425762 252000
rect 68370 251880 68376 251932
rect 68428 251920 68434 251932
rect 96614 251920 96620 251932
rect 68428 251892 96620 251920
rect 68428 251880 68434 251892
rect 96614 251880 96620 251892
rect 96672 251880 96678 251932
rect 218606 251880 218612 251932
rect 218664 251920 218670 251932
rect 233234 251920 233240 251932
rect 218664 251892 233240 251920
rect 218664 251880 218670 251892
rect 233234 251880 233240 251892
rect 233292 251880 233298 251932
rect 368382 251880 368388 251932
rect 368440 251920 368446 251932
rect 371142 251920 371148 251932
rect 368440 251892 371148 251920
rect 368440 251880 368446 251892
rect 371142 251880 371148 251892
rect 371200 251920 371206 251932
rect 421558 251920 421564 251932
rect 371200 251892 421564 251920
rect 371200 251880 371206 251892
rect 421558 251880 421564 251892
rect 421616 251880 421622 251932
rect 53834 251812 53840 251864
rect 53892 251852 53898 251864
rect 102778 251852 102784 251864
rect 53892 251824 102784 251852
rect 53892 251812 53898 251824
rect 102778 251812 102784 251824
rect 102836 251812 102842 251864
rect 216030 251812 216036 251864
rect 216088 251852 216094 251864
rect 218514 251852 218520 251864
rect 216088 251824 218520 251852
rect 216088 251812 216094 251824
rect 218514 251812 218520 251824
rect 218572 251852 218578 251864
rect 264238 251852 264244 251864
rect 218572 251824 264244 251852
rect 218572 251812 218578 251824
rect 264238 251812 264244 251824
rect 264296 251812 264302 251864
rect 343542 251812 343548 251864
rect 343600 251852 343606 251864
rect 360286 251852 360292 251864
rect 343600 251824 360292 251852
rect 343600 251812 343606 251824
rect 360286 251812 360292 251824
rect 360344 251812 360350 251864
rect 369670 251812 369676 251864
rect 369728 251852 369734 251864
rect 371050 251852 371056 251864
rect 369728 251824 371056 251852
rect 369728 251812 369734 251824
rect 371050 251812 371056 251824
rect 371108 251852 371114 251864
rect 422938 251852 422944 251864
rect 371108 251824 422944 251852
rect 371108 251812 371114 251824
rect 422938 251812 422944 251824
rect 422996 251812 423002 251864
rect 49142 250452 49148 250504
rect 49200 250492 49206 250504
rect 54846 250492 54852 250504
rect 49200 250464 54852 250492
rect 49200 250452 49206 250464
rect 54846 250452 54852 250464
rect 54904 250492 54910 250504
rect 68370 250492 68376 250504
rect 54904 250464 68376 250492
rect 54904 250452 54910 250464
rect 68370 250452 68376 250464
rect 68428 250452 68434 250504
rect 519354 183540 519360 183592
rect 519412 183580 519418 183592
rect 520182 183580 520188 183592
rect 519412 183552 520188 183580
rect 519412 183540 519418 183552
rect 520182 183540 520188 183552
rect 520240 183580 520246 183592
rect 580258 183580 580264 183592
rect 520240 183552 580264 183580
rect 520240 183540 520246 183552
rect 580258 183540 580264 183552
rect 580316 183540 580322 183592
rect 520090 183472 520096 183524
rect 520148 183512 520154 183524
rect 580350 183512 580356 183524
rect 520148 183484 580356 183512
rect 520148 183472 520154 183484
rect 580350 183472 580356 183484
rect 580408 183472 580414 183524
rect 209406 177964 209412 178016
rect 209464 178004 209470 178016
rect 216674 178004 216680 178016
rect 209464 177976 216680 178004
rect 209464 177964 209470 177976
rect 216674 177964 216680 177976
rect 216732 177964 216738 178016
rect 365346 177964 365352 178016
rect 365404 178004 365410 178016
rect 377030 178004 377036 178016
rect 365404 177976 377036 178004
rect 365404 177964 365410 177976
rect 377030 177964 377036 177976
rect 377088 177964 377094 178016
rect 360194 176604 360200 176656
rect 360252 176644 360258 176656
rect 376938 176644 376944 176656
rect 360252 176616 376944 176644
rect 360252 176604 360258 176616
rect 376938 176604 376944 176616
rect 376996 176604 377002 176656
rect 358722 176128 358728 176180
rect 358780 176168 358786 176180
rect 360194 176168 360200 176180
rect 358780 176140 360200 176168
rect 358780 176128 358786 176140
rect 360194 176128 360200 176140
rect 360252 176128 360258 176180
rect 197998 175924 198004 175976
rect 198056 175964 198062 175976
rect 198642 175964 198648 175976
rect 198056 175936 198648 175964
rect 198056 175924 198062 175936
rect 198642 175924 198648 175936
rect 198700 175964 198706 175976
rect 216674 175964 216680 175976
rect 198700 175936 216680 175964
rect 198700 175924 198706 175936
rect 216674 175924 216680 175936
rect 216732 175924 216738 175976
rect 204990 175176 204996 175228
rect 205048 175216 205054 175228
rect 216674 175216 216680 175228
rect 205048 175188 216680 175216
rect 205048 175176 205054 175188
rect 216674 175176 216680 175188
rect 216732 175176 216738 175228
rect 362402 175176 362408 175228
rect 362460 175216 362466 175228
rect 377214 175216 377220 175228
rect 362460 175188 377220 175216
rect 362460 175176 362466 175188
rect 377214 175176 377220 175188
rect 377272 175176 377278 175228
rect 52086 166948 52092 167000
rect 52144 166988 52150 167000
rect 101030 166988 101036 167000
rect 52144 166960 101036 166988
rect 52144 166948 52150 166960
rect 101030 166948 101036 166960
rect 101088 166948 101094 167000
rect 366634 166948 366640 167000
rect 366692 166988 366698 167000
rect 423398 166988 423404 167000
rect 366692 166960 423404 166988
rect 366692 166948 366698 166960
rect 423398 166948 423404 166960
rect 423456 166948 423462 167000
rect 49326 166880 49332 166932
rect 49384 166920 49390 166932
rect 98454 166920 98460 166932
rect 49384 166892 98460 166920
rect 49384 166880 49390 166892
rect 98454 166880 98460 166892
rect 98512 166880 98518 166932
rect 358262 166880 358268 166932
rect 358320 166920 358326 166932
rect 416038 166920 416044 166932
rect 358320 166892 416044 166920
rect 358320 166880 358326 166892
rect 416038 166880 416044 166892
rect 416096 166880 416102 166932
rect 52270 166812 52276 166864
rect 52328 166852 52334 166864
rect 105814 166852 105820 166864
rect 52328 166824 105820 166852
rect 52328 166812 52334 166824
rect 105814 166812 105820 166824
rect 105872 166812 105878 166864
rect 202230 166812 202236 166864
rect 202288 166852 202294 166864
rect 253566 166852 253572 166864
rect 202288 166824 253572 166852
rect 202288 166812 202294 166824
rect 253566 166812 253572 166824
rect 253624 166812 253630 166864
rect 356698 166812 356704 166864
rect 356756 166852 356762 166864
rect 418430 166852 418436 166864
rect 356756 166824 418436 166852
rect 356756 166812 356762 166824
rect 418430 166812 418436 166824
rect 418488 166812 418494 166864
rect 50706 166744 50712 166796
rect 50764 166784 50770 166796
rect 108206 166784 108212 166796
rect 50764 166756 108212 166784
rect 50764 166744 50770 166756
rect 108206 166744 108212 166756
rect 108264 166744 108270 166796
rect 209222 166744 209228 166796
rect 209280 166784 209286 166796
rect 270862 166784 270868 166796
rect 209280 166756 270868 166784
rect 209280 166744 209286 166756
rect 270862 166744 270868 166756
rect 270920 166744 270926 166796
rect 356790 166744 356796 166796
rect 356848 166784 356854 166796
rect 425974 166784 425980 166796
rect 356848 166756 425980 166784
rect 356848 166744 356854 166756
rect 425974 166744 425980 166756
rect 426032 166744 426038 166796
rect 56226 166676 56232 166728
rect 56284 166716 56290 166728
rect 138474 166716 138480 166728
rect 56284 166688 138480 166716
rect 56284 166676 56290 166688
rect 138474 166676 138480 166688
rect 138532 166676 138538 166728
rect 202414 166676 202420 166728
rect 202472 166716 202478 166728
rect 265894 166716 265900 166728
rect 202472 166688 265900 166716
rect 202472 166676 202478 166688
rect 265894 166676 265900 166688
rect 265952 166676 265958 166728
rect 370774 166676 370780 166728
rect 370832 166716 370838 166728
rect 473446 166716 473452 166728
rect 370832 166688 473452 166716
rect 370832 166676 370838 166688
rect 473446 166676 473452 166688
rect 473504 166676 473510 166728
rect 59814 166608 59820 166660
rect 59872 166648 59878 166660
rect 143534 166648 143540 166660
rect 59872 166620 143540 166648
rect 59872 166608 59878 166620
rect 143534 166608 143540 166620
rect 143592 166608 143598 166660
rect 206370 166608 206376 166660
rect 206428 166648 206434 166660
rect 288250 166648 288256 166660
rect 206428 166620 288256 166648
rect 206428 166608 206434 166620
rect 288250 166608 288256 166620
rect 288308 166608 288314 166660
rect 367830 166608 367836 166660
rect 367888 166648 367894 166660
rect 475838 166648 475844 166660
rect 367888 166620 475844 166648
rect 367888 166608 367894 166620
rect 475838 166608 475844 166620
rect 475896 166608 475902 166660
rect 59078 166540 59084 166592
rect 59136 166580 59142 166592
rect 145926 166580 145932 166592
rect 59136 166552 145932 166580
rect 59136 166540 59142 166552
rect 145926 166540 145932 166552
rect 145984 166540 145990 166592
rect 209314 166540 209320 166592
rect 209372 166580 209378 166592
rect 298462 166580 298468 166592
rect 209372 166552 298468 166580
rect 209372 166540 209378 166552
rect 298462 166540 298468 166552
rect 298520 166540 298526 166592
rect 369302 166540 369308 166592
rect 369360 166580 369366 166592
rect 478414 166580 478420 166592
rect 369360 166552 478420 166580
rect 369360 166540 369366 166552
rect 478414 166540 478420 166552
rect 478472 166540 478478 166592
rect 59906 166472 59912 166524
rect 59964 166512 59970 166524
rect 150894 166512 150900 166524
rect 59964 166484 150900 166512
rect 59964 166472 59970 166484
rect 150894 166472 150900 166484
rect 150952 166472 150958 166524
rect 211982 166472 211988 166524
rect 212040 166512 212046 166524
rect 303522 166512 303528 166524
rect 212040 166484 303528 166512
rect 212040 166472 212046 166484
rect 303522 166472 303528 166484
rect 303580 166472 303586 166524
rect 371970 166472 371976 166524
rect 372028 166512 372034 166524
rect 480898 166512 480904 166524
rect 372028 166484 480904 166512
rect 372028 166472 372034 166484
rect 480898 166472 480904 166484
rect 480956 166472 480962 166524
rect 58986 166404 58992 166456
rect 59044 166444 59050 166456
rect 153286 166444 153292 166456
rect 59044 166416 153292 166444
rect 59044 166404 59050 166416
rect 153286 166404 153292 166416
rect 153344 166404 153350 166456
rect 203610 166404 203616 166456
rect 203668 166444 203674 166456
rect 295886 166444 295892 166456
rect 203668 166416 295892 166444
rect 203668 166404 203674 166416
rect 295886 166404 295892 166416
rect 295944 166404 295950 166456
rect 361114 166404 361120 166456
rect 361172 166444 361178 166456
rect 470962 166444 470968 166456
rect 361172 166416 470968 166444
rect 361172 166404 361178 166416
rect 470962 166404 470968 166416
rect 471020 166404 471026 166456
rect 42702 166336 42708 166388
rect 42760 166376 42766 166388
rect 163314 166376 163320 166388
rect 42760 166348 163320 166376
rect 42760 166336 42766 166348
rect 163314 166336 163320 166348
rect 163372 166336 163378 166388
rect 213454 166336 213460 166388
rect 213512 166376 213518 166388
rect 308490 166376 308496 166388
rect 213512 166348 308496 166376
rect 213512 166336 213518 166348
rect 308490 166336 308496 166348
rect 308548 166336 308554 166388
rect 373350 166336 373356 166388
rect 373408 166376 373414 166388
rect 485958 166376 485964 166388
rect 373408 166348 485964 166376
rect 373408 166336 373414 166348
rect 485958 166336 485964 166348
rect 486016 166336 486022 166388
rect 41138 166268 41144 166320
rect 41196 166308 41202 166320
rect 165890 166308 165896 166320
rect 41196 166280 165896 166308
rect 41196 166268 41202 166280
rect 165890 166268 165896 166280
rect 165948 166268 165954 166320
rect 214742 166268 214748 166320
rect 214800 166308 214806 166320
rect 315850 166308 315856 166320
rect 214800 166280 315856 166308
rect 214800 166268 214806 166280
rect 315850 166268 315856 166280
rect 315908 166268 315914 166320
rect 365254 166268 365260 166320
rect 365312 166308 365318 166320
rect 483382 166308 483388 166320
rect 365312 166280 483388 166308
rect 365312 166268 365318 166280
rect 483382 166268 483388 166280
rect 483440 166268 483446 166320
rect 50798 166200 50804 166252
rect 50856 166240 50862 166252
rect 96062 166240 96068 166252
rect 50856 166212 96068 166240
rect 50856 166200 50862 166212
rect 96062 166200 96068 166212
rect 96120 166200 96126 166252
rect 374914 166200 374920 166252
rect 374972 166240 374978 166252
rect 428182 166240 428188 166252
rect 374972 166212 428188 166240
rect 374972 166200 374978 166212
rect 428182 166200 428188 166212
rect 428240 166200 428246 166252
rect 365162 166132 365168 166184
rect 365220 166172 365226 166184
rect 408126 166172 408132 166184
rect 365220 166144 408132 166172
rect 365220 166132 365226 166144
rect 408126 166132 408132 166144
rect 408184 166132 408190 166184
rect 370406 166064 370412 166116
rect 370464 166104 370470 166116
rect 380894 166104 380900 166116
rect 370464 166076 380900 166104
rect 370464 166064 370470 166076
rect 380894 166064 380900 166076
rect 380952 166064 380958 166116
rect 54386 165588 54392 165640
rect 54444 165628 54450 165640
rect 113266 165628 113272 165640
rect 54444 165600 113272 165628
rect 54444 165588 54450 165600
rect 113266 165588 113272 165600
rect 113324 165588 113330 165640
rect 55858 165520 55864 165572
rect 55916 165560 55922 165572
rect 132494 165560 132500 165572
rect 55916 165532 132500 165560
rect 55916 165520 55922 165532
rect 132494 165520 132500 165532
rect 132552 165520 132558 165572
rect 211890 165520 211896 165572
rect 211948 165560 211954 165572
rect 310974 165560 310980 165572
rect 211948 165532 310980 165560
rect 211948 165520 211954 165532
rect 310974 165520 310980 165532
rect 311032 165520 311038 165572
rect 343266 165520 343272 165572
rect 343324 165560 343330 165572
rect 357066 165560 357072 165572
rect 343324 165532 357072 165560
rect 343324 165520 343330 165532
rect 357066 165520 357072 165532
rect 357124 165560 357130 165572
rect 357526 165560 357532 165572
rect 357124 165532 357532 165560
rect 357124 165520 357130 165532
rect 357526 165520 357532 165532
rect 357584 165520 357590 165572
rect 362310 165520 362316 165572
rect 362368 165560 362374 165572
rect 452654 165560 452660 165572
rect 362368 165532 452660 165560
rect 362368 165520 362374 165532
rect 452654 165520 452660 165532
rect 452712 165520 452718 165572
rect 55122 165452 55128 165504
rect 55180 165492 55186 165504
rect 129734 165492 129740 165504
rect 55180 165464 129740 165492
rect 55180 165452 55186 165464
rect 129734 165452 129740 165464
rect 129792 165452 129798 165504
rect 210510 165452 210516 165504
rect 210568 165492 210574 165504
rect 293310 165492 293316 165504
rect 210568 165464 293316 165492
rect 210568 165452 210574 165464
rect 293310 165452 293316 165464
rect 293368 165452 293374 165504
rect 369210 165452 369216 165504
rect 369268 165492 369274 165504
rect 455414 165492 455420 165504
rect 369268 165464 455420 165492
rect 369268 165452 369274 165464
rect 455414 165452 455420 165464
rect 455472 165452 455478 165504
rect 55950 165384 55956 165436
rect 56008 165424 56014 165436
rect 128354 165424 128360 165436
rect 56008 165396 128360 165424
rect 56008 165384 56014 165396
rect 128354 165384 128360 165396
rect 128412 165384 128418 165436
rect 219066 165384 219072 165436
rect 219124 165424 219130 165436
rect 300854 165424 300860 165436
rect 219124 165396 300860 165424
rect 219124 165384 219130 165396
rect 300854 165384 300860 165396
rect 300912 165384 300918 165436
rect 358354 165384 358360 165436
rect 358412 165424 358418 165436
rect 442994 165424 443000 165436
rect 358412 165396 443000 165424
rect 358412 165384 358418 165396
rect 442994 165384 443000 165396
rect 443052 165384 443058 165436
rect 54938 165316 54944 165368
rect 54996 165356 55002 165368
rect 125870 165356 125876 165368
rect 54996 165328 125876 165356
rect 54996 165316 55002 165328
rect 125870 165316 125876 165328
rect 125928 165316 125934 165368
rect 213362 165316 213368 165368
rect 213420 165356 213426 165368
rect 285950 165356 285956 165368
rect 213420 165328 285956 165356
rect 213420 165316 213426 165328
rect 285950 165316 285956 165328
rect 286008 165316 286014 165368
rect 370590 165316 370596 165368
rect 370648 165356 370654 165368
rect 449894 165356 449900 165368
rect 370648 165328 449900 165356
rect 370648 165316 370654 165328
rect 449894 165316 449900 165328
rect 449952 165316 449958 165368
rect 56134 165248 56140 165300
rect 56192 165288 56198 165300
rect 123478 165288 123484 165300
rect 56192 165260 123484 165288
rect 56192 165248 56198 165260
rect 123478 165248 123484 165260
rect 123536 165248 123542 165300
rect 211798 165248 211804 165300
rect 211856 165288 211862 165300
rect 276014 165288 276020 165300
rect 211856 165260 276020 165288
rect 211856 165248 211862 165260
rect 276014 165248 276020 165260
rect 276072 165248 276078 165300
rect 378962 165248 378968 165300
rect 379020 165288 379026 165300
rect 458358 165288 458364 165300
rect 379020 165260 458364 165288
rect 379020 165248 379026 165260
rect 458358 165248 458364 165260
rect 458416 165248 458422 165300
rect 53374 165180 53380 165232
rect 53432 165220 53438 165232
rect 120902 165220 120908 165232
rect 53432 165192 120908 165220
rect 53432 165180 53438 165192
rect 120902 165180 120908 165192
rect 120960 165180 120966 165232
rect 214650 165180 214656 165232
rect 214708 165220 214714 165232
rect 278406 165220 278412 165232
rect 214708 165192 278412 165220
rect 214708 165180 214714 165192
rect 278406 165180 278412 165192
rect 278464 165180 278470 165232
rect 371878 165180 371884 165232
rect 371936 165220 371942 165232
rect 447318 165220 447324 165232
rect 371936 165192 447324 165220
rect 371936 165180 371942 165192
rect 447318 165180 447324 165192
rect 447376 165180 447382 165232
rect 56870 165112 56876 165164
rect 56928 165152 56934 165164
rect 57330 165152 57336 165164
rect 56928 165124 57336 165152
rect 56928 165112 56934 165124
rect 57330 165112 57336 165124
rect 57388 165112 57394 165164
rect 59814 165112 59820 165164
rect 59872 165152 59878 165164
rect 115934 165152 115940 165164
rect 59872 165124 115940 165152
rect 59872 165112 59878 165124
rect 115934 165112 115940 165124
rect 115992 165112 115998 165164
rect 183186 165112 183192 165164
rect 183244 165152 183250 165164
rect 197354 165152 197360 165164
rect 183244 165124 197360 165152
rect 183244 165112 183250 165124
rect 197354 165112 197360 165124
rect 197412 165112 197418 165164
rect 218882 165112 218888 165164
rect 218940 165152 218946 165164
rect 280798 165152 280804 165164
rect 218940 165124 280804 165152
rect 218940 165112 218946 165124
rect 280798 165112 280804 165124
rect 280856 165112 280862 165164
rect 366542 165112 366548 165164
rect 366600 165152 366606 165164
rect 440234 165152 440240 165164
rect 366600 165124 440240 165152
rect 366600 165112 366606 165124
rect 440234 165112 440240 165124
rect 440292 165112 440298 165164
rect 503622 165112 503628 165164
rect 503680 165152 503686 165164
rect 517790 165152 517796 165164
rect 503680 165124 517796 165152
rect 503680 165112 503686 165124
rect 517790 165112 517796 165124
rect 517848 165112 517854 165164
rect 55030 165044 55036 165096
rect 55088 165084 55094 165096
rect 118326 165084 118332 165096
rect 55088 165056 118332 165084
rect 55088 165044 55094 165056
rect 118326 165044 118332 165056
rect 118384 165044 118390 165096
rect 204898 165044 204904 165096
rect 204956 165084 204962 165096
rect 263594 165084 263600 165096
rect 204956 165056 263600 165084
rect 204956 165044 204962 165056
rect 263594 165044 263600 165056
rect 263652 165044 263658 165096
rect 361022 165044 361028 165096
rect 361080 165084 361086 165096
rect 422938 165084 422944 165096
rect 361080 165056 422944 165084
rect 361080 165044 361086 165056
rect 422938 165044 422944 165056
rect 422996 165044 423002 165096
rect 517882 165084 517888 165096
rect 509206 165056 517888 165084
rect 53558 164976 53564 165028
rect 53616 165016 53622 165028
rect 113542 165016 113548 165028
rect 53616 164988 113548 165016
rect 53616 164976 53622 164988
rect 113542 164976 113548 164988
rect 113600 164976 113606 165028
rect 183462 164976 183468 165028
rect 183520 165016 183526 165028
rect 201494 165016 201500 165028
rect 183520 164988 201500 165016
rect 183520 164976 183526 164988
rect 201494 164976 201500 164988
rect 201552 164976 201558 165028
rect 215938 164976 215944 165028
rect 215996 165016 216002 165028
rect 273438 165016 273444 165028
rect 215996 164988 273444 165016
rect 215996 164976 216002 164988
rect 273438 164976 273444 164988
rect 273496 164976 273502 165028
rect 373442 164976 373448 165028
rect 373500 165016 373506 165028
rect 445754 165016 445760 165028
rect 373500 164988 445760 165016
rect 373500 164976 373506 164988
rect 445754 164976 445760 164988
rect 445812 164976 445818 165028
rect 503254 164976 503260 165028
rect 503312 165016 503318 165028
rect 509206 165016 509234 165056
rect 517882 165044 517888 165056
rect 517940 165044 517946 165096
rect 516594 165016 516600 165028
rect 503312 164988 509234 165016
rect 510080 164988 516600 165016
rect 503312 164976 503318 164988
rect 51994 164908 52000 164960
rect 52052 164948 52058 164960
rect 59814 164948 59820 164960
rect 52052 164920 59820 164948
rect 52052 164908 52058 164920
rect 59814 164908 59820 164920
rect 59872 164908 59878 164960
rect 59906 164908 59912 164960
rect 59964 164948 59970 164960
rect 103514 164948 103520 164960
rect 59964 164920 103520 164948
rect 59964 164908 59970 164920
rect 103514 164908 103520 164920
rect 103572 164908 103578 164960
rect 116026 164908 116032 164960
rect 116084 164948 116090 164960
rect 196710 164948 196716 164960
rect 116084 164920 196716 164948
rect 116084 164908 116090 164920
rect 196710 164908 196716 164920
rect 196768 164908 196774 164960
rect 210602 164908 210608 164960
rect 210660 164948 210666 164960
rect 267734 164948 267740 164960
rect 210660 164920 267740 164948
rect 210660 164908 210666 164920
rect 267734 164908 267740 164920
rect 267792 164908 267798 164960
rect 363874 164908 363880 164960
rect 363932 164948 363938 164960
rect 434806 164948 434812 164960
rect 363932 164920 434812 164948
rect 363932 164908 363938 164920
rect 434806 164908 434812 164920
rect 434864 164908 434870 164960
rect 440234 164908 440240 164960
rect 440292 164948 440298 164960
rect 510080 164948 510108 164988
rect 516594 164976 516600 164988
rect 516652 164976 516658 165028
rect 440292 164920 510108 164948
rect 440292 164908 440298 164920
rect 510522 164908 510528 164960
rect 510580 164948 510586 164960
rect 517514 164948 517520 164960
rect 510580 164920 517520 164948
rect 510580 164908 510586 164920
rect 517514 164908 517520 164920
rect 517572 164908 517578 164960
rect 57330 164840 57336 164892
rect 57388 164880 57394 164892
rect 104894 164880 104900 164892
rect 57388 164852 104900 164880
rect 57388 164840 57394 164852
rect 104894 164840 104900 164852
rect 104952 164840 104958 164892
rect 114554 164840 114560 164892
rect 114612 164880 114618 164892
rect 196618 164880 196624 164892
rect 114612 164852 196624 164880
rect 114612 164840 114618 164852
rect 196618 164840 196624 164852
rect 196676 164840 196682 164892
rect 207658 164840 207664 164892
rect 207716 164880 207722 164892
rect 258074 164880 258080 164892
rect 207716 164852 258080 164880
rect 207716 164840 207722 164852
rect 258074 164840 258080 164852
rect 258132 164840 258138 164892
rect 343542 164840 343548 164892
rect 343600 164880 343606 164892
rect 360286 164880 360292 164892
rect 343600 164852 360292 164880
rect 343600 164840 343606 164852
rect 360286 164840 360292 164852
rect 360344 164840 360350 164892
rect 369118 164840 369124 164892
rect 369176 164880 369182 164892
rect 437750 164880 437756 164892
rect 369176 164852 437756 164880
rect 369176 164840 369182 164852
rect 437750 164840 437756 164852
rect 437808 164840 437814 164892
rect 50890 164772 50896 164824
rect 50948 164812 50954 164824
rect 59906 164812 59912 164824
rect 50948 164784 59912 164812
rect 50948 164772 50954 164784
rect 59906 164772 59912 164784
rect 59964 164772 59970 164824
rect 89898 164812 89904 164824
rect 60016 164784 89904 164812
rect 49418 164636 49424 164688
rect 49476 164676 49482 164688
rect 60016 164676 60044 164784
rect 89898 164772 89904 164784
rect 89956 164772 89962 164824
rect 206278 164772 206284 164824
rect 206336 164812 206342 164824
rect 255314 164812 255320 164824
rect 206336 164784 255320 164812
rect 206336 164772 206342 164784
rect 255314 164772 255320 164784
rect 255372 164772 255378 164824
rect 378870 164772 378876 164824
rect 378928 164812 378934 164824
rect 420914 164812 420920 164824
rect 378928 164784 420920 164812
rect 378928 164772 378934 164784
rect 420914 164772 420920 164784
rect 420972 164772 420978 164824
rect 422938 164772 422944 164824
rect 422996 164812 423002 164824
rect 433334 164812 433340 164824
rect 422996 164784 433340 164812
rect 422996 164772 423002 164784
rect 433334 164772 433340 164784
rect 433392 164772 433398 164824
rect 88334 164744 88340 164756
rect 49476 164648 60044 164676
rect 64846 164716 88340 164744
rect 49476 164636 49482 164648
rect 56042 164568 56048 164620
rect 56100 164608 56106 164620
rect 64846 164608 64874 164716
rect 88334 164704 88340 164716
rect 88392 164704 88398 164756
rect 209130 164704 209136 164756
rect 209188 164744 209194 164756
rect 249794 164744 249800 164756
rect 209188 164716 249800 164744
rect 209188 164704 209194 164716
rect 249794 164704 249800 164716
rect 249852 164704 249858 164756
rect 378778 164704 378784 164756
rect 378836 164744 378842 164756
rect 413554 164744 413560 164756
rect 378836 164716 413560 164744
rect 378836 164704 378842 164716
rect 413554 164704 413560 164716
rect 413612 164704 413618 164756
rect 214558 164636 214564 164688
rect 214616 164676 214622 164688
rect 247034 164676 247040 164688
rect 214616 164648 247040 164676
rect 214616 164636 214622 164648
rect 247034 164636 247040 164648
rect 247092 164636 247098 164688
rect 376110 164636 376116 164688
rect 376168 164676 376174 164688
rect 410426 164676 410432 164688
rect 376168 164648 410432 164676
rect 376168 164636 376174 164648
rect 410426 164636 410432 164648
rect 410484 164636 410490 164688
rect 56100 164580 64874 164608
rect 56100 164568 56106 164580
rect 428826 164500 428832 164552
rect 428884 164540 428890 164552
rect 433334 164540 433340 164552
rect 428884 164512 433340 164540
rect 428884 164500 428890 164512
rect 433334 164500 433340 164512
rect 433392 164500 433398 164552
rect 83458 164432 83464 164484
rect 83516 164472 83522 164484
rect 107746 164472 107752 164484
rect 83516 164444 107752 164472
rect 83516 164432 83522 164444
rect 107746 164432 107752 164444
rect 107804 164432 107810 164484
rect 97258 164364 97264 164416
rect 97316 164404 97322 164416
rect 100754 164404 100760 164416
rect 97316 164376 100760 164404
rect 97316 164364 97322 164376
rect 100754 164364 100760 164376
rect 100812 164364 100818 164416
rect 88978 164296 88984 164348
rect 89036 164336 89042 164348
rect 106274 164336 106280 164348
rect 89036 164308 106280 164336
rect 89036 164296 89042 164308
rect 106274 164296 106280 164308
rect 106332 164296 106338 164348
rect 269758 164228 269764 164280
rect 269816 164268 269822 164280
rect 273806 164268 273812 164280
rect 269816 164240 273812 164268
rect 269816 164228 269822 164240
rect 273806 164228 273812 164240
rect 273864 164228 273870 164280
rect 47578 164160 47584 164212
rect 47636 164200 47642 164212
rect 52270 164200 52276 164212
rect 47636 164172 52276 164200
rect 47636 164160 47642 164172
rect 52270 164160 52276 164172
rect 52328 164160 52334 164212
rect 54570 164160 54576 164212
rect 54628 164200 54634 164212
rect 57514 164200 57520 164212
rect 54628 164172 57520 164200
rect 54628 164160 54634 164172
rect 57514 164160 57520 164172
rect 57572 164200 57578 164212
rect 116394 164200 116400 164212
rect 57572 164172 116400 164200
rect 57572 164160 57578 164172
rect 116394 164160 116400 164172
rect 116452 164160 116458 164212
rect 214282 164160 214288 164212
rect 214340 164200 214346 164212
rect 215754 164200 215760 164212
rect 214340 164172 215760 164200
rect 214340 164160 214346 164172
rect 215754 164160 215760 164172
rect 215812 164160 215818 164212
rect 219526 164160 219532 164212
rect 219584 164200 219590 164212
rect 219986 164200 219992 164212
rect 219584 164172 219992 164200
rect 219584 164160 219590 164172
rect 219986 164160 219992 164172
rect 220044 164200 220050 164212
rect 267734 164200 267740 164212
rect 220044 164172 267740 164200
rect 220044 164160 220050 164172
rect 267734 164160 267740 164172
rect 267792 164160 267798 164212
rect 377306 164160 377312 164212
rect 377364 164200 377370 164212
rect 437842 164200 437848 164212
rect 377364 164172 437848 164200
rect 377364 164160 377370 164172
rect 437842 164160 437848 164172
rect 437900 164160 437906 164212
rect 55674 164092 55680 164144
rect 55732 164132 55738 164144
rect 59630 164132 59636 164144
rect 55732 164104 59636 164132
rect 55732 164092 55738 164104
rect 59630 164092 59636 164104
rect 59688 164132 59694 164144
rect 117866 164132 117872 164144
rect 59688 164104 117872 164132
rect 59688 164092 59694 164104
rect 117866 164092 117872 164104
rect 117924 164092 117930 164144
rect 370682 164092 370688 164144
rect 370740 164132 370746 164144
rect 430574 164132 430580 164144
rect 370740 164104 430580 164132
rect 370740 164092 370746 164104
rect 430574 164092 430580 164104
rect 430632 164092 430638 164144
rect 53466 164024 53472 164076
rect 53524 164064 53530 164076
rect 110874 164064 110880 164076
rect 53524 164036 110880 164064
rect 53524 164024 53530 164036
rect 110874 164024 110880 164036
rect 110932 164024 110938 164076
rect 376386 164024 376392 164076
rect 376444 164064 376450 164076
rect 429286 164064 429292 164076
rect 376444 164036 429292 164064
rect 376444 164024 376450 164036
rect 429286 164024 429292 164036
rect 429344 164024 429350 164076
rect 53006 163956 53012 164008
rect 53064 163996 53070 164008
rect 109678 163996 109684 164008
rect 53064 163968 109684 163996
rect 53064 163956 53070 163968
rect 109678 163956 109684 163968
rect 109736 163956 109742 164008
rect 379790 163956 379796 164008
rect 379848 163996 379854 164008
rect 426434 163996 426440 164008
rect 379848 163968 426440 163996
rect 379848 163956 379854 163968
rect 426434 163956 426440 163968
rect 426492 163956 426498 164008
rect 379698 163888 379704 163940
rect 379756 163928 379762 163940
rect 425054 163928 425060 163940
rect 379756 163900 425060 163928
rect 379756 163888 379762 163900
rect 425054 163888 425060 163900
rect 425112 163888 425118 163940
rect 379146 163820 379152 163872
rect 379204 163860 379210 163872
rect 416866 163860 416872 163872
rect 379204 163832 416872 163860
rect 379204 163820 379210 163832
rect 416866 163820 416872 163832
rect 416924 163820 416930 163872
rect 59078 163752 59084 163804
rect 59136 163792 59142 163804
rect 95234 163792 95240 163804
rect 59136 163764 95240 163792
rect 59136 163752 59142 163764
rect 95234 163752 95240 163764
rect 95292 163752 95298 163804
rect 374546 163752 374552 163804
rect 374604 163792 374610 163804
rect 396074 163792 396080 163804
rect 374604 163764 396080 163792
rect 374604 163752 374610 163764
rect 396074 163752 396080 163764
rect 396132 163752 396138 163804
rect 50982 163684 50988 163736
rect 51040 163724 51046 163736
rect 55030 163724 55036 163736
rect 51040 163696 55036 163724
rect 51040 163684 51046 163696
rect 55030 163684 55036 163696
rect 55088 163724 55094 163736
rect 97994 163724 98000 163736
rect 55088 163696 98000 163724
rect 55088 163684 55094 163696
rect 97994 163684 98000 163696
rect 98052 163684 98058 163736
rect 217134 163684 217140 163736
rect 217192 163724 217198 163736
rect 219066 163724 219072 163736
rect 217192 163696 219072 163724
rect 217192 163684 217198 163696
rect 219066 163684 219072 163696
rect 219124 163724 219130 163736
rect 263778 163724 263784 163736
rect 219124 163696 263784 163724
rect 219124 163684 219130 163696
rect 263778 163684 263784 163696
rect 263836 163684 263842 163736
rect 374362 163684 374368 163736
rect 374420 163724 374426 163736
rect 396166 163724 396172 163736
rect 374420 163696 396172 163724
rect 374420 163684 374426 163696
rect 396166 163684 396172 163696
rect 396224 163684 396230 163736
rect 52270 163616 52276 163668
rect 52328 163656 52334 163668
rect 111150 163656 111156 163668
rect 52328 163628 111156 163656
rect 52328 163616 52334 163628
rect 111150 163616 111156 163628
rect 111208 163616 111214 163668
rect 215754 163616 215760 163668
rect 215812 163656 215818 163668
rect 262214 163656 262220 163668
rect 215812 163628 262220 163656
rect 215812 163616 215818 163628
rect 262214 163616 262220 163628
rect 262272 163616 262278 163668
rect 50338 163548 50344 163600
rect 50396 163588 50402 163600
rect 53558 163588 53564 163600
rect 50396 163560 53564 163588
rect 50396 163548 50402 163560
rect 53558 163548 53564 163560
rect 53616 163588 53622 163600
rect 111886 163588 111892 163600
rect 53616 163560 111892 163588
rect 53616 163548 53622 163560
rect 111886 163548 111892 163560
rect 111944 163548 111950 163600
rect 220722 163548 220728 163600
rect 220780 163588 220786 163600
rect 266446 163588 266452 163600
rect 220780 163560 266452 163588
rect 220780 163548 220786 163560
rect 266446 163548 266452 163560
rect 266504 163548 266510 163600
rect 375190 163548 375196 163600
rect 375248 163588 375254 163600
rect 430666 163588 430672 163600
rect 375248 163560 430672 163588
rect 375248 163548 375254 163560
rect 430666 163548 430672 163560
rect 430724 163548 430730 163600
rect 52730 163480 52736 163532
rect 52788 163520 52794 163532
rect 59078 163520 59084 163532
rect 52788 163492 59084 163520
rect 52788 163480 52794 163492
rect 59078 163480 59084 163492
rect 59136 163480 59142 163532
rect 59446 163480 59452 163532
rect 59504 163520 59510 163532
rect 118878 163520 118884 163532
rect 59504 163492 118884 163520
rect 59504 163480 59510 163492
rect 118878 163480 118884 163492
rect 118936 163480 118942 163532
rect 218882 163480 218888 163532
rect 218940 163520 218946 163532
rect 219250 163520 219256 163532
rect 218940 163492 219256 163520
rect 218940 163480 218946 163492
rect 219250 163480 219256 163492
rect 219308 163520 219314 163532
rect 266538 163520 266544 163532
rect 219308 163492 266544 163520
rect 219308 163480 219314 163492
rect 266538 163480 266544 163492
rect 266596 163480 266602 163532
rect 371142 163480 371148 163532
rect 371200 163520 371206 163532
rect 375834 163520 375840 163532
rect 371200 163492 375840 163520
rect 371200 163480 371206 163492
rect 375834 163480 375840 163492
rect 375892 163520 375898 163532
rect 436094 163520 436100 163532
rect 375892 163492 436100 163520
rect 375892 163480 375898 163492
rect 436094 163480 436100 163492
rect 436152 163480 436158 163532
rect 372154 163140 372160 163192
rect 372212 163180 372218 163192
rect 374270 163180 374276 163192
rect 372212 163152 374276 163180
rect 372212 163140 372218 163152
rect 374270 163140 374276 163152
rect 374328 163180 374334 163192
rect 375190 163180 375196 163192
rect 374328 163152 375196 163180
rect 374328 163140 374334 163152
rect 375190 163140 375196 163152
rect 375248 163140 375254 163192
rect 218514 162936 218520 162988
rect 218572 162976 218578 162988
rect 219526 162976 219532 162988
rect 218572 162948 219532 162976
rect 218572 162936 218578 162948
rect 219526 162936 219532 162948
rect 219584 162976 219590 162988
rect 220722 162976 220728 162988
rect 219584 162948 220728 162976
rect 219584 162936 219590 162948
rect 220722 162936 220728 162948
rect 220780 162936 220786 162988
rect 217226 162800 217232 162852
rect 217284 162840 217290 162852
rect 217962 162840 217968 162852
rect 217284 162812 217968 162840
rect 217284 162800 217290 162812
rect 217962 162800 217968 162812
rect 218020 162800 218026 162852
rect 260834 162840 260840 162852
rect 218072 162812 260840 162840
rect 216122 162732 216128 162784
rect 216180 162772 216186 162784
rect 218072 162772 218100 162812
rect 260834 162800 260840 162812
rect 260892 162800 260898 162852
rect 375098 162800 375104 162852
rect 375156 162840 375162 162852
rect 379606 162840 379612 162852
rect 375156 162812 379612 162840
rect 375156 162800 375162 162812
rect 379606 162800 379612 162812
rect 379664 162800 379670 162852
rect 434806 162840 434812 162852
rect 379716 162812 434812 162840
rect 259546 162772 259552 162784
rect 216180 162744 218100 162772
rect 218532 162744 259552 162772
rect 216180 162732 216186 162744
rect 214650 162528 214656 162580
rect 214708 162568 214714 162580
rect 216214 162568 216220 162580
rect 214708 162540 216220 162568
rect 214708 162528 214714 162540
rect 216214 162528 216220 162540
rect 216272 162568 216278 162580
rect 218532 162568 218560 162744
rect 259546 162732 259552 162744
rect 259604 162732 259610 162784
rect 375006 162732 375012 162784
rect 375064 162772 375070 162784
rect 379716 162772 379744 162812
rect 434806 162800 434812 162812
rect 434864 162800 434870 162852
rect 375064 162744 379744 162772
rect 375064 162732 375070 162744
rect 379882 162732 379888 162784
rect 379940 162772 379946 162784
rect 428826 162772 428832 162784
rect 379940 162744 428832 162772
rect 379940 162732 379946 162744
rect 428826 162732 428832 162744
rect 428884 162732 428890 162784
rect 218882 162664 218888 162716
rect 218940 162704 218946 162716
rect 259454 162704 259460 162716
rect 218940 162676 259460 162704
rect 218940 162664 218946 162676
rect 259454 162664 259460 162676
rect 259512 162664 259518 162716
rect 374454 162664 374460 162716
rect 374512 162704 374518 162716
rect 420914 162704 420920 162716
rect 374512 162676 420920 162704
rect 374512 162664 374518 162676
rect 420914 162664 420920 162676
rect 420972 162664 420978 162716
rect 218606 162596 218612 162648
rect 218664 162636 218670 162648
rect 258166 162636 258172 162648
rect 218664 162608 258172 162636
rect 218664 162596 218670 162608
rect 258166 162596 258172 162608
rect 258224 162596 258230 162648
rect 419534 162636 419540 162648
rect 383626 162608 419540 162636
rect 216272 162540 218560 162568
rect 216272 162528 216278 162540
rect 376754 162460 376760 162512
rect 376812 162500 376818 162512
rect 378042 162500 378048 162512
rect 376812 162472 378048 162500
rect 376812 162460 376818 162472
rect 378042 162460 378048 162472
rect 378100 162460 378106 162512
rect 378134 162460 378140 162512
rect 378192 162500 378198 162512
rect 383626 162500 383654 162608
rect 419534 162596 419540 162608
rect 419592 162596 419598 162648
rect 378192 162472 383654 162500
rect 378192 162460 378198 162472
rect 376478 162392 376484 162444
rect 376536 162432 376542 162444
rect 379882 162432 379888 162444
rect 376536 162404 379888 162432
rect 376536 162392 376542 162404
rect 379882 162392 379888 162404
rect 379940 162392 379946 162444
rect 379606 162188 379612 162240
rect 379664 162228 379670 162240
rect 418246 162228 418252 162240
rect 379664 162200 418252 162228
rect 379664 162188 379670 162200
rect 418246 162188 418252 162200
rect 418304 162188 418310 162240
rect 220170 162120 220176 162172
rect 220228 162160 220234 162172
rect 256694 162160 256700 162172
rect 220228 162132 256700 162160
rect 220228 162120 220234 162132
rect 256694 162120 256700 162132
rect 256752 162120 256758 162172
rect 373534 162120 373540 162172
rect 373592 162160 373598 162172
rect 375190 162160 375196 162172
rect 373592 162132 375196 162160
rect 373592 162120 373598 162132
rect 375190 162120 375196 162132
rect 375248 162160 375254 162172
rect 431954 162160 431960 162172
rect 375248 162132 431960 162160
rect 375248 162120 375254 162132
rect 431954 162120 431960 162132
rect 432012 162120 432018 162172
rect 214742 161848 214748 161900
rect 214800 161888 214806 161900
rect 216674 161888 216680 161900
rect 214800 161860 216680 161888
rect 214800 161848 214806 161860
rect 216674 161848 216680 161860
rect 216732 161848 216738 161900
rect 378042 161508 378048 161560
rect 378100 161548 378106 161560
rect 395338 161548 395344 161560
rect 378100 161520 395344 161548
rect 378100 161508 378106 161520
rect 395338 161508 395344 161520
rect 395396 161508 395402 161560
rect 217962 161440 217968 161492
rect 218020 161480 218026 161492
rect 235258 161480 235264 161492
rect 218020 161452 235264 161480
rect 218020 161440 218026 161452
rect 235258 161440 235264 161452
rect 235316 161440 235322 161492
rect 376662 161440 376668 161492
rect 376720 161480 376726 161492
rect 396718 161480 396724 161492
rect 376720 161452 396724 161480
rect 376720 161440 376726 161452
rect 396718 161440 396724 161452
rect 396776 161440 396782 161492
rect 205542 161372 205548 161424
rect 205600 161412 205606 161424
rect 220170 161412 220176 161424
rect 205600 161384 220176 161412
rect 205600 161372 205606 161384
rect 220170 161372 220176 161384
rect 220228 161372 220234 161424
rect 219802 156612 219808 156664
rect 219860 156652 219866 156664
rect 220078 156652 220084 156664
rect 219860 156624 220084 156652
rect 219860 156612 219866 156624
rect 220078 156612 220084 156624
rect 220136 156612 220142 156664
rect 219434 156476 219440 156528
rect 219492 156516 219498 156528
rect 219802 156516 219808 156528
rect 219492 156488 219808 156516
rect 219492 156476 219498 156488
rect 219802 156476 219808 156488
rect 219860 156476 219866 156528
rect 219434 156340 219440 156392
rect 219492 156380 219498 156392
rect 220170 156380 220176 156392
rect 219492 156352 220176 156380
rect 219492 156340 219498 156352
rect 220170 156340 220176 156352
rect 220228 156340 220234 156392
rect 57974 148996 57980 149048
rect 58032 149036 58038 149048
rect 103606 149036 103612 149048
rect 58032 149008 103612 149036
rect 58032 148996 58038 149008
rect 103606 148996 103612 149008
rect 103664 148996 103670 149048
rect 212810 148996 212816 149048
rect 212868 149036 212874 149048
rect 274634 149036 274640 149048
rect 212868 149008 274640 149036
rect 212868 148996 212874 149008
rect 274634 148996 274640 149008
rect 274692 148996 274698 149048
rect 274726 148996 274732 149048
rect 274784 149036 274790 149048
rect 275278 149036 275284 149048
rect 274784 149008 275284 149036
rect 274784 148996 274790 149008
rect 275278 148996 275284 149008
rect 275336 149036 275342 149048
rect 356882 149036 356888 149048
rect 275336 149008 356888 149036
rect 275336 148996 275342 149008
rect 356882 148996 356888 149008
rect 356940 148996 356946 149048
rect 379514 148996 379520 149048
rect 379572 149036 379578 149048
rect 412726 149036 412732 149048
rect 379572 149008 412732 149036
rect 379572 148996 379578 149008
rect 412726 148996 412732 149008
rect 412784 148996 412790 149048
rect 58802 148928 58808 148980
rect 58860 148968 58866 148980
rect 102134 148968 102140 148980
rect 58860 148940 102140 148968
rect 58860 148928 58866 148940
rect 102134 148928 102140 148940
rect 102192 148928 102198 148980
rect 212166 148928 212172 148980
rect 212224 148968 212230 148980
rect 269758 148968 269764 148980
rect 212224 148940 269764 148968
rect 212224 148928 212230 148940
rect 269758 148928 269764 148940
rect 269816 148928 269822 148980
rect 375282 148928 375288 148980
rect 375340 148968 375346 148980
rect 401594 148968 401600 148980
rect 375340 148940 401600 148968
rect 375340 148928 375346 148940
rect 401594 148928 401600 148940
rect 401652 148928 401658 148980
rect 213638 148860 213644 148912
rect 213696 148900 213702 148912
rect 240134 148900 240140 148912
rect 213696 148872 240140 148900
rect 213696 148860 213702 148872
rect 240134 148860 240140 148872
rect 240192 148860 240198 148912
rect 47762 148792 47768 148844
rect 47820 148832 47826 148844
rect 59906 148832 59912 148844
rect 47820 148804 59912 148832
rect 47820 148792 47826 148804
rect 59906 148792 59912 148804
rect 59964 148832 59970 148844
rect 83458 148832 83464 148844
rect 59964 148804 83464 148832
rect 59964 148792 59970 148804
rect 83458 148792 83464 148804
rect 83516 148792 83522 148844
rect 47946 148724 47952 148776
rect 48004 148764 48010 148776
rect 52086 148764 52092 148776
rect 48004 148736 52092 148764
rect 48004 148724 48010 148736
rect 52086 148724 52092 148736
rect 52144 148764 52150 148776
rect 78674 148764 78680 148776
rect 52144 148736 78680 148764
rect 52144 148724 52150 148736
rect 78674 148724 78680 148736
rect 78732 148724 78738 148776
rect 47854 148656 47860 148708
rect 47912 148696 47918 148708
rect 51994 148696 52000 148708
rect 47912 148668 52000 148696
rect 47912 148656 47918 148668
rect 51994 148656 52000 148668
rect 52052 148696 52058 148708
rect 80054 148696 80060 148708
rect 52052 148668 80060 148696
rect 52052 148656 52058 148668
rect 80054 148656 80060 148668
rect 80112 148656 80118 148708
rect 49050 148588 49056 148640
rect 49108 148628 49114 148640
rect 53374 148628 53380 148640
rect 49108 148600 53380 148628
rect 49108 148588 49114 148600
rect 53374 148588 53380 148600
rect 53432 148628 53438 148640
rect 81434 148628 81440 148640
rect 53432 148600 81440 148628
rect 53432 148588 53438 148600
rect 81434 148588 81440 148600
rect 81492 148588 81498 148640
rect 374914 148588 374920 148640
rect 374972 148628 374978 148640
rect 375282 148628 375288 148640
rect 374972 148600 375288 148628
rect 374972 148588 374978 148600
rect 375282 148588 375288 148600
rect 375340 148588 375346 148640
rect 56042 148520 56048 148572
rect 56100 148560 56106 148572
rect 58802 148560 58808 148572
rect 56100 148532 58808 148560
rect 56100 148520 56106 148532
rect 58802 148520 58808 148532
rect 58860 148520 58866 148572
rect 58986 148520 58992 148572
rect 59044 148560 59050 148572
rect 88978 148560 88984 148572
rect 59044 148532 88984 148560
rect 59044 148520 59050 148532
rect 88978 148520 88984 148532
rect 89036 148520 89042 148572
rect 212902 148520 212908 148572
rect 212960 148560 212966 148572
rect 213638 148560 213644 148572
rect 212960 148532 213644 148560
rect 212960 148520 212966 148532
rect 213638 148520 213644 148532
rect 213696 148520 213702 148572
rect 58526 148452 58532 148504
rect 58584 148492 58590 148504
rect 59814 148492 59820 148504
rect 58584 148464 59820 148492
rect 58584 148452 58590 148464
rect 59814 148452 59820 148464
rect 59872 148492 59878 148504
rect 107654 148492 107660 148504
rect 59872 148464 107660 148492
rect 59872 148452 59878 148464
rect 107654 148452 107660 148464
rect 107712 148452 107718 148504
rect 210878 148452 210884 148504
rect 210936 148492 210942 148504
rect 213454 148492 213460 148504
rect 210936 148464 213460 148492
rect 210936 148452 210942 148464
rect 213454 148452 213460 148464
rect 213512 148492 213518 148504
rect 238754 148492 238760 148504
rect 213512 148464 238760 148492
rect 213512 148452 213518 148464
rect 238754 148452 238760 148464
rect 238812 148452 238818 148504
rect 375282 148452 375288 148504
rect 375340 148492 375346 148504
rect 398834 148492 398840 148504
rect 375340 148464 398840 148492
rect 375340 148452 375346 148464
rect 398834 148452 398840 148464
rect 398892 148452 398898 148504
rect 54938 148384 54944 148436
rect 54996 148424 55002 148436
rect 116026 148424 116032 148436
rect 54996 148396 116032 148424
rect 54996 148384 55002 148396
rect 116026 148384 116032 148396
rect 116084 148384 116090 148436
rect 213730 148384 213736 148436
rect 213788 148424 213794 148436
rect 241514 148424 241520 148436
rect 213788 148396 241520 148424
rect 213788 148384 213794 148396
rect 241514 148384 241520 148396
rect 241572 148384 241578 148436
rect 372062 148384 372068 148436
rect 372120 148424 372126 148436
rect 373350 148424 373356 148436
rect 372120 148396 373356 148424
rect 372120 148384 372126 148396
rect 373350 148384 373356 148396
rect 373408 148424 373414 148436
rect 400214 148424 400220 148436
rect 373408 148396 400220 148424
rect 373408 148384 373414 148396
rect 400214 148384 400220 148396
rect 400272 148384 400278 148436
rect 53190 148316 53196 148368
rect 53248 148356 53254 148368
rect 114554 148356 114560 148368
rect 53248 148328 114560 148356
rect 53248 148316 53254 148328
rect 114554 148316 114560 148328
rect 114612 148316 114618 148368
rect 213086 148316 213092 148368
rect 213144 148356 213150 148368
rect 274726 148356 274732 148368
rect 213144 148328 274732 148356
rect 213144 148316 213150 148328
rect 274726 148316 274732 148328
rect 274784 148316 274790 148368
rect 373166 148316 373172 148368
rect 373224 148356 373230 148368
rect 374546 148356 374552 148368
rect 373224 148328 374552 148356
rect 373224 148316 373230 148328
rect 374546 148316 374552 148328
rect 374604 148356 374610 148368
rect 434714 148356 434720 148368
rect 374604 148328 434720 148356
rect 374604 148316 374610 148328
rect 434714 148316 434720 148328
rect 434772 148316 434778 148368
rect 47670 148248 47676 148300
rect 47728 148288 47734 148300
rect 58526 148288 58532 148300
rect 47728 148260 58532 148288
rect 47728 148248 47734 148260
rect 58526 148248 58532 148260
rect 58584 148288 58590 148300
rect 58986 148288 58992 148300
rect 58584 148260 58992 148288
rect 58584 148248 58590 148260
rect 58986 148248 58992 148260
rect 59044 148248 59050 148300
rect 56134 147636 56140 147688
rect 56192 147676 56198 147688
rect 57974 147676 57980 147688
rect 56192 147648 57980 147676
rect 56192 147636 56198 147648
rect 57974 147636 57980 147648
rect 58032 147636 58038 147688
rect 212810 147636 212816 147688
rect 212868 147676 212874 147688
rect 212868 147648 213868 147676
rect 212868 147636 212874 147648
rect 208118 147568 208124 147620
rect 208176 147608 208182 147620
rect 213362 147608 213368 147620
rect 208176 147580 213368 147608
rect 208176 147568 208182 147580
rect 213362 147568 213368 147580
rect 213420 147608 213426 147620
rect 213730 147608 213736 147620
rect 213420 147580 213736 147608
rect 213420 147568 213426 147580
rect 213730 147568 213736 147580
rect 213788 147568 213794 147620
rect 213840 147540 213868 147648
rect 379330 147636 379336 147688
rect 379388 147676 379394 147688
rect 379514 147676 379520 147688
rect 379388 147648 379520 147676
rect 379388 147636 379394 147648
rect 379514 147636 379520 147648
rect 379572 147636 379578 147688
rect 213748 147512 213868 147540
rect 213748 147484 213776 147512
rect 368290 147500 368296 147552
rect 368348 147540 368354 147552
rect 374822 147540 374828 147552
rect 368348 147512 374828 147540
rect 368348 147500 368354 147512
rect 374822 147500 374828 147512
rect 374880 147540 374886 147552
rect 375282 147540 375288 147552
rect 374880 147512 375288 147540
rect 374880 147500 374886 147512
rect 375282 147500 375288 147512
rect 375340 147500 375346 147552
rect 213730 147432 213736 147484
rect 213788 147432 213794 147484
rect 60090 146316 60096 146328
rect 58912 146288 60096 146316
rect 58912 146260 58940 146288
rect 60090 146276 60096 146288
rect 60148 146276 60154 146328
rect 215846 146276 215852 146328
rect 215904 146316 215910 146328
rect 277394 146316 277400 146328
rect 215904 146288 277400 146316
rect 215904 146276 215910 146288
rect 277366 146276 277400 146288
rect 277452 146276 277458 146328
rect 46658 146208 46664 146260
rect 46716 146248 46722 146260
rect 51902 146248 51908 146260
rect 46716 146220 51908 146248
rect 46716 146208 46722 146220
rect 51902 146208 51908 146220
rect 51960 146208 51966 146260
rect 55766 146208 55772 146260
rect 55824 146248 55830 146260
rect 56226 146248 56232 146260
rect 55824 146220 56232 146248
rect 55824 146208 55830 146220
rect 56226 146208 56232 146220
rect 56284 146208 56290 146260
rect 58618 146208 58624 146260
rect 58676 146248 58682 146260
rect 58894 146248 58900 146260
rect 58676 146220 58900 146248
rect 58676 146208 58682 146220
rect 58894 146208 58900 146220
rect 58952 146208 58958 146260
rect 58986 146208 58992 146260
rect 59044 146248 59050 146260
rect 59354 146248 59360 146260
rect 59044 146220 59360 146248
rect 59044 146208 59050 146220
rect 59354 146208 59360 146220
rect 59412 146248 59418 146260
rect 92474 146248 92480 146260
rect 59412 146220 92480 146248
rect 59412 146208 59418 146220
rect 92474 146208 92480 146220
rect 92532 146208 92538 146260
rect 179046 146208 179052 146260
rect 179104 146248 179110 146260
rect 197538 146248 197544 146260
rect 179104 146220 197544 146248
rect 179104 146208 179110 146220
rect 197538 146208 197544 146220
rect 197596 146208 197602 146260
rect 219710 146208 219716 146260
rect 219768 146248 219774 146260
rect 253934 146248 253940 146260
rect 219768 146220 253940 146248
rect 219768 146208 219774 146220
rect 253934 146208 253940 146220
rect 253992 146208 253998 146260
rect 277366 146248 277394 146276
rect 357434 146248 357440 146260
rect 277366 146220 357440 146248
rect 357434 146208 357440 146220
rect 357492 146208 357498 146260
rect 358722 146208 358728 146260
rect 358780 146248 358786 146260
rect 510614 146248 510620 146260
rect 358780 146220 510620 146248
rect 358780 146208 358786 146220
rect 510614 146208 510620 146220
rect 510672 146208 510678 146260
rect 54202 146140 54208 146192
rect 54260 146180 54266 146192
rect 56318 146180 56324 146192
rect 54260 146152 56324 146180
rect 54260 146140 54266 146152
rect 56318 146140 56324 146152
rect 56376 146140 56382 146192
rect 58710 146140 58716 146192
rect 58768 146180 58774 146192
rect 59630 146180 59636 146192
rect 58768 146152 59636 146180
rect 58768 146140 58774 146152
rect 59630 146140 59636 146152
rect 59688 146140 59694 146192
rect 85574 146180 85580 146192
rect 59740 146152 85580 146180
rect 53282 146004 53288 146056
rect 53340 146044 53346 146056
rect 59740 146044 59768 146152
rect 85574 146140 85580 146152
rect 85632 146140 85638 146192
rect 179690 146140 179696 146192
rect 179748 146180 179754 146192
rect 197446 146180 197452 146192
rect 179748 146152 197452 146180
rect 179748 146140 179754 146152
rect 197446 146140 197452 146152
rect 197504 146140 197510 146192
rect 219802 146140 219808 146192
rect 219860 146180 219866 146192
rect 219860 146152 229094 146180
rect 219860 146140 219866 146152
rect 60918 146072 60924 146124
rect 60976 146112 60982 146124
rect 86954 146112 86960 146124
rect 60976 146084 86960 146112
rect 60976 146072 60982 146084
rect 86954 146072 86960 146084
rect 87012 146072 87018 146124
rect 229066 146112 229094 146152
rect 235258 146140 235264 146192
rect 235316 146180 235322 146192
rect 255406 146180 255412 146192
rect 235316 146152 255412 146180
rect 235316 146140 235322 146152
rect 255406 146140 255412 146152
rect 255464 146140 255470 146192
rect 338482 146140 338488 146192
rect 338540 146180 338546 146192
rect 357710 146180 357716 146192
rect 338540 146152 357716 146180
rect 338540 146140 338546 146152
rect 357710 146140 357716 146152
rect 357768 146140 357774 146192
rect 374454 146140 374460 146192
rect 374512 146180 374518 146192
rect 375742 146180 375748 146192
rect 374512 146152 375748 146180
rect 374512 146140 374518 146152
rect 375742 146140 375748 146152
rect 375800 146140 375806 146192
rect 375926 146140 375932 146192
rect 375984 146180 375990 146192
rect 376294 146180 376300 146192
rect 375984 146152 376300 146180
rect 375984 146140 375990 146152
rect 376294 146140 376300 146152
rect 376352 146140 376358 146192
rect 378870 146140 378876 146192
rect 378928 146180 378934 146192
rect 379238 146180 379244 146192
rect 378928 146152 379244 146180
rect 378928 146140 378934 146152
rect 379238 146140 379244 146152
rect 379296 146140 379302 146192
rect 396718 146140 396724 146192
rect 396776 146180 396782 146192
rect 418154 146180 418160 146192
rect 396776 146152 418160 146180
rect 396776 146140 396782 146152
rect 418154 146140 418160 146152
rect 418212 146140 418218 146192
rect 498654 146140 498660 146192
rect 498712 146180 498718 146192
rect 517606 146180 517612 146192
rect 498712 146152 517612 146180
rect 498712 146140 498718 146152
rect 517606 146140 517612 146152
rect 517664 146180 517670 146192
rect 518434 146180 518440 146192
rect 517664 146152 518440 146180
rect 517664 146140 517670 146152
rect 518434 146140 518440 146152
rect 518492 146140 518498 146192
rect 252554 146112 252560 146124
rect 229066 146084 252560 146112
rect 252554 146072 252560 146084
rect 252612 146072 252618 146124
rect 340230 146072 340236 146124
rect 340288 146112 340294 146124
rect 357618 146112 357624 146124
rect 340288 146084 357624 146112
rect 340288 146072 340294 146084
rect 357618 146072 357624 146084
rect 357676 146072 357682 146124
rect 379974 146072 379980 146124
rect 380032 146112 380038 146124
rect 414014 146112 414020 146124
rect 380032 146084 414020 146112
rect 380032 146072 380038 146084
rect 414014 146072 414020 146084
rect 414072 146072 414078 146124
rect 499850 146072 499856 146124
rect 499908 146112 499914 146124
rect 517514 146112 517520 146124
rect 499908 146084 517520 146112
rect 499908 146072 499914 146084
rect 517514 146072 517520 146084
rect 517572 146112 517578 146124
rect 517698 146112 517704 146124
rect 517572 146084 517704 146112
rect 517572 146072 517578 146084
rect 517698 146072 517704 146084
rect 517756 146072 517762 146124
rect 53340 146016 59768 146044
rect 53340 146004 53346 146016
rect 60090 146004 60096 146056
rect 60148 146044 60154 146056
rect 89806 146044 89812 146056
rect 60148 146016 89812 146044
rect 60148 146004 60154 146016
rect 89806 146004 89812 146016
rect 89864 146004 89870 146056
rect 216490 146004 216496 146056
rect 216548 146044 216554 146056
rect 248414 146044 248420 146056
rect 216548 146016 248420 146044
rect 216548 146004 216554 146016
rect 248414 146004 248420 146016
rect 248472 146004 248478 146056
rect 375926 146004 375932 146056
rect 375984 146044 375990 146056
rect 377950 146044 377956 146056
rect 375984 146016 377956 146044
rect 375984 146004 375990 146016
rect 377950 146004 377956 146016
rect 378008 146004 378014 146056
rect 378962 146004 378968 146056
rect 379020 146044 379026 146056
rect 411254 146044 411260 146056
rect 379020 146016 411260 146044
rect 379020 146004 379026 146016
rect 411254 146004 411260 146016
rect 411312 146004 411318 146056
rect 54110 145936 54116 145988
rect 54168 145976 54174 145988
rect 54754 145976 54760 145988
rect 54168 145948 54760 145976
rect 54168 145936 54174 145948
rect 54754 145936 54760 145948
rect 54812 145976 54818 145988
rect 84286 145976 84292 145988
rect 54812 145948 84292 145976
rect 54812 145936 54818 145948
rect 84286 145936 84292 145948
rect 84344 145936 84350 145988
rect 220078 145936 220084 145988
rect 220136 145976 220142 145988
rect 251174 145976 251180 145988
rect 220136 145948 251180 145976
rect 220136 145936 220142 145948
rect 251174 145936 251180 145948
rect 251232 145936 251238 145988
rect 376294 145936 376300 145988
rect 376352 145976 376358 145988
rect 407114 145976 407120 145988
rect 376352 145948 407120 145976
rect 376352 145936 376358 145948
rect 407114 145936 407120 145948
rect 407172 145936 407178 145988
rect 54294 145868 54300 145920
rect 54352 145908 54358 145920
rect 54478 145908 54484 145920
rect 54352 145880 54484 145908
rect 54352 145868 54358 145880
rect 54478 145868 54484 145880
rect 54536 145908 54542 145920
rect 82814 145908 82820 145920
rect 54536 145880 82820 145908
rect 54536 145868 54542 145880
rect 82814 145868 82820 145880
rect 82872 145868 82878 145920
rect 219894 145868 219900 145920
rect 219952 145908 219958 145920
rect 251266 145908 251272 145920
rect 219952 145880 251272 145908
rect 219952 145868 219958 145880
rect 251266 145868 251272 145880
rect 251324 145868 251330 145920
rect 377306 145868 377312 145920
rect 377364 145908 377370 145920
rect 379054 145908 379060 145920
rect 377364 145880 379060 145908
rect 377364 145868 377370 145880
rect 379054 145868 379060 145880
rect 379112 145908 379118 145920
rect 409966 145908 409972 145920
rect 379112 145880 409972 145908
rect 379112 145868 379118 145880
rect 409966 145868 409972 145880
rect 410024 145868 410030 145920
rect 56410 145800 56416 145852
rect 56468 145840 56474 145852
rect 84194 145840 84200 145852
rect 56468 145812 84200 145840
rect 56468 145800 56474 145812
rect 84194 145800 84200 145812
rect 84252 145800 84258 145852
rect 214374 145800 214380 145852
rect 214432 145840 214438 145852
rect 215202 145840 215208 145852
rect 214432 145812 215208 145840
rect 214432 145800 214438 145812
rect 215202 145800 215208 145812
rect 215260 145800 215266 145852
rect 219158 145800 219164 145852
rect 219216 145840 219222 145852
rect 249886 145840 249892 145852
rect 219216 145812 249892 145840
rect 219216 145800 219222 145812
rect 249886 145800 249892 145812
rect 249944 145800 249950 145852
rect 377950 145800 377956 145852
rect 378008 145840 378014 145852
rect 408494 145840 408500 145852
rect 378008 145812 408500 145840
rect 378008 145800 378014 145812
rect 408494 145800 408500 145812
rect 408552 145800 408558 145852
rect 56318 145732 56324 145784
rect 56376 145772 56382 145784
rect 88426 145772 88432 145784
rect 56376 145744 88432 145772
rect 56376 145732 56382 145744
rect 88426 145732 88432 145744
rect 88484 145732 88490 145784
rect 217226 145732 217232 145784
rect 217284 145772 217290 145784
rect 245654 145772 245660 145784
rect 217284 145744 245660 145772
rect 217284 145732 217290 145744
rect 245654 145732 245660 145744
rect 245712 145732 245718 145784
rect 375742 145732 375748 145784
rect 375800 145772 375806 145784
rect 402974 145772 402980 145784
rect 375800 145744 402980 145772
rect 375800 145732 375806 145744
rect 402974 145732 402980 145744
rect 403032 145732 403038 145784
rect 57514 145664 57520 145716
rect 57572 145704 57578 145716
rect 91186 145704 91192 145716
rect 57572 145676 91192 145704
rect 57572 145664 57578 145676
rect 91186 145664 91192 145676
rect 91244 145664 91250 145716
rect 216214 145664 216220 145716
rect 216272 145704 216278 145716
rect 242894 145704 242900 145716
rect 216272 145676 242900 145704
rect 216272 145664 216278 145676
rect 242894 145664 242900 145676
rect 242952 145664 242958 145716
rect 343542 145664 343548 145716
rect 343600 145704 343606 145716
rect 356606 145704 356612 145716
rect 343600 145676 356612 145704
rect 343600 145664 343606 145676
rect 356606 145664 356612 145676
rect 356664 145664 356670 145716
rect 378870 145664 378876 145716
rect 378928 145704 378934 145716
rect 403066 145704 403072 145716
rect 378928 145676 403072 145704
rect 378928 145664 378934 145676
rect 403066 145664 403072 145676
rect 403124 145664 403130 145716
rect 503622 145664 503628 145716
rect 503680 145704 503686 145716
rect 517790 145704 517796 145716
rect 503680 145676 517796 145704
rect 503680 145664 503686 145676
rect 517790 145664 517796 145676
rect 517848 145664 517854 145716
rect 59630 145596 59636 145648
rect 59688 145636 59694 145648
rect 93854 145636 93860 145648
rect 59688 145608 93860 145636
rect 59688 145596 59694 145608
rect 93854 145596 93860 145608
rect 93912 145596 93918 145648
rect 183462 145596 183468 145648
rect 183520 145636 183526 145648
rect 197446 145636 197452 145648
rect 183520 145608 197452 145636
rect 183520 145596 183526 145608
rect 197446 145596 197452 145608
rect 197504 145596 197510 145648
rect 218514 145596 218520 145648
rect 218572 145636 218578 145648
rect 244366 145636 244372 145648
rect 218572 145608 244372 145636
rect 218572 145596 218578 145608
rect 244366 145596 244372 145608
rect 244424 145596 244430 145648
rect 280062 145596 280068 145648
rect 280120 145636 280126 145648
rect 356698 145636 356704 145648
rect 280120 145608 356704 145636
rect 280120 145596 280126 145608
rect 356698 145596 356704 145608
rect 356756 145636 356762 145648
rect 358814 145636 358820 145648
rect 356756 145608 358820 145636
rect 356756 145596 356762 145608
rect 358814 145596 358820 145608
rect 358872 145596 358878 145648
rect 378778 145596 378784 145648
rect 378836 145636 378842 145648
rect 405734 145636 405740 145648
rect 378836 145608 405740 145636
rect 378836 145596 378842 145608
rect 405734 145596 405740 145608
rect 405792 145596 405798 145648
rect 517514 145596 517520 145648
rect 517572 145636 517578 145648
rect 580258 145636 580264 145648
rect 517572 145608 580264 145636
rect 517572 145596 517578 145608
rect 580258 145596 580264 145608
rect 580316 145596 580322 145648
rect 58618 145528 58624 145580
rect 58676 145568 58682 145580
rect 100754 145568 100760 145580
rect 58676 145540 100760 145568
rect 58676 145528 58682 145540
rect 100754 145528 100760 145540
rect 100812 145528 100818 145580
rect 191742 145528 191748 145580
rect 191800 145568 191806 145580
rect 197998 145568 198004 145580
rect 191800 145540 198004 145568
rect 191800 145528 191806 145540
rect 197998 145528 198004 145540
rect 198056 145568 198062 145580
rect 214558 145568 214564 145580
rect 198056 145540 214564 145568
rect 198056 145528 198062 145540
rect 214558 145528 214564 145540
rect 214616 145528 214622 145580
rect 216490 145528 216496 145580
rect 216548 145568 216554 145580
rect 244274 145568 244280 145580
rect 216548 145540 244280 145568
rect 216548 145528 216554 145540
rect 244274 145528 244280 145540
rect 244332 145528 244338 145580
rect 351638 145528 351644 145580
rect 351696 145568 351702 145580
rect 358722 145568 358728 145580
rect 351696 145540 358728 145568
rect 351696 145528 351702 145540
rect 358722 145528 358728 145540
rect 358780 145528 358786 145580
rect 376570 145528 376576 145580
rect 376628 145568 376634 145580
rect 404354 145568 404360 145580
rect 376628 145540 404360 145568
rect 376628 145528 376634 145540
rect 404354 145528 404360 145540
rect 404412 145528 404418 145580
rect 518434 145528 518440 145580
rect 518492 145568 518498 145580
rect 580350 145568 580356 145580
rect 518492 145540 580356 145568
rect 518492 145528 518498 145540
rect 580350 145528 580356 145540
rect 580408 145528 580414 145580
rect 51902 145460 51908 145512
rect 51960 145500 51966 145512
rect 77294 145500 77300 145512
rect 51960 145472 77300 145500
rect 51960 145460 51966 145472
rect 77294 145460 77300 145472
rect 77352 145460 77358 145512
rect 214282 145460 214288 145512
rect 214340 145500 214346 145512
rect 235994 145500 236000 145512
rect 214340 145472 236000 145500
rect 214340 145460 214346 145472
rect 235994 145460 236000 145472
rect 236052 145460 236058 145512
rect 371694 145460 371700 145512
rect 371752 145500 371758 145512
rect 373442 145500 373448 145512
rect 371752 145472 373448 145500
rect 371752 145460 371758 145472
rect 373442 145460 373448 145472
rect 373500 145500 373506 145512
rect 397454 145500 397460 145512
rect 373500 145472 397460 145500
rect 373500 145460 373506 145472
rect 397454 145460 397460 145472
rect 397512 145460 397518 145512
rect 48038 145392 48044 145444
rect 48096 145432 48102 145444
rect 54662 145432 54668 145444
rect 48096 145404 54668 145432
rect 48096 145392 48102 145404
rect 54662 145392 54668 145404
rect 54720 145432 54726 145444
rect 76006 145432 76012 145444
rect 54720 145404 76012 145432
rect 54720 145392 54726 145404
rect 76006 145392 76012 145404
rect 76064 145392 76070 145444
rect 215662 145392 215668 145444
rect 215720 145432 215726 145444
rect 236086 145432 236092 145444
rect 215720 145404 236092 145432
rect 215720 145392 215726 145404
rect 236086 145392 236092 145404
rect 236144 145392 236150 145444
rect 378594 145392 378600 145444
rect 378652 145432 378658 145444
rect 396166 145432 396172 145444
rect 378652 145404 396172 145432
rect 378652 145392 378658 145404
rect 396166 145392 396172 145404
rect 396224 145392 396230 145444
rect 46474 145324 46480 145376
rect 46532 145364 46538 145376
rect 54846 145364 54852 145376
rect 46532 145336 54852 145364
rect 46532 145324 46538 145336
rect 54846 145324 54852 145336
rect 54904 145364 54910 145376
rect 75914 145364 75920 145376
rect 54904 145336 75920 145364
rect 54904 145324 54910 145336
rect 75914 145324 75920 145336
rect 75972 145324 75978 145376
rect 215202 145324 215208 145376
rect 215260 145364 215266 145376
rect 247126 145364 247132 145376
rect 215260 145336 247132 145364
rect 215260 145324 215266 145336
rect 247126 145324 247132 145336
rect 247184 145324 247190 145376
rect 378686 145324 378692 145376
rect 378744 145364 378750 145376
rect 396074 145364 396080 145376
rect 378744 145336 396080 145364
rect 378744 145324 378750 145336
rect 396074 145324 396080 145336
rect 396132 145324 396138 145376
rect 56226 145256 56232 145308
rect 56284 145296 56290 145308
rect 60918 145296 60924 145308
rect 56284 145268 60924 145296
rect 56284 145256 56290 145268
rect 60918 145256 60924 145268
rect 60976 145256 60982 145308
rect 377030 145256 377036 145308
rect 377088 145296 377094 145308
rect 411346 145296 411352 145308
rect 377088 145268 411352 145296
rect 377088 145256 377094 145268
rect 411346 145256 411352 145268
rect 411404 145256 411410 145308
rect 217134 145052 217140 145104
rect 217192 145092 217198 145104
rect 220078 145092 220084 145104
rect 217192 145064 220084 145092
rect 217192 145052 217198 145064
rect 220078 145052 220084 145064
rect 220136 145052 220142 145104
rect 218606 144984 218612 145036
rect 218664 145024 218670 145036
rect 219802 145024 219808 145036
rect 218664 144996 219808 145024
rect 218664 144984 218670 144996
rect 219802 144984 219808 144996
rect 219860 144984 219866 145036
rect 218882 144916 218888 144968
rect 218940 144956 218946 144968
rect 219894 144956 219900 144968
rect 218940 144928 219900 144956
rect 218940 144916 218946 144928
rect 219894 144916 219900 144928
rect 219952 144916 219958 144968
rect 51718 144848 51724 144900
rect 51776 144888 51782 144900
rect 55950 144888 55956 144900
rect 51776 144860 55956 144888
rect 51776 144848 51782 144860
rect 55950 144848 55956 144860
rect 56008 144888 56014 144900
rect 56410 144888 56416 144900
rect 56008 144860 56416 144888
rect 56008 144848 56014 144860
rect 56410 144848 56416 144860
rect 56468 144848 56474 144900
rect 210786 144848 210792 144900
rect 210844 144888 210850 144900
rect 211798 144888 211804 144900
rect 210844 144860 211804 144888
rect 210844 144848 210850 144860
rect 211798 144848 211804 144860
rect 211856 144848 211862 144900
rect 213546 144848 213552 144900
rect 213604 144888 213610 144900
rect 218514 144888 218520 144900
rect 213604 144860 218520 144888
rect 213604 144848 213610 144860
rect 218514 144848 218520 144860
rect 218572 144848 218578 144900
rect 373626 144848 373632 144900
rect 373684 144888 373690 144900
rect 378778 144888 378784 144900
rect 373684 144860 378784 144888
rect 373684 144848 373690 144860
rect 378778 144848 378784 144860
rect 378836 144848 378842 144900
rect 50522 144780 50528 144832
rect 50580 144820 50586 144832
rect 55858 144820 55864 144832
rect 50580 144792 55864 144820
rect 50580 144780 50586 144792
rect 55858 144780 55864 144792
rect 55916 144820 55922 144832
rect 56502 144820 56508 144832
rect 55916 144792 56508 144820
rect 55916 144780 55922 144792
rect 56502 144780 56508 144792
rect 56560 144780 56566 144832
rect 212994 144780 213000 144832
rect 213052 144820 213058 144832
rect 215938 144820 215944 144832
rect 213052 144792 215944 144820
rect 213052 144780 213058 144792
rect 215938 144780 215944 144792
rect 215996 144820 216002 144832
rect 216398 144820 216404 144832
rect 215996 144792 216404 144820
rect 215996 144780 216002 144792
rect 216398 144780 216404 144792
rect 216456 144780 216462 144832
rect 373718 144780 373724 144832
rect 373776 144820 373782 144832
rect 376110 144820 376116 144832
rect 373776 144792 376116 144820
rect 373776 144780 373782 144792
rect 376110 144780 376116 144792
rect 376168 144820 376174 144832
rect 376570 144820 376576 144832
rect 376168 144792 376576 144820
rect 376168 144780 376174 144792
rect 376570 144780 376576 144792
rect 376628 144780 376634 144832
rect 51626 144712 51632 144764
rect 51684 144752 51690 144764
rect 58618 144752 58624 144764
rect 51684 144724 58624 144752
rect 51684 144712 51690 144724
rect 58618 144712 58624 144724
rect 58676 144712 58682 144764
rect 212258 144712 212264 144764
rect 212316 144752 212322 144764
rect 216030 144752 216036 144764
rect 212316 144724 216036 144752
rect 212316 144712 212322 144724
rect 216030 144712 216036 144724
rect 216088 144752 216094 144764
rect 216490 144752 216496 144764
rect 216088 144724 216496 144752
rect 216088 144712 216094 144724
rect 216490 144712 216496 144724
rect 216548 144712 216554 144764
rect 48130 144644 48136 144696
rect 48188 144684 48194 144696
rect 56962 144684 56968 144696
rect 48188 144656 56968 144684
rect 48188 144644 48194 144656
rect 56962 144644 56968 144656
rect 57020 144684 57026 144696
rect 57514 144684 57520 144696
rect 57020 144656 57520 144684
rect 57020 144644 57026 144656
rect 57514 144644 57520 144656
rect 57572 144644 57578 144696
rect 48222 144576 48228 144628
rect 48280 144616 48286 144628
rect 58710 144616 58716 144628
rect 48280 144588 58716 144616
rect 48280 144576 48286 144588
rect 58710 144576 58716 144588
rect 58768 144576 58774 144628
rect 215662 143692 215668 143744
rect 215720 143732 215726 143744
rect 216490 143732 216496 143744
rect 215720 143704 216496 143732
rect 215720 143692 215726 143704
rect 216490 143692 216496 143704
rect 216548 143692 216554 143744
rect 55674 96568 55680 96620
rect 55732 96608 55738 96620
rect 57054 96608 57060 96620
rect 55732 96580 57060 96608
rect 55732 96568 55738 96580
rect 57054 96568 57060 96580
rect 57112 96568 57118 96620
rect 215846 96568 215852 96620
rect 215904 96608 215910 96620
rect 217502 96608 217508 96620
rect 215904 96580 217508 96608
rect 215904 96568 215910 96580
rect 217502 96568 217508 96580
rect 217560 96568 217566 96620
rect 520182 79976 520188 80028
rect 520240 80016 520246 80028
rect 580442 80016 580448 80028
rect 520240 79988 580448 80016
rect 520240 79976 520246 79988
rect 580442 79976 580448 79988
rect 580500 79976 580506 80028
rect 41322 70320 41328 70372
rect 41380 70360 41386 70372
rect 57514 70360 57520 70372
rect 41380 70332 57520 70360
rect 41380 70320 41386 70332
rect 57514 70320 57520 70332
rect 57572 70320 57578 70372
rect 370498 70320 370504 70372
rect 370556 70360 370562 70372
rect 376938 70360 376944 70372
rect 370556 70332 376944 70360
rect 370556 70320 370562 70332
rect 376938 70320 376944 70332
rect 376996 70320 377002 70372
rect 214558 68960 214564 69012
rect 214616 69000 214622 69012
rect 215202 69000 215208 69012
rect 214616 68972 215208 69000
rect 214616 68960 214622 68972
rect 215202 68960 215208 68972
rect 215260 68960 215266 69012
rect 213270 68892 213276 68944
rect 213328 68932 213334 68944
rect 216766 68932 216772 68944
rect 213328 68904 216772 68932
rect 213328 68892 213334 68904
rect 216766 68892 216772 68904
rect 216824 68892 216830 68944
rect 215202 68348 215208 68400
rect 215260 68388 215266 68400
rect 216674 68388 216680 68400
rect 215260 68360 216680 68388
rect 215260 68348 215266 68360
rect 216674 68348 216680 68360
rect 216732 68348 216738 68400
rect 358722 68280 358728 68332
rect 358780 68320 358786 68332
rect 376938 68320 376944 68332
rect 358780 68292 376944 68320
rect 358780 68280 358786 68292
rect 376938 68280 376944 68292
rect 376996 68280 377002 68332
rect 358078 68144 358084 68196
rect 358136 68184 358142 68196
rect 358722 68184 358728 68196
rect 358136 68156 358728 68184
rect 358136 68144 358142 68156
rect 358722 68144 358728 68156
rect 358780 68144 358786 68196
rect 214742 61956 214748 62008
rect 214800 61996 214806 62008
rect 214926 61996 214932 62008
rect 214800 61968 214932 61996
rect 214800 61956 214806 61968
rect 214926 61956 214932 61968
rect 214984 61956 214990 62008
rect 378962 60664 378968 60716
rect 379020 60704 379026 60716
rect 379238 60704 379244 60716
rect 379020 60676 379244 60704
rect 379020 60664 379026 60676
rect 379238 60664 379244 60676
rect 379296 60664 379302 60716
rect 54662 59780 54668 59832
rect 54720 59820 54726 59832
rect 77110 59820 77116 59832
rect 54720 59792 77116 59820
rect 54720 59780 54726 59792
rect 77110 59780 77116 59792
rect 77168 59780 77174 59832
rect 55950 59712 55956 59764
rect 56008 59752 56014 59764
rect 84194 59752 84200 59764
rect 56008 59724 84200 59752
rect 56008 59712 56014 59724
rect 84194 59712 84200 59724
rect 84252 59712 84258 59764
rect 378686 59712 378692 59764
rect 378744 59752 378750 59764
rect 396074 59752 396080 59764
rect 378744 59724 396080 59752
rect 378744 59712 378750 59724
rect 396074 59712 396080 59724
rect 396132 59712 396138 59764
rect 55858 59644 55864 59696
rect 55916 59684 55922 59696
rect 100754 59684 100760 59696
rect 55916 59656 100760 59684
rect 55916 59644 55922 59656
rect 100754 59644 100760 59656
rect 100812 59644 100818 59696
rect 217962 59644 217968 59696
rect 218020 59684 218026 59696
rect 255866 59684 255872 59696
rect 218020 59656 255872 59684
rect 218020 59644 218026 59656
rect 255866 59644 255872 59656
rect 255924 59644 255930 59696
rect 378594 59644 378600 59696
rect 378652 59684 378658 59696
rect 397086 59684 397092 59696
rect 378652 59656 397092 59684
rect 378652 59644 378658 59656
rect 397086 59644 397092 59656
rect 397144 59644 397150 59696
rect 54478 59576 54484 59628
rect 54536 59616 54542 59628
rect 83090 59616 83096 59628
rect 54536 59588 83096 59616
rect 54536 59576 54542 59588
rect 83090 59576 83096 59588
rect 83148 59576 83154 59628
rect 219066 59576 219072 59628
rect 219124 59616 219130 59628
rect 263870 59616 263876 59628
rect 219124 59588 263876 59616
rect 219124 59576 219130 59588
rect 263870 59576 263876 59588
rect 263928 59576 263934 59628
rect 378870 59576 378876 59628
rect 378928 59616 378934 59628
rect 403066 59616 403072 59628
rect 378928 59588 403072 59616
rect 378928 59576 378934 59588
rect 403066 59576 403072 59588
rect 403124 59576 403130 59628
rect 54570 59508 54576 59560
rect 54628 59548 54634 59560
rect 99466 59548 99472 59560
rect 54628 59520 99472 59548
rect 54628 59508 54634 59520
rect 99466 59508 99472 59520
rect 99524 59508 99530 59560
rect 216122 59508 216128 59560
rect 216180 59548 216186 59560
rect 261754 59548 261760 59560
rect 216180 59520 261760 59548
rect 216180 59508 216186 59520
rect 261754 59508 261760 59520
rect 261812 59508 261818 59560
rect 378042 59508 378048 59560
rect 378100 59548 378106 59560
rect 415854 59548 415860 59560
rect 378100 59520 415860 59548
rect 378100 59508 378106 59520
rect 415854 59508 415860 59520
rect 415912 59508 415918 59560
rect 56042 59440 56048 59492
rect 56100 59480 56106 59492
rect 102778 59480 102784 59492
rect 56100 59452 102784 59480
rect 56100 59440 56106 59452
rect 102778 59440 102784 59452
rect 102836 59440 102842 59492
rect 214650 59440 214656 59492
rect 214708 59480 214714 59492
rect 260650 59480 260656 59492
rect 214708 59452 260656 59480
rect 214708 59440 214714 59452
rect 260650 59440 260656 59452
rect 260708 59440 260714 59492
rect 376662 59440 376668 59492
rect 376720 59480 376726 59492
rect 419442 59480 419448 59492
rect 376720 59452 419448 59480
rect 376720 59440 376726 59452
rect 419442 59440 419448 59452
rect 419500 59440 419506 59492
rect 58802 59372 58808 59424
rect 58860 59412 58866 59424
rect 107562 59412 107568 59424
rect 58860 59384 107568 59412
rect 58860 59372 58866 59384
rect 107562 59372 107568 59384
rect 107620 59372 107626 59424
rect 215754 59372 215760 59424
rect 215812 59412 215818 59424
rect 262858 59412 262864 59424
rect 215812 59384 262864 59412
rect 215812 59372 215818 59384
rect 262858 59372 262864 59384
rect 262916 59372 262922 59424
rect 360930 59372 360936 59424
rect 360988 59412 360994 59424
rect 413554 59412 413560 59424
rect 360988 59384 413560 59412
rect 360988 59372 360994 59384
rect 413554 59372 413560 59384
rect 413612 59372 413618 59424
rect 54754 59304 54760 59356
rect 54812 59344 54818 59356
rect 85390 59344 85396 59356
rect 54812 59316 85396 59344
rect 54812 59304 54818 59316
rect 85390 59304 85396 59316
rect 85448 59304 85454 59356
rect 214742 59304 214748 59356
rect 214800 59344 214806 59356
rect 215202 59344 215208 59356
rect 214800 59316 215208 59344
rect 214800 59304 214806 59316
rect 215202 59304 215208 59316
rect 215260 59344 215266 59356
rect 358078 59344 358084 59356
rect 215260 59316 358084 59344
rect 215260 59304 215266 59316
rect 358078 59304 358084 59316
rect 358136 59304 358142 59356
rect 373442 59304 373448 59356
rect 373500 59344 373506 59356
rect 398190 59344 398196 59356
rect 373500 59316 398196 59344
rect 373500 59304 373506 59316
rect 398190 59304 398196 59316
rect 398248 59304 398254 59356
rect 59078 59236 59084 59288
rect 59136 59276 59142 59288
rect 95878 59276 95884 59288
rect 59136 59248 95884 59276
rect 59136 59236 59142 59248
rect 95878 59236 95884 59248
rect 95936 59236 95942 59288
rect 374638 59236 374644 59288
rect 374696 59276 374702 59288
rect 410702 59276 410708 59288
rect 374696 59248 410708 59276
rect 374696 59236 374702 59248
rect 410702 59236 410708 59248
rect 410760 59236 410766 59288
rect 55030 59168 55036 59220
rect 55088 59208 55094 59220
rect 98086 59208 98092 59220
rect 55088 59180 98092 59208
rect 55088 59168 55094 59180
rect 98086 59168 98092 59180
rect 98144 59168 98150 59220
rect 219434 59168 219440 59220
rect 219492 59208 219498 59220
rect 256970 59208 256976 59220
rect 219492 59180 256976 59208
rect 219492 59168 219498 59180
rect 256970 59168 256976 59180
rect 257028 59168 257034 59220
rect 379146 59168 379152 59220
rect 379204 59208 379210 59220
rect 416958 59208 416964 59220
rect 379204 59180 416964 59208
rect 379204 59168 379210 59180
rect 416958 59168 416964 59180
rect 417016 59168 417022 59220
rect 59814 59100 59820 59152
rect 59872 59140 59878 59152
rect 106366 59140 106372 59152
rect 59872 59112 106372 59140
rect 59872 59100 59878 59112
rect 106366 59100 106372 59112
rect 106424 59100 106430 59152
rect 214926 59100 214932 59152
rect 214984 59140 214990 59152
rect 259454 59140 259460 59152
rect 214984 59112 259460 59140
rect 214984 59100 214990 59112
rect 259454 59100 259460 59112
rect 259512 59100 259518 59152
rect 379606 59100 379612 59152
rect 379664 59140 379670 59152
rect 418154 59140 418160 59152
rect 379664 59112 418160 59140
rect 379664 59100 379670 59112
rect 418154 59100 418160 59112
rect 418212 59100 418218 59152
rect 56134 59032 56140 59084
rect 56192 59072 56198 59084
rect 103882 59072 103888 59084
rect 56192 59044 103888 59072
rect 56192 59032 56198 59044
rect 103882 59032 103888 59044
rect 103940 59032 103946 59084
rect 213822 59032 213828 59084
rect 213880 59072 213886 59084
rect 298462 59072 298468 59084
rect 213880 59044 298468 59072
rect 213880 59032 213886 59044
rect 298462 59032 298468 59044
rect 298520 59032 298526 59084
rect 379698 59032 379704 59084
rect 379756 59072 379762 59084
rect 425238 59072 425244 59084
rect 379756 59044 425244 59072
rect 379756 59032 379762 59044
rect 425238 59032 425244 59044
rect 425296 59032 425302 59084
rect 57330 58964 57336 59016
rect 57388 59004 57394 59016
rect 105262 59004 105268 59016
rect 57388 58976 105268 59004
rect 57388 58964 57394 58976
rect 105262 58964 105268 58976
rect 105320 58964 105326 59016
rect 198550 58964 198556 59016
rect 198608 59004 198614 59016
rect 295886 59004 295892 59016
rect 198608 58976 295892 59004
rect 198608 58964 198614 58976
rect 295886 58964 295892 58976
rect 295944 58964 295950 59016
rect 374362 58964 374368 59016
rect 374420 59004 374426 59016
rect 421742 59004 421748 59016
rect 374420 58976 421748 59004
rect 374420 58964 374426 58976
rect 421742 58964 421748 58976
rect 421800 58964 421806 59016
rect 53190 58896 53196 58948
rect 53248 58936 53254 58948
rect 114370 58936 114376 58948
rect 53248 58908 114376 58936
rect 53248 58896 53254 58908
rect 114370 58896 114376 58908
rect 114428 58896 114434 58948
rect 209038 58896 209044 58948
rect 209096 58936 209102 58948
rect 308490 58936 308496 58948
rect 209096 58908 308496 58936
rect 209096 58896 209102 58908
rect 308490 58896 308496 58908
rect 308548 58896 308554 58948
rect 358170 58896 358176 58948
rect 358228 58936 358234 58948
rect 423490 58936 423496 58948
rect 358228 58908 423496 58936
rect 358228 58896 358234 58908
rect 423490 58896 423496 58908
rect 423548 58896 423554 58948
rect 55582 58828 55588 58880
rect 55640 58868 55646 58880
rect 138382 58868 138388 58880
rect 55640 58840 138388 58868
rect 55640 58828 55646 58840
rect 138382 58828 138388 58840
rect 138440 58828 138446 58880
rect 201402 58828 201408 58880
rect 201460 58868 201466 58880
rect 303430 58868 303436 58880
rect 201460 58840 303436 58868
rect 201460 58828 201466 58840
rect 303430 58828 303436 58840
rect 303488 58828 303494 58880
rect 363690 58828 363696 58880
rect 363748 58868 363754 58880
rect 468478 58868 468484 58880
rect 363748 58840 468484 58868
rect 363748 58828 363754 58840
rect 468478 58828 468484 58840
rect 468536 58828 468542 58880
rect 52178 58760 52184 58812
rect 52236 58800 52242 58812
rect 143534 58800 143540 58812
rect 52236 58772 143540 58800
rect 52236 58760 52242 58772
rect 143534 58760 143540 58772
rect 143592 58760 143598 58812
rect 219342 58760 219348 58812
rect 219400 58800 219406 58812
rect 425974 58800 425980 58812
rect 219400 58772 425980 58800
rect 219400 58760 219406 58772
rect 425974 58760 425980 58772
rect 426032 58760 426038 58812
rect 55490 58692 55496 58744
rect 55548 58732 55554 58744
rect 150894 58732 150900 58744
rect 55548 58704 150900 58732
rect 55548 58692 55554 58704
rect 150894 58692 150900 58704
rect 150952 58692 150958 58744
rect 219618 58692 219624 58744
rect 219676 58732 219682 58744
rect 421006 58732 421012 58744
rect 219676 58704 421012 58732
rect 219676 58692 219682 58704
rect 421006 58692 421012 58704
rect 421064 58692 421070 58744
rect 50062 58624 50068 58676
rect 50120 58664 50126 58676
rect 148502 58664 148508 58676
rect 50120 58636 148508 58664
rect 50120 58624 50126 58636
rect 148502 58624 148508 58636
rect 148560 58624 148566 58676
rect 219066 58624 219072 58676
rect 219124 58664 219130 58676
rect 428182 58664 428188 58676
rect 219124 58636 428188 58664
rect 219124 58624 219130 58636
rect 428182 58624 428188 58636
rect 428240 58624 428246 58676
rect 219342 57944 219348 57996
rect 219400 57984 219406 57996
rect 430942 57984 430948 57996
rect 219400 57956 430948 57984
rect 219400 57944 219406 57956
rect 430942 57944 430948 57956
rect 431000 57944 431006 57996
rect 57238 57876 57244 57928
rect 57296 57916 57302 57928
rect 57882 57916 57888 57928
rect 57296 57888 57888 57916
rect 57296 57876 57302 57888
rect 57882 57876 57888 57888
rect 57940 57916 57946 57928
rect 214742 57916 214748 57928
rect 57940 57888 214748 57916
rect 57940 57876 57946 57888
rect 214742 57876 214748 57888
rect 214800 57876 214806 57928
rect 343174 57876 343180 57928
rect 343232 57916 343238 57928
rect 357526 57916 357532 57928
rect 343232 57888 357532 57916
rect 343232 57876 343238 57888
rect 357526 57876 357532 57888
rect 357584 57876 357590 57928
rect 361482 57876 361488 57928
rect 361540 57916 361546 57928
rect 475838 57916 475844 57928
rect 361540 57888 475844 57916
rect 361540 57876 361546 57888
rect 475838 57876 475844 57888
rect 475896 57876 475902 57928
rect 503346 57876 503352 57928
rect 503404 57916 503410 57928
rect 517790 57916 517796 57928
rect 503404 57888 517796 57916
rect 503404 57876 503410 57888
rect 517790 57876 517796 57888
rect 517848 57876 517854 57928
rect 53742 57808 53748 57860
rect 53800 57848 53806 57860
rect 145558 57848 145564 57860
rect 53800 57820 145564 57848
rect 53800 57808 53806 57820
rect 145558 57808 145564 57820
rect 145616 57808 145622 57860
rect 183462 57808 183468 57860
rect 183520 57848 183526 57860
rect 197446 57848 197452 57860
rect 183520 57820 197452 57848
rect 183520 57808 183526 57820
rect 197446 57808 197452 57820
rect 197504 57808 197510 57860
rect 209682 57808 209688 57860
rect 209740 57848 209746 57860
rect 325878 57848 325884 57860
rect 209740 57820 325884 57848
rect 209740 57808 209746 57820
rect 325878 57808 325884 57820
rect 325936 57808 325942 57860
rect 343450 57808 343456 57860
rect 343508 57848 343514 57860
rect 356606 57848 356612 57860
rect 343508 57820 356612 57848
rect 343508 57808 343514 57820
rect 356606 57808 356612 57820
rect 356664 57808 356670 57860
rect 373902 57808 373908 57860
rect 373960 57848 373966 57860
rect 480622 57848 480628 57860
rect 373960 57820 480628 57848
rect 373960 57808 373966 57820
rect 480622 57808 480628 57820
rect 480680 57808 480686 57860
rect 503254 57808 503260 57860
rect 503312 57848 503318 57860
rect 517882 57848 517888 57860
rect 503312 57820 517888 57848
rect 503312 57808 503318 57820
rect 517882 57808 517888 57820
rect 517940 57808 517946 57860
rect 53650 57740 53656 57792
rect 53708 57780 53714 57792
rect 130838 57780 130844 57792
rect 53708 57752 130844 57780
rect 53708 57740 53714 57752
rect 130838 57740 130844 57752
rect 130896 57740 130902 57792
rect 183186 57740 183192 57792
rect 183244 57780 183250 57792
rect 197354 57780 197360 57792
rect 183244 57752 197360 57780
rect 183244 57740 183250 57752
rect 197354 57740 197360 57752
rect 197412 57740 197418 57792
rect 215018 57740 215024 57792
rect 215076 57780 215082 57792
rect 313366 57780 313372 57792
rect 215076 57752 313372 57780
rect 215076 57740 215082 57752
rect 313366 57740 313372 57752
rect 313424 57740 313430 57792
rect 378962 57740 378968 57792
rect 379020 57780 379026 57792
rect 483382 57780 483388 57792
rect 379020 57752 483388 57780
rect 379020 57740 379026 57752
rect 483382 57740 483388 57752
rect 483440 57740 483446 57792
rect 49602 57672 49608 57724
rect 49660 57712 49666 57724
rect 120718 57712 120724 57724
rect 49660 57684 120724 57712
rect 49660 57672 49666 57684
rect 120718 57672 120724 57684
rect 120776 57672 120782 57724
rect 212442 57672 212448 57724
rect 212500 57712 212506 57724
rect 310974 57712 310980 57724
rect 212500 57684 310980 57712
rect 212500 57672 212506 57684
rect 310974 57672 310980 57684
rect 311032 57672 311038 57724
rect 364978 57672 364984 57724
rect 365036 57712 365042 57724
rect 465902 57712 465908 57724
rect 365036 57684 465908 57712
rect 365036 57672 365042 57684
rect 465902 57672 465908 57684
rect 465960 57672 465966 57724
rect 49510 57604 49516 57656
rect 49568 57644 49574 57656
rect 113542 57644 113548 57656
rect 49568 57616 113548 57644
rect 49568 57604 49574 57616
rect 113542 57604 113548 57616
rect 113600 57604 113606 57656
rect 218974 57604 218980 57656
rect 219032 57644 219038 57656
rect 305822 57644 305828 57656
rect 219032 57616 305828 57644
rect 219032 57604 219038 57616
rect 305822 57604 305828 57616
rect 305880 57604 305886 57656
rect 366450 57604 366456 57656
rect 366508 57644 366514 57656
rect 460934 57644 460940 57656
rect 366508 57616 460940 57644
rect 366508 57604 366514 57616
rect 460934 57604 460940 57616
rect 460992 57604 460998 57656
rect 57054 57536 57060 57588
rect 57112 57576 57118 57588
rect 117958 57576 117964 57588
rect 57112 57548 117964 57576
rect 57112 57536 57118 57548
rect 117958 57536 117964 57548
rect 118016 57536 118022 57588
rect 216582 57536 216588 57588
rect 216640 57576 216646 57588
rect 300854 57576 300860 57588
rect 216640 57548 300860 57576
rect 216640 57536 216646 57548
rect 300854 57536 300860 57548
rect 300912 57536 300918 57588
rect 379422 57536 379428 57588
rect 379480 57576 379486 57588
rect 470870 57576 470876 57588
rect 379480 57548 470876 57576
rect 379480 57536 379486 57548
rect 470870 57536 470876 57548
rect 470928 57536 470934 57588
rect 59906 57468 59912 57520
rect 59964 57508 59970 57520
rect 108574 57508 108580 57520
rect 59964 57480 108580 57508
rect 59964 57468 59970 57480
rect 108574 57468 108580 57480
rect 108632 57468 108638 57520
rect 211062 57468 211068 57520
rect 211120 57508 211126 57520
rect 293310 57508 293316 57520
rect 211120 57480 293316 57508
rect 211120 57468 211126 57480
rect 293310 57468 293316 57480
rect 293368 57468 293374 57520
rect 362218 57468 362224 57520
rect 362276 57508 362282 57520
rect 433518 57508 433524 57520
rect 362276 57480 433524 57508
rect 362276 57468 362282 57480
rect 433518 57468 433524 57480
rect 433576 57468 433582 57520
rect 59998 57400 60004 57452
rect 60056 57440 60062 57452
rect 98454 57440 98460 57452
rect 60056 57412 98460 57440
rect 60056 57400 60062 57412
rect 98454 57400 98460 57412
rect 98512 57400 98518 57452
rect 213178 57400 213184 57452
rect 213236 57440 213242 57452
rect 268194 57440 268200 57452
rect 213236 57412 268200 57440
rect 213236 57400 213242 57412
rect 268194 57400 268200 57412
rect 268252 57400 268258 57452
rect 279050 57400 279056 57452
rect 279108 57440 279114 57452
rect 356698 57440 356704 57452
rect 279108 57412 356704 57440
rect 279108 57400 279114 57412
rect 356698 57400 356704 57412
rect 356756 57400 356762 57452
rect 367738 57400 367744 57452
rect 367796 57440 367802 57452
rect 438486 57440 438492 57452
rect 367796 57412 438492 57440
rect 367796 57400 367802 57412
rect 438486 57400 438492 57412
rect 438544 57400 438550 57452
rect 51534 57332 51540 57384
rect 51592 57372 51598 57384
rect 88426 57372 88432 57384
rect 51592 57344 88432 57372
rect 51592 57332 51598 57344
rect 88426 57332 88432 57344
rect 88484 57332 88490 57384
rect 215110 57332 215116 57384
rect 215168 57372 215174 57384
rect 287606 57372 287612 57384
rect 215168 57344 287612 57372
rect 215168 57332 215174 57344
rect 287606 57332 287612 57344
rect 287664 57332 287670 57384
rect 374730 57332 374736 57384
rect 374788 57372 374794 57384
rect 435910 57372 435916 57384
rect 374788 57344 435916 57372
rect 374788 57332 374794 57344
rect 435910 57332 435916 57344
rect 435968 57332 435974 57384
rect 59170 57264 59176 57316
rect 59228 57304 59234 57316
rect 93670 57304 93676 57316
rect 59228 57276 93676 57304
rect 59228 57264 59234 57276
rect 93670 57264 93676 57276
rect 93728 57264 93734 57316
rect 218790 57264 218796 57316
rect 218848 57304 218854 57316
rect 263594 57304 263600 57316
rect 218848 57276 263600 57304
rect 218848 57264 218854 57276
rect 263594 57264 263600 57276
rect 263652 57264 263658 57316
rect 373258 57264 373264 57316
rect 373316 57304 373322 57316
rect 418430 57304 418436 57316
rect 373316 57276 418436 57304
rect 373316 57264 373322 57276
rect 418430 57264 418436 57276
rect 418488 57264 418494 57316
rect 59262 57196 59268 57248
rect 59320 57236 59326 57248
rect 90726 57236 90732 57248
rect 59320 57208 90732 57236
rect 59320 57196 59326 57208
rect 90726 57196 90732 57208
rect 90784 57196 90790 57248
rect 218698 57196 218704 57248
rect 218756 57236 218762 57248
rect 248138 57236 248144 57248
rect 218756 57208 248144 57236
rect 218756 57196 218762 57208
rect 248138 57196 248144 57208
rect 248196 57196 248202 57248
rect 365070 57196 365076 57248
rect 365128 57236 365134 57248
rect 408310 57236 408316 57248
rect 365128 57208 408316 57236
rect 365128 57196 365134 57208
rect 408310 57196 408316 57208
rect 408368 57196 408374 57248
rect 54846 57128 54852 57180
rect 54904 57168 54910 57180
rect 76006 57168 76012 57180
rect 54904 57140 76012 57168
rect 54904 57128 54910 57140
rect 76006 57128 76012 57140
rect 76064 57128 76070 57180
rect 214098 57128 214104 57180
rect 214156 57168 214162 57180
rect 318242 57168 318248 57180
rect 214156 57140 318248 57168
rect 214156 57128 214162 57140
rect 318242 57128 318248 57140
rect 318300 57128 318306 57180
rect 41230 56516 41236 56568
rect 41288 56556 41294 56568
rect 123478 56556 123484 56568
rect 41288 56528 123484 56556
rect 41288 56516 41294 56528
rect 123478 56516 123484 56528
rect 123536 56516 123542 56568
rect 213086 56516 213092 56568
rect 213144 56556 213150 56568
rect 275646 56556 275652 56568
rect 213144 56528 275652 56556
rect 213144 56516 213150 56528
rect 275646 56516 275652 56528
rect 275704 56516 275710 56568
rect 375006 56516 375012 56568
rect 375064 56556 375070 56568
rect 435082 56556 435088 56568
rect 375064 56528 435088 56556
rect 375064 56516 375070 56528
rect 435082 56516 435088 56528
rect 435140 56516 435146 56568
rect 52270 56448 52276 56500
rect 52328 56488 52334 56500
rect 111150 56488 111156 56500
rect 52328 56460 111156 56488
rect 52328 56448 52334 56460
rect 111150 56448 111156 56460
rect 111208 56448 111214 56500
rect 217502 56448 217508 56500
rect 217560 56488 217566 56500
rect 278038 56488 278044 56500
rect 217560 56460 278044 56488
rect 217560 56448 217566 56460
rect 278038 56448 278044 56460
rect 278096 56448 278102 56500
rect 374546 56448 374552 56500
rect 374604 56488 374610 56500
rect 433334 56488 433340 56500
rect 374604 56460 433340 56488
rect 374604 56448 374610 56460
rect 433334 56448 433340 56460
rect 433392 56448 433398 56500
rect 53006 56380 53012 56432
rect 53064 56420 53070 56432
rect 109494 56420 109500 56432
rect 53064 56392 109500 56420
rect 53064 56380 53070 56392
rect 109494 56380 109500 56392
rect 109552 56380 109558 56432
rect 213730 56380 213736 56432
rect 213788 56420 213794 56432
rect 273254 56420 273260 56432
rect 213788 56392 273260 56420
rect 213788 56380 213794 56392
rect 273254 56380 273260 56392
rect 273312 56380 273318 56432
rect 374270 56380 374276 56432
rect 374328 56420 374334 56432
rect 430574 56420 430580 56432
rect 374328 56392 430580 56420
rect 374328 56380 374334 56392
rect 430574 56380 430580 56392
rect 430632 56380 430638 56432
rect 58618 56312 58624 56364
rect 58676 56352 58682 56364
rect 101766 56352 101772 56364
rect 58676 56324 101772 56352
rect 58676 56312 58682 56324
rect 101766 56312 101772 56324
rect 101824 56312 101830 56364
rect 215938 56312 215944 56364
rect 215996 56352 216002 56364
rect 271230 56352 271236 56364
rect 215996 56324 271236 56352
rect 215996 56312 216002 56324
rect 271230 56312 271236 56324
rect 271288 56312 271294 56364
rect 376386 56312 376392 56364
rect 376444 56352 376450 56364
rect 429654 56352 429660 56364
rect 376444 56324 429660 56352
rect 376444 56312 376450 56324
rect 429654 56312 429660 56324
rect 429712 56312 429718 56364
rect 59722 56244 59728 56296
rect 59780 56284 59786 56296
rect 94406 56284 94412 56296
rect 59780 56256 94412 56284
rect 59780 56244 59786 56256
rect 94406 56244 94412 56256
rect 94464 56244 94470 56296
rect 219986 56244 219992 56296
rect 220044 56284 220050 56296
rect 268654 56284 268660 56296
rect 220044 56256 268660 56284
rect 220044 56244 220050 56256
rect 268654 56244 268660 56256
rect 268712 56244 268718 56296
rect 379790 56244 379796 56296
rect 379848 56284 379854 56296
rect 427630 56284 427636 56296
rect 379848 56256 427636 56284
rect 379848 56244 379854 56256
rect 427630 56244 427636 56256
rect 427688 56244 427694 56296
rect 58710 56176 58716 56228
rect 58768 56216 58774 56228
rect 92198 56216 92204 56228
rect 58768 56188 92204 56216
rect 58768 56176 58774 56188
rect 92198 56176 92204 56188
rect 92256 56176 92262 56228
rect 219526 56176 219532 56228
rect 219584 56216 219590 56228
rect 266354 56216 266360 56228
rect 219584 56188 266360 56216
rect 219584 56176 219590 56188
rect 266354 56176 266360 56188
rect 266412 56176 266418 56228
rect 376202 56176 376208 56228
rect 376260 56216 376266 56228
rect 422846 56216 422852 56228
rect 376260 56188 422852 56216
rect 376260 56176 376266 56188
rect 422846 56176 422852 56188
rect 422904 56176 422910 56228
rect 53282 56108 53288 56160
rect 53340 56148 53346 56160
rect 86494 56148 86500 56160
rect 53340 56120 86500 56148
rect 53340 56108 53346 56120
rect 86494 56108 86500 56120
rect 86552 56108 86558 56160
rect 217134 56108 217140 56160
rect 217192 56148 217198 56160
rect 251174 56148 251180 56160
rect 217192 56120 251180 56148
rect 217192 56108 217198 56120
rect 251174 56108 251180 56120
rect 251232 56108 251238 56160
rect 379974 56108 379980 56160
rect 380032 56148 380038 56160
rect 414566 56148 414572 56160
rect 380032 56120 414572 56148
rect 380032 56108 380038 56120
rect 414566 56108 414572 56120
rect 414624 56108 414630 56160
rect 58894 56040 58900 56092
rect 58952 56080 58958 56092
rect 89990 56080 89996 56092
rect 58952 56052 89996 56080
rect 58952 56040 58958 56052
rect 89990 56040 89996 56052
rect 90048 56040 90054 56092
rect 218606 56040 218612 56092
rect 218664 56080 218670 56092
rect 253382 56080 253388 56092
rect 218664 56052 253388 56080
rect 218664 56040 218670 56052
rect 253382 56040 253388 56052
rect 253440 56040 253446 56092
rect 379330 56040 379336 56092
rect 379388 56080 379394 56092
rect 413462 56080 413468 56092
rect 379388 56052 413468 56080
rect 379388 56040 379394 56052
rect 413462 56040 413468 56052
rect 413520 56040 413526 56092
rect 51994 55972 52000 56024
rect 52052 56012 52058 56024
rect 80422 56012 80428 56024
rect 52052 55984 80428 56012
rect 52052 55972 52058 55984
rect 80422 55972 80428 55984
rect 80480 55972 80486 56024
rect 214374 55972 214380 56024
rect 214432 56012 214438 56024
rect 247678 56012 247684 56024
rect 214432 55984 247684 56012
rect 214432 55972 214438 55984
rect 247678 55972 247684 55984
rect 247736 55972 247742 56024
rect 375926 55972 375932 56024
rect 375984 56012 375990 56024
rect 408678 56012 408684 56024
rect 375984 55984 408684 56012
rect 375984 55972 375990 55984
rect 408678 55972 408684 55984
rect 408736 55972 408742 56024
rect 51902 55904 51908 55956
rect 51960 55944 51966 55956
rect 78214 55944 78220 55956
rect 51960 55916 78220 55944
rect 51960 55904 51966 55916
rect 78214 55904 78220 55916
rect 78272 55904 78278 55956
rect 216030 55904 216036 55956
rect 216088 55944 216094 55956
rect 245286 55944 245292 55956
rect 216088 55916 245292 55944
rect 216088 55904 216094 55916
rect 245286 55904 245292 55916
rect 245344 55904 245350 55956
rect 379238 55904 379244 55956
rect 379296 55944 379302 55956
rect 411254 55944 411260 55956
rect 379296 55916 411260 55944
rect 379296 55904 379302 55916
rect 411254 55904 411260 55916
rect 411312 55904 411318 55956
rect 211798 55836 211804 55888
rect 211856 55876 211862 55888
rect 238110 55876 238116 55888
rect 211856 55848 238116 55876
rect 211856 55836 211862 55848
rect 238110 55836 238116 55848
rect 238168 55836 238174 55888
rect 374454 55836 374460 55888
rect 374512 55876 374518 55888
rect 404078 55876 404084 55888
rect 374512 55848 404084 55876
rect 374512 55836 374518 55848
rect 404078 55836 404084 55848
rect 404136 55836 404142 55888
rect 213638 55768 213644 55820
rect 213696 55808 213702 55820
rect 240502 55808 240508 55820
rect 213696 55780 240508 55808
rect 213696 55768 213702 55780
rect 240502 55768 240508 55780
rect 240560 55768 240566 55820
rect 373350 55768 373356 55820
rect 373408 55808 373414 55820
rect 400398 55808 400404 55820
rect 373408 55780 400404 55808
rect 373408 55768 373414 55780
rect 400398 55768 400404 55780
rect 400456 55768 400462 55820
rect 54938 55156 54944 55208
rect 54996 55196 55002 55208
rect 114554 55196 114560 55208
rect 54996 55168 114560 55196
rect 54996 55156 55002 55168
rect 114554 55156 114560 55168
rect 114612 55156 114618 55208
rect 218514 55156 218520 55208
rect 218572 55196 218578 55208
rect 244366 55196 244372 55208
rect 218572 55168 244372 55196
rect 218572 55156 218578 55168
rect 244366 55156 244372 55168
rect 244424 55156 244430 55208
rect 375834 55156 375840 55208
rect 375892 55196 375898 55208
rect 436094 55196 436100 55208
rect 375892 55168 436100 55196
rect 375892 55156 375898 55168
rect 436094 55156 436100 55168
rect 436152 55156 436158 55208
rect 53558 55088 53564 55140
rect 53616 55128 53622 55140
rect 111794 55128 111800 55140
rect 53616 55100 111800 55128
rect 53616 55088 53622 55100
rect 111794 55088 111800 55100
rect 111852 55088 111858 55140
rect 214282 55088 214288 55140
rect 214340 55128 214346 55140
rect 235994 55128 236000 55140
rect 214340 55100 236000 55128
rect 214340 55088 214346 55100
rect 235994 55088 236000 55100
rect 236052 55088 236058 55140
rect 376478 55088 376484 55140
rect 376536 55128 376542 55140
rect 433702 55128 433708 55140
rect 376536 55100 433708 55128
rect 376536 55088 376542 55100
rect 433702 55088 433708 55100
rect 433760 55088 433766 55140
rect 54386 55020 54392 55072
rect 54444 55060 54450 55072
rect 113174 55060 113180 55072
rect 54444 55032 113180 55060
rect 54444 55020 54450 55032
rect 113174 55020 113180 55032
rect 113232 55020 113238 55072
rect 219250 55020 219256 55072
rect 219308 55060 219314 55072
rect 266446 55060 266452 55072
rect 219308 55032 266452 55060
rect 219308 55020 219314 55032
rect 266446 55020 266452 55032
rect 266504 55020 266510 55072
rect 375190 55020 375196 55072
rect 375248 55060 375254 55072
rect 431954 55060 431960 55072
rect 375248 55032 431960 55060
rect 375248 55020 375254 55032
rect 431954 55020 431960 55032
rect 432012 55020 432018 55072
rect 56962 54952 56968 55004
rect 57020 54992 57026 55004
rect 91186 54992 91192 55004
rect 57020 54964 91192 54992
rect 57020 54952 57026 54964
rect 91186 54952 91192 54964
rect 91244 54952 91250 55004
rect 219710 54952 219716 55004
rect 219768 54992 219774 55004
rect 253934 54992 253940 55004
rect 219768 54964 253940 54992
rect 219768 54952 219774 54964
rect 253934 54952 253940 54964
rect 253992 54952 253998 55004
rect 379054 54952 379060 55004
rect 379112 54992 379118 55004
rect 426526 54992 426532 55004
rect 379112 54964 426532 54992
rect 379112 54952 379118 54964
rect 426526 54952 426532 54964
rect 426584 54952 426590 55004
rect 58986 54884 58992 54936
rect 59044 54924 59050 54936
rect 92474 54924 92480 54936
rect 59044 54896 92480 54924
rect 59044 54884 59050 54896
rect 92474 54884 92480 54896
rect 92532 54884 92538 54936
rect 218882 54884 218888 54936
rect 218940 54924 218946 54936
rect 251358 54924 251364 54936
rect 218940 54896 251364 54924
rect 218940 54884 218946 54896
rect 251358 54884 251364 54896
rect 251416 54884 251422 54936
rect 378410 54884 378416 54936
rect 378468 54924 378474 54936
rect 423674 54924 423680 54936
rect 378468 54896 423680 54924
rect 378468 54884 378474 54896
rect 423674 54884 423680 54896
rect 423732 54884 423738 54936
rect 56318 54816 56324 54868
rect 56376 54856 56382 54868
rect 88334 54856 88340 54868
rect 56376 54828 88340 54856
rect 56376 54816 56382 54828
rect 88334 54816 88340 54828
rect 88392 54816 88398 54868
rect 216398 54816 216404 54868
rect 216456 54856 216462 54868
rect 248414 54856 248420 54868
rect 216456 54828 248420 54856
rect 216456 54816 216462 54828
rect 248414 54816 248420 54828
rect 248472 54816 248478 54868
rect 377214 54816 377220 54868
rect 377272 54856 377278 54868
rect 411346 54856 411352 54868
rect 377272 54828 411352 54856
rect 377272 54816 377278 54828
rect 411346 54816 411352 54828
rect 411404 54816 411410 54868
rect 56226 54748 56232 54800
rect 56284 54788 56290 54800
rect 86954 54788 86960 54800
rect 56284 54760 86960 54788
rect 56284 54748 56290 54760
rect 86954 54748 86960 54760
rect 87012 54748 87018 54800
rect 219158 54748 219164 54800
rect 219216 54788 219222 54800
rect 249794 54788 249800 54800
rect 219216 54760 249800 54788
rect 219216 54748 219222 54760
rect 249794 54748 249800 54760
rect 249852 54748 249858 54800
rect 377306 54748 377312 54800
rect 377364 54788 377370 54800
rect 409874 54788 409880 54800
rect 377364 54760 409880 54788
rect 377364 54748 377370 54760
rect 409874 54748 409880 54760
rect 409932 54748 409938 54800
rect 53374 54680 53380 54732
rect 53432 54720 53438 54732
rect 81434 54720 81440 54732
rect 53432 54692 81440 54720
rect 53432 54680 53438 54692
rect 81434 54680 81440 54692
rect 81492 54680 81498 54732
rect 217226 54680 217232 54732
rect 217284 54720 217290 54732
rect 245654 54720 245660 54732
rect 217284 54692 245660 54720
rect 217284 54680 217290 54692
rect 245654 54680 245660 54692
rect 245712 54680 245718 54732
rect 376294 54680 376300 54732
rect 376352 54720 376358 54732
rect 407114 54720 407120 54732
rect 376352 54692 407120 54720
rect 376352 54680 376358 54692
rect 407114 54680 407120 54692
rect 407172 54680 407178 54732
rect 52086 54612 52092 54664
rect 52144 54652 52150 54664
rect 78674 54652 78680 54664
rect 52144 54624 78680 54652
rect 52144 54612 52150 54624
rect 78674 54612 78680 54624
rect 78732 54612 78738 54664
rect 213362 54612 213368 54664
rect 213420 54652 213426 54664
rect 241514 54652 241520 54664
rect 213420 54624 241520 54652
rect 213420 54612 213426 54624
rect 241514 54612 241520 54624
rect 241572 54612 241578 54664
rect 376110 54612 376116 54664
rect 376168 54652 376174 54664
rect 404354 54652 404360 54664
rect 376168 54624 404360 54652
rect 376168 54612 376174 54624
rect 404354 54612 404360 54624
rect 404412 54612 404418 54664
rect 216306 54544 216312 54596
rect 216364 54584 216370 54596
rect 242894 54584 242900 54596
rect 216364 54556 242900 54584
rect 216364 54544 216370 54556
rect 242894 54544 242900 54556
rect 242952 54544 242958 54596
rect 378778 54544 378784 54596
rect 378836 54584 378842 54596
rect 405826 54584 405832 54596
rect 378836 54556 405832 54584
rect 378836 54544 378842 54556
rect 405826 54544 405832 54556
rect 405884 54544 405890 54596
rect 214834 54476 214840 54528
rect 214892 54516 214898 54528
rect 271874 54516 271880 54528
rect 214892 54488 271880 54516
rect 214892 54476 214898 54488
rect 271874 54476 271880 54488
rect 271932 54476 271938 54528
rect 374914 54476 374920 54528
rect 374972 54516 374978 54528
rect 401594 54516 401600 54528
rect 374972 54488 401600 54516
rect 374972 54476 374978 54488
rect 401594 54476 401600 54488
rect 401652 54476 401658 54528
rect 214190 54408 214196 54460
rect 214248 54448 214254 54460
rect 269114 54448 269120 54460
rect 214248 54420 269120 54448
rect 214248 54408 214254 54420
rect 269114 54408 269120 54420
rect 269172 54408 269178 54460
rect 374822 54408 374828 54460
rect 374880 54448 374886 54460
rect 398834 54448 398840 54460
rect 374880 54420 398840 54448
rect 374880 54408 374886 54420
rect 398834 54408 398840 54420
rect 398892 54408 398898 54460
rect 213454 54340 213460 54392
rect 213512 54380 213518 54392
rect 238754 54380 238760 54392
rect 213512 54352 238760 54380
rect 213512 54340 213518 54352
rect 238754 54340 238760 54352
rect 238812 54340 238818 54392
rect 216490 54272 216496 54324
rect 216548 54312 216554 54324
rect 236086 54312 236092 54324
rect 216548 54284 236092 54312
rect 216548 54272 216554 54284
rect 236086 54272 236092 54284
rect 236144 54272 236150 54324
rect 2774 20340 2780 20392
rect 2832 20380 2838 20392
rect 4798 20380 4804 20392
rect 2832 20352 4804 20380
rect 2832 20340 2838 20352
rect 4798 20340 4804 20352
rect 4856 20340 4862 20392
rect 147122 3476 147128 3528
rect 147180 3516 147186 3528
rect 363598 3516 363604 3528
rect 147180 3488 363604 3516
rect 147180 3476 147186 3488
rect 363598 3476 363604 3488
rect 363656 3476 363662 3528
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 57238 3448 57244 3460
rect 624 3420 57244 3448
rect 624 3408 630 3420
rect 57238 3408 57244 3420
rect 57296 3408 57302 3460
rect 125870 3408 125876 3460
rect 125928 3448 125934 3460
rect 366358 3448 366364 3460
rect 125928 3420 366364 3448
rect 125928 3408 125934 3420
rect 366358 3408 366364 3420
rect 366416 3408 366422 3460
<< via1 >>
rect 235172 700340 235224 700392
rect 307024 700340 307076 700392
rect 429844 700340 429896 700392
rect 434720 700340 434772 700392
rect 170312 700272 170364 700324
rect 434812 700272 434864 700324
rect 364340 692044 364392 692096
rect 427820 692044 427872 692096
rect 147312 683136 147364 683188
rect 580172 683136 580224 683188
rect 59176 654780 59228 654832
rect 542360 654780 542412 654832
rect 104900 653352 104952 653404
rect 434904 653352 434956 653404
rect 299480 651992 299532 652044
rect 405832 651992 405884 652044
rect 324228 649272 324280 649324
rect 494060 649272 494112 649324
rect 311164 648116 311216 648168
rect 337568 648116 337620 648168
rect 316776 648048 316828 648100
rect 342260 648048 342312 648100
rect 323768 647980 323820 648032
rect 401692 647980 401744 648032
rect 322388 647912 322440 647964
rect 346584 647912 346636 647964
rect 322296 647844 322348 647896
rect 355600 647844 355652 647896
rect 323584 647776 323636 647828
rect 369124 647776 369176 647828
rect 318156 647708 318208 647760
rect 364616 647708 364668 647760
rect 320916 647640 320968 647692
rect 374000 647640 374052 647692
rect 324872 647572 324924 647624
rect 378140 647572 378192 647624
rect 324780 647504 324832 647556
rect 387800 647504 387852 647556
rect 313924 647436 313976 647488
rect 383660 647436 383712 647488
rect 320824 647368 320876 647420
rect 392308 647368 392360 647420
rect 322204 647300 322256 647352
rect 432880 647300 432932 647352
rect 323676 647232 323728 647284
rect 328552 647232 328604 647284
rect 391940 647232 391992 647284
rect 396816 647232 396868 647284
rect 419540 647232 419592 647284
rect 457444 647232 457496 647284
rect 235080 646484 235132 646536
rect 391940 646484 391992 646536
rect 322572 646416 322624 646468
rect 436192 646416 436244 646468
rect 322480 646348 322532 646400
rect 436100 646348 436152 646400
rect 319444 646280 319496 646332
rect 436284 646280 436336 646332
rect 234344 646212 234396 646264
rect 360200 646212 360252 646264
rect 316868 646144 316920 646196
rect 457536 646144 457588 646196
rect 319536 646076 319588 646128
rect 494796 646076 494848 646128
rect 239404 646008 239456 646060
rect 433340 646008 433392 646060
rect 18604 645940 18656 645992
rect 414848 645940 414900 645992
rect 238024 645872 238076 645924
rect 419540 645872 419592 645924
rect 147496 645328 147548 645380
rect 164516 645328 164568 645380
rect 145472 645260 145524 645312
rect 144920 645124 144972 645176
rect 156604 645124 156656 645176
rect 196072 645124 196124 645176
rect 238852 645124 238904 645176
rect 580356 645124 580408 645176
rect 142804 645056 142856 645108
rect 161480 645056 161532 645108
rect 215024 645056 215076 645108
rect 245660 645056 245712 645108
rect 322664 645056 322716 645108
rect 457720 645056 457772 645108
rect 115388 644988 115440 645040
rect 124588 644988 124640 645040
rect 148784 644988 148836 645040
rect 86408 644920 86460 644972
rect 124220 644920 124272 644972
rect 148968 644920 149020 644972
rect 156420 644920 156472 644972
rect 94780 644852 94832 644904
rect 120908 644852 120960 644904
rect 147588 644852 147640 644904
rect 155224 644852 155276 644904
rect 156696 644988 156748 645040
rect 207664 644988 207716 645040
rect 226432 644988 226484 645040
rect 300308 644988 300360 645040
rect 314108 644988 314160 645040
rect 456984 644988 457036 645040
rect 156604 644920 156656 644972
rect 172888 644920 172940 644972
rect 214288 644920 214340 644972
rect 289268 644920 289320 644972
rect 318064 644920 318116 644972
rect 471612 644920 471664 644972
rect 176108 644852 176160 644904
rect 232504 644852 232556 644904
rect 271972 644852 272024 644904
rect 304264 644852 304316 644904
rect 457628 644852 457680 644904
rect 106372 644784 106424 644836
rect 121644 644784 121696 644836
rect 143356 644784 143408 644836
rect 184480 644784 184532 644836
rect 231124 644784 231176 644836
rect 248788 644784 248840 644836
rect 249156 644784 249208 644836
rect 295524 644784 295576 644836
rect 314016 644784 314068 644836
rect 483204 644784 483256 644836
rect 109592 644716 109644 644768
rect 126980 644716 127032 644768
rect 149704 644716 149756 644768
rect 190460 644716 190512 644768
rect 222936 644716 222988 644768
rect 277676 644716 277728 644768
rect 319628 644716 319680 644768
rect 512000 644716 512052 644768
rect 55128 644648 55180 644700
rect 80612 644648 80664 644700
rect 103796 644648 103848 644700
rect 121460 644648 121512 644700
rect 149796 644648 149848 644700
rect 199292 644648 199344 644700
rect 239680 644648 239732 644700
rect 297732 644648 297784 644700
rect 316960 644648 317012 644700
rect 512092 644648 512144 644700
rect 54944 644580 54996 644632
rect 92204 644580 92256 644632
rect 100576 644580 100628 644632
rect 124404 644580 124456 644632
rect 148876 644580 148928 644632
rect 55036 644512 55088 644564
rect 88984 644512 89036 644564
rect 112168 644512 112220 644564
rect 121000 644512 121052 644564
rect 148416 644512 148468 644564
rect 153200 644512 153252 644564
rect 155224 644512 155276 644564
rect 158720 644512 158772 644564
rect 239588 644580 239640 644632
rect 251364 644580 251416 644632
rect 317052 644580 317104 644632
rect 512184 644580 512236 644632
rect 201868 644512 201920 644564
rect 237472 644512 237524 644564
rect 254492 644512 254544 644564
rect 305644 644512 305696 644564
rect 501236 644512 501288 644564
rect 59360 644444 59412 644496
rect 98000 644444 98052 644496
rect 117964 644444 118016 644496
rect 124496 644444 124548 644496
rect 134064 644444 134116 644496
rect 149980 644444 150032 644496
rect 205548 644444 205600 644496
rect 211160 644444 211212 644496
rect 239496 644444 239548 644496
rect 242900 644444 242952 644496
rect 3424 643696 3476 643748
rect 321008 643696 321060 643748
rect 238116 643560 238168 643612
rect 268660 643560 268712 643612
rect 126244 643492 126296 643544
rect 187700 643492 187752 643544
rect 220084 643492 220136 643544
rect 257068 643492 257120 643544
rect 149888 643424 149940 643476
rect 170312 643424 170364 643476
rect 228364 643424 228416 643476
rect 266544 643424 266596 643476
rect 56324 643356 56376 643408
rect 71596 643356 71648 643408
rect 141884 643356 141936 643408
rect 167092 643356 167144 643408
rect 220176 643356 220228 643408
rect 260380 643356 260432 643408
rect 56508 643288 56560 643340
rect 65800 643288 65852 643340
rect 137652 643288 137704 643340
rect 179006 643288 179058 643340
rect 231216 643288 231268 643340
rect 280252 643288 280304 643340
rect 59268 643220 59320 643272
rect 74816 643220 74868 643272
rect 144184 643220 144236 643272
rect 193818 643220 193870 643272
rect 236644 643220 236696 643272
rect 291844 643220 291896 643272
rect 56416 643152 56468 643204
rect 77392 643152 77444 643204
rect 83188 643152 83240 643204
rect 124312 643152 124364 643204
rect 125416 643152 125468 643204
rect 182226 643152 182278 643204
rect 215944 643152 215996 643204
rect 274640 643152 274692 643204
rect 69296 643084 69348 643136
rect 122840 643084 122892 643136
rect 146116 643084 146168 643136
rect 155500 643084 155552 643136
rect 217324 643084 217376 643136
rect 286140 643084 286192 643136
rect 312544 643084 312596 643136
rect 321560 643084 321612 643136
rect 54852 642336 54904 642388
rect 62948 642336 63000 642388
rect 223580 642336 223632 642388
rect 249156 642336 249208 642388
rect 222844 641860 222896 641912
rect 262956 642336 263008 642388
rect 214564 641792 214616 641844
rect 283564 642336 283616 642388
rect 57888 641724 57940 641776
rect 146208 641724 146260 641776
rect 238024 641724 238076 641776
rect 140044 640296 140096 640348
rect 146300 640296 146352 640348
rect 235264 640296 235316 640348
rect 237380 640296 237432 640348
rect 465172 640296 465224 640348
rect 580264 640296 580316 640348
rect 309876 638936 309928 638988
rect 321560 638936 321612 638988
rect 238944 638596 238996 638648
rect 239772 638596 239824 638648
rect 215760 638188 215812 638240
rect 237472 638188 237524 638240
rect 233608 633428 233660 633480
rect 237380 633428 237432 633480
rect 307116 633428 307168 633480
rect 321560 633428 321612 633480
rect 141240 630640 141292 630692
rect 146300 630640 146352 630692
rect 232596 630640 232648 630692
rect 237380 630640 237432 630692
rect 309784 629280 309836 629332
rect 321560 629280 321612 629332
rect 132592 627920 132644 627972
rect 146300 627920 146352 627972
rect 224316 625132 224368 625184
rect 237380 625132 237432 625184
rect 305736 625132 305788 625184
rect 321560 625132 321612 625184
rect 218612 620984 218664 621036
rect 237380 620984 237432 621036
rect 312636 619624 312688 619676
rect 321560 619624 321612 619676
rect 314200 615476 314252 615528
rect 321560 615476 321612 615528
rect 233884 612756 233936 612808
rect 237380 612756 237432 612808
rect 129096 609968 129148 610020
rect 146300 609968 146352 610020
rect 217416 609968 217468 610020
rect 237380 609968 237432 610020
rect 311256 609968 311308 610020
rect 321560 609968 321612 610020
rect 302792 609220 302844 609272
rect 303160 609220 303212 609272
rect 322664 609220 322716 609272
rect 124036 608608 124088 608660
rect 145564 608608 145616 608660
rect 220268 607180 220320 607232
rect 237380 607180 237432 607232
rect 229744 603100 229796 603152
rect 237380 603100 237432 603152
rect 232872 600312 232924 600364
rect 237380 600312 237432 600364
rect 308404 600312 308456 600364
rect 321560 600312 321612 600364
rect 126888 597524 126940 597576
rect 146300 597524 146352 597576
rect 235356 597524 235408 597576
rect 237380 597524 237432 597576
rect 305828 596164 305880 596216
rect 321560 596164 321612 596216
rect 144276 594804 144328 594856
rect 146944 594804 146996 594856
rect 216036 594804 216088 594856
rect 237380 594804 237432 594856
rect 513288 592016 513340 592068
rect 578884 592016 578936 592068
rect 139768 590656 139820 590708
rect 146300 590656 146352 590708
rect 217508 590656 217560 590708
rect 237380 590656 237432 590708
rect 317144 590656 317196 590708
rect 321560 590656 321612 590708
rect 227168 587868 227220 587920
rect 237380 587868 237432 587920
rect 219256 585148 219308 585200
rect 237380 585148 237432 585200
rect 123116 584944 123168 584996
rect 123576 584944 123628 584996
rect 148324 583040 148376 583092
rect 148784 583040 148836 583092
rect 148784 582904 148836 582956
rect 148968 582904 149020 582956
rect 223488 582360 223540 582412
rect 237380 582360 237432 582412
rect 120724 581748 120776 581800
rect 121184 581748 121236 581800
rect 57428 581204 57480 581256
rect 59912 581204 59964 581256
rect 3148 580932 3200 580984
rect 305828 580932 305880 580984
rect 145564 580864 145616 580916
rect 213920 580864 213972 580916
rect 302792 580864 302844 580916
rect 58808 580660 58860 580712
rect 60924 580660 60976 580712
rect 119344 580660 119396 580712
rect 123116 580660 123168 580712
rect 147128 580660 147180 580712
rect 151084 580660 151136 580712
rect 57336 580592 57388 580644
rect 61384 580592 61436 580644
rect 112536 580252 112588 580304
rect 123576 580252 123628 580304
rect 199384 580252 199436 580304
rect 212632 580252 212684 580304
rect 59176 579572 59228 579624
rect 62396 579572 62448 579624
rect 148600 579572 148652 579624
rect 150532 579572 150584 579624
rect 295248 579572 295300 579624
rect 319628 579572 319680 579624
rect 289544 579504 289596 579556
rect 316868 579504 316920 579556
rect 107568 579436 107620 579488
rect 124588 579436 124640 579488
rect 288808 579436 288860 579488
rect 317052 579436 317104 579488
rect 97448 579368 97500 579420
rect 121000 579368 121052 579420
rect 288072 579368 288124 579420
rect 316960 579368 317012 579420
rect 98184 579300 98236 579352
rect 126980 579300 127032 579352
rect 148876 579300 148928 579352
rect 155500 579300 155552 579352
rect 286324 579300 286376 579352
rect 319444 579300 319496 579352
rect 93952 579232 94004 579284
rect 124404 579232 124456 579284
rect 149796 579232 149848 579284
rect 156236 579232 156288 579284
rect 165528 579232 165580 579284
rect 211160 579232 211212 579284
rect 258724 579232 258776 579284
rect 322480 579232 322532 579284
rect 58440 579164 58492 579216
rect 68836 579164 68888 579216
rect 87420 579164 87472 579216
rect 121644 579164 121696 579216
rect 123116 579164 123168 579216
rect 211712 579164 211764 579216
rect 245844 579164 245896 579216
rect 322572 579164 322624 579216
rect 57704 579096 57756 579148
rect 71044 579096 71096 579148
rect 88156 579096 88208 579148
rect 124496 579096 124548 579148
rect 148968 579096 149020 579148
rect 159088 579096 159140 579148
rect 200672 579096 200724 579148
rect 301412 579096 301464 579148
rect 57612 579028 57664 579080
rect 83188 579028 83240 579080
rect 84568 579028 84620 579080
rect 122104 579028 122156 579080
rect 148324 579028 148376 579080
rect 161940 579028 161992 579080
rect 196348 579028 196400 579080
rect 302608 579028 302660 579080
rect 66720 578960 66772 579012
rect 120724 578960 120776 579012
rect 148784 578960 148836 579012
rect 164884 578960 164936 579012
rect 184204 578960 184256 579012
rect 301044 578960 301096 579012
rect 63776 578892 63828 578944
rect 122288 578892 122340 578944
rect 149704 578892 149756 578944
rect 151820 578892 151872 578944
rect 179880 578892 179932 578944
rect 301596 578892 301648 578944
rect 147220 578824 147272 578876
rect 166264 578824 166316 578876
rect 290188 578824 290240 578876
rect 314016 578824 314068 578876
rect 297364 578756 297416 578808
rect 319536 578756 319588 578808
rect 292396 578688 292448 578740
rect 314108 578688 314160 578740
rect 106924 578144 106976 578196
rect 108580 578144 108632 578196
rect 116584 578144 116636 578196
rect 117412 578144 117464 578196
rect 191104 578144 191156 578196
rect 195428 578144 195480 578196
rect 192484 578076 192536 578128
rect 198740 578076 198792 578128
rect 174176 577940 174228 577992
rect 189632 577940 189684 577992
rect 162676 577872 162728 577924
rect 178040 577872 178092 577924
rect 164148 577804 164200 577856
rect 183836 577804 183888 577856
rect 227904 577804 227956 577856
rect 265532 577804 265584 577856
rect 77024 577736 77076 577788
rect 86776 577736 86828 577788
rect 94504 577736 94556 577788
rect 104164 577736 104216 577788
rect 150348 577736 150400 577788
rect 151176 577736 151228 577788
rect 154856 577736 154908 577788
rect 181260 577736 181312 577788
rect 232228 577736 232280 577788
rect 279700 577736 279752 577788
rect 60280 577668 60332 577720
rect 71136 577668 71188 577720
rect 75276 577668 75328 577720
rect 96988 577668 97040 577720
rect 100208 577668 100260 577720
rect 115204 577668 115256 577720
rect 159824 577668 159876 577720
rect 192852 577668 192904 577720
rect 198004 577668 198056 577720
rect 210240 577668 210292 577720
rect 220728 577668 220780 577720
rect 268108 577668 268160 577720
rect 273904 577668 273956 577720
rect 282920 577668 282972 577720
rect 289084 577668 289136 577720
rect 300308 577668 300360 577720
rect 58900 577600 58952 577652
rect 74540 577600 74592 577652
rect 86040 577600 86092 577652
rect 108304 577600 108356 577652
rect 116676 577600 116728 577652
rect 120172 577600 120224 577652
rect 130476 577600 130528 577652
rect 163872 577600 163924 577652
rect 169852 577600 169904 577652
rect 175464 577600 175516 577652
rect 183468 577600 183520 577652
rect 232504 577600 232556 577652
rect 235448 577600 235500 577652
rect 242348 577600 242400 577652
rect 249064 577600 249116 577652
rect 259644 577600 259696 577652
rect 280804 577600 280856 577652
rect 296996 577600 297048 577652
rect 68744 577532 68796 577584
rect 105544 577532 105596 577584
rect 133328 577532 133380 577584
rect 187056 577532 187108 577584
rect 195244 577532 195296 577584
rect 212724 577532 212776 577584
rect 222200 577532 222252 577584
rect 273812 577532 273864 577584
rect 280896 577532 280948 577584
rect 322388 577532 322440 577584
rect 71320 577464 71372 577516
rect 108396 577464 108448 577516
rect 110420 577464 110472 577516
rect 121184 577464 121236 577516
rect 134708 577464 134760 577516
rect 207020 577464 207072 577516
rect 217140 577464 217192 577516
rect 223488 577464 223540 577516
rect 231308 577464 231360 577516
rect 239772 577464 239824 577516
rect 257988 577464 258040 577516
rect 324780 577464 324832 577516
rect 202236 577192 202288 577244
rect 204444 577192 204496 577244
rect 269764 577192 269816 577244
rect 271236 577192 271288 577244
rect 242164 576920 242216 576972
rect 248512 576920 248564 576972
rect 64144 576852 64196 576904
rect 64972 576852 65024 576904
rect 199476 576852 199528 576904
rect 201500 576852 201552 576904
rect 244924 576852 244976 576904
rect 250628 576852 250680 576904
rect 282184 576852 282236 576904
rect 288716 576852 288768 576904
rect 160744 576376 160796 576428
rect 213000 576376 213052 576428
rect 122564 576308 122616 576360
rect 211252 576308 211304 576360
rect 228640 576308 228692 576360
rect 300952 576308 301004 576360
rect 57244 576240 57296 576292
rect 79324 576240 79376 576292
rect 91100 576240 91152 576292
rect 96804 576240 96856 576292
rect 100392 576240 100444 576292
rect 123300 576240 123352 576292
rect 206284 576240 206336 576292
rect 302976 576240 303028 576292
rect 65248 576172 65300 576224
rect 122012 576172 122064 576224
rect 180616 576172 180668 576224
rect 300860 576172 300912 576224
rect 3424 576104 3476 576156
rect 323860 576104 323912 576156
rect 128268 574948 128320 575000
rect 211804 574948 211856 575000
rect 266544 574948 266596 575000
rect 322296 574948 322348 575000
rect 58624 574880 58676 574932
rect 91008 574880 91060 574932
rect 187792 574880 187844 574932
rect 302332 574880 302384 574932
rect 70308 574812 70360 574864
rect 122196 574812 122248 574864
rect 181352 574812 181404 574864
rect 301320 574812 301372 574864
rect 4804 574744 4856 574796
rect 321836 574744 321888 574796
rect 204260 573520 204312 573572
rect 239680 573520 239732 573572
rect 59084 573452 59136 573504
rect 92480 573452 92532 573504
rect 177028 573452 177080 573504
rect 217416 573452 217468 573504
rect 240784 573452 240836 573504
rect 320916 573452 320968 573504
rect 59452 573384 59504 573436
rect 76012 573384 76064 573436
rect 80336 573384 80388 573436
rect 120816 573384 120868 573436
rect 126152 573384 126204 573436
rect 211344 573384 211396 573436
rect 216404 573384 216456 573436
rect 301504 573384 301556 573436
rect 64512 573316 64564 573368
rect 122932 573316 122984 573368
rect 181996 573316 182048 573368
rect 301136 573316 301188 573368
rect 68100 572228 68152 572280
rect 121828 572228 121880 572280
rect 189908 572228 189960 572280
rect 239588 572228 239640 572280
rect 139032 572160 139084 572212
rect 213092 572160 213144 572212
rect 121828 572092 121880 572144
rect 211896 572092 211948 572144
rect 267280 572092 267332 572144
rect 313924 572092 313976 572144
rect 70952 572024 71004 572076
rect 121920 572024 121972 572076
rect 209780 572024 209832 572076
rect 301228 572024 301280 572076
rect 65984 571956 66036 572008
rect 123208 571956 123260 572008
rect 147036 571956 147088 572008
rect 169116 571956 169168 572008
rect 194968 571956 195020 572008
rect 302884 571956 302936 572008
rect 268016 571344 268068 571396
rect 321560 571344 321612 571396
rect 192116 570800 192168 570852
rect 238944 570800 238996 570852
rect 269488 570800 269540 570852
rect 317144 570800 317196 570852
rect 136916 570732 136968 570784
rect 213184 570732 213236 570784
rect 253664 570732 253716 570784
rect 323768 570732 323820 570784
rect 57520 570664 57572 570716
rect 87604 570664 87656 570716
rect 89628 570664 89680 570716
rect 104900 570664 104952 570716
rect 119712 570664 119764 570716
rect 154672 570664 154724 570716
rect 197084 570664 197136 570716
rect 302700 570664 302752 570716
rect 78864 570596 78916 570648
rect 123484 570596 123536 570648
rect 185584 570596 185636 570648
rect 293960 570596 294012 570648
rect 81440 569304 81492 569356
rect 90364 569304 90416 569356
rect 98644 569304 98696 569356
rect 123392 569304 123444 569356
rect 204996 569304 205048 569356
rect 239496 569304 239548 569356
rect 274456 569304 274508 569356
rect 322204 569304 322256 569356
rect 80980 569236 81032 569288
rect 121092 569236 121144 569288
rect 178500 569236 178552 569288
rect 216036 569236 216088 569288
rect 250812 569236 250864 569288
rect 323676 569236 323728 569288
rect 57152 569168 57204 569220
rect 103244 569168 103296 569220
rect 124036 569168 124088 569220
rect 211528 569168 211580 569220
rect 229284 569168 229336 569220
rect 303068 569168 303120 569220
rect 199200 567944 199252 567996
rect 232596 567944 232648 567996
rect 263692 567944 263744 567996
rect 311164 567944 311216 567996
rect 78680 567876 78732 567928
rect 115388 567876 115440 567928
rect 147036 567876 147088 567928
rect 212816 567876 212868 567928
rect 247960 567876 248012 567928
rect 324872 567876 324924 567928
rect 57060 567808 57112 567860
rect 101036 567808 101088 567860
rect 205640 567808 205692 567860
rect 285864 567808 285916 567860
rect 3424 567196 3476 567248
rect 321560 567196 321612 567248
rect 177764 566652 177816 566704
rect 244280 566652 244332 566704
rect 259460 566652 259512 566704
rect 312544 566652 312596 566704
rect 129004 566584 129056 566636
rect 211436 566584 211488 566636
rect 250076 566584 250128 566636
rect 314200 566584 314252 566636
rect 86040 566516 86092 566568
rect 121552 566516 121604 566568
rect 151176 566516 151228 566568
rect 163412 566516 163464 566568
rect 191380 566516 191432 566568
rect 277400 566516 277452 566568
rect 279516 566516 279568 566568
rect 307116 566516 307168 566568
rect 58992 566448 59044 566500
rect 102508 566448 102560 566500
rect 160100 566448 160152 566500
rect 172704 566448 172756 566500
rect 198556 566448 198608 566500
rect 289084 566448 289136 566500
rect 202788 565292 202840 565344
rect 256700 565292 256752 565344
rect 152648 565224 152700 565276
rect 212908 565224 212960 565276
rect 275192 565224 275244 565276
rect 316776 565224 316828 565276
rect 124680 565156 124732 565208
rect 210884 565156 210936 565208
rect 246488 565156 246540 565208
rect 305736 565156 305788 565208
rect 71136 565088 71188 565140
rect 105360 565088 105412 565140
rect 149060 565088 149112 565140
rect 161296 565088 161348 565140
rect 179144 565088 179196 565140
rect 291200 565088 291252 565140
rect 193496 563864 193548 563916
rect 235264 563864 235316 563916
rect 245108 563864 245160 563916
rect 318156 563864 318208 563916
rect 82452 563796 82504 563848
rect 116676 563796 116728 563848
rect 142620 563796 142672 563848
rect 211620 563796 211672 563848
rect 242900 563796 242952 563848
rect 320824 563796 320876 563848
rect 62212 563728 62264 563780
rect 109684 563728 109736 563780
rect 131212 563728 131264 563780
rect 192484 563728 192536 563780
rect 192760 563728 192812 563780
rect 280804 563728 280856 563780
rect 71688 563660 71740 563712
rect 121736 563660 121788 563712
rect 187056 563660 187108 563712
rect 302424 563660 302476 563712
rect 40040 562980 40092 563032
rect 321560 562980 321612 563032
rect 207112 562436 207164 562488
rect 229744 562436 229796 562488
rect 88340 562368 88392 562420
rect 104624 562368 104676 562420
rect 158352 562368 158404 562420
rect 213276 562368 213328 562420
rect 57796 562300 57848 562352
rect 116676 562300 116728 562352
rect 147312 562300 147364 562352
rect 174912 562300 174964 562352
rect 189172 562300 189224 562352
rect 282184 562300 282236 562352
rect 169852 562164 169904 562216
rect 170036 562164 170088 562216
rect 121092 561076 121144 561128
rect 199476 561076 199528 561128
rect 206376 561076 206428 561128
rect 262220 561076 262272 561128
rect 76748 561008 76800 561060
rect 116584 561008 116636 561060
rect 129740 561008 129792 561060
rect 212540 561008 212592 561060
rect 251548 561008 251600 561060
rect 323584 561008 323636 561060
rect 63132 560940 63184 560992
rect 110512 560940 110564 560992
rect 182732 560940 182784 560992
rect 300676 560940 300728 560992
rect 217876 559716 217928 559768
rect 273904 559716 273956 559768
rect 73252 559648 73304 559700
rect 106924 559648 106976 559700
rect 197820 559648 197872 559700
rect 217508 559648 217560 559700
rect 256516 559648 256568 559700
rect 316684 559648 316736 559700
rect 69572 559580 69624 559632
rect 114560 559580 114612 559632
rect 120448 559580 120500 559632
rect 144276 559580 144328 559632
rect 148692 559580 148744 559632
rect 160560 559580 160612 559632
rect 184940 559580 184992 559632
rect 235356 559580 235408 559632
rect 260104 559580 260156 559632
rect 321100 559580 321152 559632
rect 58716 559512 58768 559564
rect 111064 559512 111116 559564
rect 140504 559512 140556 559564
rect 198004 559512 198056 559564
rect 202144 559512 202196 559564
rect 302240 559512 302292 559564
rect 148508 558832 148560 558884
rect 149796 558832 149848 558884
rect 208584 558356 208636 558408
rect 238208 558356 238260 558408
rect 148324 558288 148376 558340
rect 172520 558288 172572 558340
rect 190644 558288 190696 558340
rect 238300 558288 238352 558340
rect 283748 558288 283800 558340
rect 312636 558288 312688 558340
rect 147404 558220 147456 558272
rect 169760 558220 169812 558272
rect 171324 558220 171376 558272
rect 210792 558220 210844 558272
rect 212816 558220 212868 558272
rect 269764 558220 269816 558272
rect 271604 558220 271656 558272
rect 309876 558220 309928 558272
rect 58532 558152 58584 558204
rect 108212 558152 108264 558204
rect 131856 558152 131908 558204
rect 142804 558152 142856 558204
rect 144736 558152 144788 558204
rect 165712 558152 165764 558204
rect 168380 558152 168432 558204
rect 210700 558152 210752 558204
rect 212172 558152 212224 558204
rect 302516 558152 302568 558204
rect 287336 557880 287388 557932
rect 316776 557880 316828 557932
rect 283104 557812 283156 557864
rect 319444 557812 319496 557864
rect 284944 557744 284996 557796
rect 322204 557744 322256 557796
rect 252284 557676 252336 557728
rect 321560 557676 321612 557728
rect 248696 557608 248748 557660
rect 319720 557608 319772 557660
rect 237932 557540 237984 557592
rect 322296 557540 322348 557592
rect 146944 557132 146996 557184
rect 148416 557132 148468 557184
rect 147680 556996 147732 557048
rect 191104 556996 191156 557048
rect 211436 556996 211488 557048
rect 220268 556996 220320 557048
rect 176292 556928 176344 556980
rect 222936 556928 222988 556980
rect 188528 556860 188580 556912
rect 253940 556860 253992 556912
rect 282368 556860 282420 556912
rect 308404 556860 308456 556912
rect 94596 556792 94648 556844
rect 123024 556792 123076 556844
rect 127624 556792 127676 556844
rect 202236 556792 202288 556844
rect 207848 556792 207900 556844
rect 233884 556792 233936 556844
rect 270132 556792 270184 556844
rect 311256 556792 311308 556844
rect 291660 556656 291712 556708
rect 316868 556656 316920 556708
rect 285220 556588 285272 556640
rect 316684 556588 316736 556640
rect 255872 556520 255924 556572
rect 304356 556520 304408 556572
rect 273720 556452 273772 556504
rect 323676 556452 323728 556504
rect 264428 556384 264480 556436
rect 320824 556384 320876 556436
rect 265900 556316 265952 556368
rect 324872 556316 324924 556368
rect 263048 556248 263100 556300
rect 323584 556248 323636 556300
rect 135444 556180 135496 556232
rect 140044 556180 140096 556232
rect 148232 556180 148284 556232
rect 149060 556180 149112 556232
rect 254400 556180 254452 556232
rect 318156 556180 318208 556232
rect 136180 556112 136232 556164
rect 144184 556112 144236 556164
rect 169944 556112 169996 556164
rect 173440 556112 173492 556164
rect 54944 556044 54996 556096
rect 67364 556044 67416 556096
rect 71044 556044 71096 556096
rect 77392 556044 77444 556096
rect 108396 556044 108448 556096
rect 114652 556044 114704 556096
rect 151084 556044 151136 556096
rect 153384 556044 153436 556096
rect 55036 555976 55088 556028
rect 79600 555976 79652 556028
rect 54852 555908 54904 555960
rect 88892 555908 88944 555960
rect 203524 555908 203576 555960
rect 217324 555908 217376 555960
rect 60372 555840 60424 555892
rect 95332 555840 95384 555892
rect 118240 555840 118292 555892
rect 126244 555840 126296 555892
rect 201408 555840 201460 555892
rect 215944 555840 215996 555892
rect 225788 555840 225840 555892
rect 235448 555840 235500 555892
rect 56416 555772 56468 555824
rect 83924 555772 83976 555824
rect 85304 555772 85356 555824
rect 120908 555772 120960 555824
rect 157340 555772 157392 555824
rect 167000 555772 167052 555824
rect 186320 555772 186372 555824
rect 206284 555772 206336 555824
rect 209228 555772 209280 555824
rect 220176 555772 220228 555824
rect 221464 555772 221516 555824
rect 231308 555772 231360 555824
rect 55128 555704 55180 555756
rect 93216 555704 93268 555756
rect 114008 555704 114060 555756
rect 122840 555704 122892 555756
rect 146116 555704 146168 555756
rect 156972 555704 157024 555756
rect 199936 555704 199988 555756
rect 220084 555704 220136 555756
rect 230756 555704 230808 555756
rect 244924 555704 244976 555756
rect 278044 555704 278096 555756
rect 300308 555704 300360 555756
rect 59268 555636 59320 555688
rect 99656 555636 99708 555688
rect 106832 555636 106884 555688
rect 124312 555636 124364 555688
rect 147496 555636 147548 555688
rect 157708 555636 157760 555688
rect 169760 555636 169812 555688
rect 175556 555636 175608 555688
rect 194232 555636 194284 555688
rect 214564 555636 214616 555688
rect 225052 555636 225104 555688
rect 242164 555636 242216 555688
rect 270868 555636 270920 555688
rect 324688 555636 324740 555688
rect 56508 555568 56560 555620
rect 98920 555568 98972 555620
rect 103980 555568 104032 555620
rect 124220 555568 124272 555620
rect 152004 555568 152056 555620
rect 167736 555568 167788 555620
rect 170588 555568 170640 555620
rect 199384 555568 199436 555620
rect 209964 555568 210016 555620
rect 231216 555568 231268 555620
rect 231492 555568 231544 555620
rect 249064 555568 249116 555620
rect 252928 555568 252980 555620
rect 323768 555568 323820 555620
rect 61660 555500 61712 555552
rect 64144 555500 64196 555552
rect 56324 555364 56376 555416
rect 73804 555500 73856 555552
rect 78128 555500 78180 555552
rect 121460 555500 121512 555552
rect 138296 555500 138348 555552
rect 147036 555500 147088 555552
rect 147588 555500 147640 555552
rect 171968 555500 172020 555552
rect 195612 555500 195664 555552
rect 238116 555500 238168 555552
rect 261576 555500 261628 555552
rect 286324 555500 286376 555552
rect 298652 555500 298704 555552
rect 302056 555500 302108 555552
rect 61384 555296 61436 555348
rect 116860 555432 116912 555484
rect 118976 555432 119028 555484
rect 129096 555432 129148 555484
rect 144092 555432 144144 555484
rect 195244 555432 195296 555484
rect 213552 555432 213604 555484
rect 236644 555432 236696 555484
rect 237196 555432 237248 555484
rect 284944 555432 284996 555484
rect 299572 555432 299624 555484
rect 318064 555432 318116 555484
rect 72424 555364 72476 555416
rect 73160 555364 73212 555416
rect 113272 555364 113324 555416
rect 119344 555364 119396 555416
rect 242256 555364 242308 555416
rect 324136 555364 324188 555416
rect 276572 555296 276624 555348
rect 300400 555296 300452 555348
rect 79324 555228 79376 555280
rect 81716 555228 81768 555280
rect 87604 555228 87656 555280
rect 91744 555228 91796 555280
rect 96068 555228 96120 555280
rect 98644 555228 98696 555280
rect 104164 555228 104216 555280
rect 106096 555228 106148 555280
rect 108304 555228 108356 555280
rect 111800 555228 111852 555280
rect 115204 555228 115256 555280
rect 116124 555228 116176 555280
rect 116676 555228 116728 555280
rect 117596 555228 117648 555280
rect 144920 555228 144972 555280
rect 146208 555228 146260 555280
rect 149888 555228 149940 555280
rect 151268 555228 151320 555280
rect 154120 555228 154172 555280
rect 160744 555228 160796 555280
rect 219992 555228 220044 555280
rect 228364 555228 228416 555280
rect 230020 555228 230072 555280
rect 231124 555228 231176 555280
rect 277308 555228 277360 555280
rect 105544 555160 105596 555212
rect 108948 555160 109000 555212
rect 275928 555160 275980 555212
rect 298652 555160 298704 555212
rect 298836 555228 298888 555280
rect 304264 555228 304316 555280
rect 301872 555160 301924 555212
rect 290924 555092 290976 555144
rect 322480 555092 322532 555144
rect 280160 555024 280212 555076
rect 322664 555024 322716 555076
rect 257252 554956 257304 555008
rect 300492 554956 300544 555008
rect 265164 554888 265216 554940
rect 274640 554888 274692 554940
rect 281632 554820 281684 554872
rect 301504 554888 301556 554940
rect 295984 554752 296036 554804
rect 301596 554820 301648 554872
rect 296812 554752 296864 554804
rect 300124 554752 300176 554804
rect 240048 554276 240100 554328
rect 303068 554276 303120 554328
rect 236460 554208 236512 554260
rect 321652 554208 321704 554260
rect 235816 554140 235868 554192
rect 324044 554140 324096 554192
rect 268752 554072 268804 554124
rect 302976 554072 303028 554124
rect 274640 554004 274692 554056
rect 324320 554004 324372 554056
rect 260840 553936 260892 553988
rect 305644 553936 305696 553988
rect 272340 553868 272392 553920
rect 324596 553868 324648 553920
rect 247224 553800 247276 553852
rect 301780 553800 301832 553852
rect 243636 553732 243688 553784
rect 300676 553732 300728 553784
rect 262312 553664 262364 553716
rect 324780 553664 324832 553716
rect 284484 553596 284536 553648
rect 319536 553596 319588 553648
rect 244372 553528 244424 553580
rect 322572 553528 322624 553580
rect 278780 553460 278832 553512
rect 299388 553460 299440 553512
rect 273076 553392 273128 553444
rect 301688 553392 301740 553444
rect 299388 553324 299440 553376
rect 321560 553324 321612 553376
rect 3516 553052 3568 553104
rect 322756 553052 322808 553104
rect 302240 545096 302292 545148
rect 304264 545096 304316 545148
rect 300676 543668 300728 543720
rect 321560 543668 321612 543720
rect 436836 543192 436888 543244
rect 436284 543056 436336 543108
rect 436836 542988 436888 543040
rect 436652 542852 436704 542904
rect 303068 539520 303120 539572
rect 321560 539520 321612 539572
rect 324136 535372 324188 535424
rect 436560 535372 436612 535424
rect 324320 534556 324372 534608
rect 325148 534556 325200 534608
rect 300216 534012 300268 534064
rect 436284 534012 436336 534064
rect 300308 533944 300360 533996
rect 436100 533944 436152 533996
rect 300492 533876 300544 533928
rect 436836 533876 436888 533928
rect 301872 533808 301924 533860
rect 436376 533808 436428 533860
rect 319720 533740 319772 533792
rect 433340 533740 433392 533792
rect 322664 533672 322716 533724
rect 434628 533672 434680 533724
rect 323768 533604 323820 533656
rect 436744 533604 436796 533656
rect 323952 533536 324004 533588
rect 436928 533536 436980 533588
rect 324688 533468 324740 533520
rect 436652 533468 436704 533520
rect 322296 533400 322348 533452
rect 433800 533400 433852 533452
rect 302056 532856 302108 532908
rect 356244 532856 356296 532908
rect 307024 532788 307076 532840
rect 374276 532788 374328 532840
rect 300400 532720 300452 532772
rect 420000 532720 420052 532772
rect 324044 532652 324096 532704
rect 338212 532652 338264 532704
rect 322572 532584 322624 532636
rect 424508 532584 424560 532636
rect 324780 532516 324832 532568
rect 334072 532516 334124 532568
rect 302976 532448 303028 532500
rect 393320 532448 393372 532500
rect 323584 532380 323636 532432
rect 406476 532380 406528 532432
rect 323676 532312 323728 532364
rect 401968 532312 402020 532364
rect 301688 532244 301740 532296
rect 369860 532244 369912 532296
rect 324872 532176 324924 532228
rect 388444 532176 388496 532228
rect 301780 532108 301832 532160
rect 365260 532108 365312 532160
rect 320824 532040 320876 532092
rect 379520 532040 379572 532092
rect 318156 531972 318208 532024
rect 351920 531972 351972 532024
rect 305644 531904 305696 531956
rect 347228 531904 347280 531956
rect 304356 531836 304408 531888
rect 411352 531836 411404 531888
rect 324596 531768 324648 531820
rect 415492 531768 415544 531820
rect 302884 531224 302936 531276
rect 495440 531224 495492 531276
rect 322388 531156 322440 531208
rect 512184 531156 512236 531208
rect 322480 531088 322532 531140
rect 488540 531088 488592 531140
rect 300124 531020 300176 531072
rect 459560 531020 459612 531072
rect 316776 530952 316828 531004
rect 476120 530952 476172 531004
rect 301596 530884 301648 530936
rect 457444 530884 457496 530936
rect 316868 530816 316920 530868
rect 457628 530816 457680 530868
rect 301504 530748 301556 530800
rect 436468 530748 436520 530800
rect 302424 529932 302476 529984
rect 520924 529932 520976 529984
rect 316960 529864 317012 529916
rect 512276 529864 512328 529916
rect 319628 529796 319680 529848
rect 500960 529796 501012 529848
rect 316684 529728 316736 529780
rect 470600 529728 470652 529780
rect 319812 529660 319864 529712
rect 465080 529660 465132 529712
rect 319444 529592 319496 529644
rect 433524 529592 433576 529644
rect 319536 529524 319588 529576
rect 433708 529524 433760 529576
rect 322204 529456 322256 529508
rect 433432 529456 433484 529508
rect 329748 529388 329800 529440
rect 434720 529388 434772 529440
rect 363604 527824 363656 527876
rect 506480 527824 506532 527876
rect 53748 521704 53800 521756
rect 57704 521704 57756 521756
rect 302884 499536 302936 499588
rect 518164 499536 518216 499588
rect 304264 494708 304316 494760
rect 580264 494708 580316 494760
rect 49424 492124 49476 492176
rect 82176 492124 82228 492176
rect 50988 492056 51040 492108
rect 84384 492056 84436 492108
rect 140780 492056 140832 492108
rect 198924 492056 198976 492108
rect 51908 491988 51960 492040
rect 99380 491988 99432 492040
rect 109040 491988 109092 492040
rect 197452 491988 197504 492040
rect 15844 491920 15896 491972
rect 383660 491920 383712 491972
rect 214012 491512 214064 491564
rect 214932 491512 214984 491564
rect 59360 491444 59412 491496
rect 60280 491444 60332 491496
rect 204444 491444 204496 491496
rect 204812 491444 204864 491496
rect 207020 491444 207072 491496
rect 207756 491444 207808 491496
rect 209780 491444 209832 491496
rect 210516 491444 210568 491496
rect 213920 491444 213972 491496
rect 214380 491444 214432 491496
rect 215300 491444 215352 491496
rect 216220 491444 216272 491496
rect 219900 491444 219952 491496
rect 220084 491444 220136 491496
rect 64144 491240 64196 491292
rect 86224 491240 86276 491292
rect 153476 491240 153528 491292
rect 212540 491240 212592 491292
rect 213828 491240 213880 491292
rect 219256 491240 219308 491292
rect 68284 491172 68336 491224
rect 95332 491172 95384 491224
rect 150900 491172 150952 491224
rect 62856 491104 62908 491156
rect 91376 491104 91428 491156
rect 152188 491104 152240 491156
rect 72424 491036 72476 491088
rect 103336 491036 103388 491088
rect 149520 491036 149572 491088
rect 201592 491036 201644 491088
rect 50896 490968 50948 491020
rect 68928 490968 68980 491020
rect 72516 490968 72568 491020
rect 104624 490968 104676 491020
rect 157892 490968 157944 491020
rect 201684 490968 201736 491020
rect 52276 490900 52328 490952
rect 84844 490900 84896 490952
rect 149980 490900 150032 490952
rect 200764 490900 200816 490952
rect 201960 491172 202012 491224
rect 206652 491172 206704 491224
rect 211620 491172 211672 491224
rect 218152 491172 218204 491224
rect 290004 491172 290056 491224
rect 356980 491172 357032 491224
rect 248604 491104 248656 491156
rect 361120 491104 361172 491156
rect 205640 491036 205692 491088
rect 240692 491036 240744 491088
rect 356796 491036 356848 491088
rect 239404 490968 239456 491020
rect 356704 490968 356756 491020
rect 204260 490900 204312 490952
rect 238944 490900 238996 490952
rect 358268 490900 358320 490952
rect 53564 490832 53616 490884
rect 86132 490832 86184 490884
rect 156604 490832 156656 490884
rect 205640 490832 205692 490884
rect 207940 490832 207992 490884
rect 217416 490832 217468 490884
rect 237656 490832 237708 490884
rect 365168 490832 365220 490884
rect 59084 490764 59136 490816
rect 91836 490764 91888 490816
rect 155316 490764 155368 490816
rect 209044 490764 209096 490816
rect 233240 490764 233292 490816
rect 363696 490764 363748 490816
rect 55128 490696 55180 490748
rect 89168 490696 89220 490748
rect 139400 490696 139452 490748
rect 193956 490696 194008 490748
rect 194876 490696 194928 490748
rect 196808 490696 196860 490748
rect 206560 490696 206612 490748
rect 217784 490696 217836 490748
rect 225328 490696 225380 490748
rect 358176 490696 358228 490748
rect 49056 490628 49108 490680
rect 97172 490628 97224 490680
rect 138940 490628 138992 490680
rect 193864 490628 193916 490680
rect 195336 490628 195388 490680
rect 199384 490628 199436 490680
rect 201684 490628 201736 490680
rect 208400 490628 208452 490680
rect 209412 490628 209464 490680
rect 210056 490628 210108 490680
rect 223580 490628 223632 490680
rect 360936 490628 360988 490680
rect 41052 490560 41104 490612
rect 100208 490560 100260 490612
rect 110328 490560 110380 490612
rect 180064 490560 180116 490612
rect 200672 490560 200724 490612
rect 217416 490560 217468 490612
rect 223120 490560 223172 490612
rect 374644 490560 374696 490612
rect 58532 490492 58584 490544
rect 81256 490492 81308 490544
rect 157432 490492 157484 490544
rect 204260 490492 204312 490544
rect 53656 490424 53708 490476
rect 74264 490424 74316 490476
rect 154396 490424 154448 490476
rect 200580 490424 200632 490476
rect 204076 490424 204128 490476
rect 219164 490424 219216 490476
rect 56324 490356 56376 490408
rect 71780 490356 71832 490408
rect 153108 490356 153160 490408
rect 197360 490356 197412 490408
rect 68376 490288 68428 490340
rect 85212 490288 85264 490340
rect 203248 490288 203300 490340
rect 212264 490288 212316 490340
rect 67732 489948 67784 490000
rect 68192 489948 68244 490000
rect 218704 489948 218756 490000
rect 219624 489948 219676 490000
rect 50068 489880 50120 489932
rect 72240 489880 72292 489932
rect 208584 489880 208636 489932
rect 211252 489880 211304 489932
rect 283840 489336 283892 489388
rect 359740 489336 359792 489388
rect 257896 489268 257948 489320
rect 373540 489268 373592 489320
rect 167644 489200 167696 489252
rect 210516 489200 210568 489252
rect 242072 489200 242124 489252
rect 361028 489200 361080 489252
rect 59452 489132 59504 489184
rect 160744 489132 160796 489184
rect 164056 489132 164108 489184
rect 215944 489132 215996 489184
rect 222200 489132 222252 489184
rect 376024 489132 376076 489184
rect 47952 488452 48004 488504
rect 98000 488452 98052 488504
rect 59728 488384 59780 488436
rect 119620 488384 119672 488436
rect 48044 488316 48096 488368
rect 111708 488316 111760 488368
rect 46388 488248 46440 488300
rect 111248 488248 111300 488300
rect 160100 488248 160152 488300
rect 209136 488248 209188 488300
rect 50528 488180 50580 488232
rect 116032 488180 116084 488232
rect 138572 488180 138624 488232
rect 196992 488180 197044 488232
rect 46296 488112 46348 488164
rect 112076 488112 112128 488164
rect 137652 488112 137704 488164
rect 197728 488112 197780 488164
rect 48964 488044 49016 488096
rect 115204 488044 115256 488096
rect 136732 488044 136784 488096
rect 197636 488044 197688 488096
rect 46848 487976 46900 488028
rect 115664 487976 115716 488028
rect 136364 487976 136416 488028
rect 198096 487976 198148 488028
rect 59360 487908 59412 487960
rect 133144 487908 133196 487960
rect 138112 487908 138164 487960
rect 200304 487908 200356 487960
rect 256976 487908 257028 487960
rect 367928 487908 367980 487960
rect 56416 487840 56468 487892
rect 131948 487840 132000 487892
rect 135444 487840 135496 487892
rect 198188 487840 198240 487892
rect 246856 487840 246908 487892
rect 363788 487840 363840 487892
rect 48872 487772 48924 487824
rect 134616 487772 134668 487824
rect 144736 487772 144788 487824
rect 218704 487772 218756 487824
rect 236736 487772 236788 487824
rect 370504 487772 370556 487824
rect 50436 487704 50488 487756
rect 97540 487704 97592 487756
rect 51816 487636 51868 487688
rect 98460 487636 98512 487688
rect 54852 487568 54904 487620
rect 96804 487568 96856 487620
rect 177304 486548 177356 486600
rect 203708 486548 203760 486600
rect 260932 486548 260984 486600
rect 366732 486548 366784 486600
rect 164516 486480 164568 486532
rect 211804 486480 211856 486532
rect 242440 486480 242492 486532
rect 363880 486480 363932 486532
rect 144276 486412 144328 486464
rect 213276 486412 213328 486464
rect 247776 486412 247828 486464
rect 374828 486412 374880 486464
rect 57152 485732 57204 485784
rect 132408 485732 132460 485784
rect 58624 485664 58676 485716
rect 132776 485664 132828 485716
rect 44088 485596 44140 485648
rect 119160 485596 119212 485648
rect 54484 485528 54536 485580
rect 129740 485528 129792 485580
rect 57888 485460 57940 485512
rect 135904 485460 135956 485512
rect 47768 485392 47820 485444
rect 129280 485392 129332 485444
rect 47860 485324 47912 485376
rect 131028 485324 131080 485376
rect 50160 485256 50212 485308
rect 131488 485256 131540 485308
rect 44640 485188 44692 485240
rect 130200 485188 130252 485240
rect 284300 485188 284352 485240
rect 359832 485188 359884 485240
rect 44824 485120 44876 485172
rect 130568 485120 130620 485172
rect 261392 485120 261444 485172
rect 368020 485120 368072 485172
rect 46204 485052 46256 485104
rect 133236 485052 133288 485104
rect 159640 485052 159692 485104
rect 214564 485052 214616 485104
rect 242900 485052 242952 485104
rect 369124 485052 369176 485104
rect 46756 484984 46808 485036
rect 116952 484984 117004 485036
rect 48228 484916 48280 484968
rect 117872 484916 117924 484968
rect 58808 484848 58860 484900
rect 110788 484848 110840 484900
rect 292212 484304 292264 484356
rect 368204 484304 368256 484356
rect 270224 484236 270276 484288
rect 357072 484236 357124 484288
rect 269764 484168 269816 484220
rect 358728 484168 358780 484220
rect 280804 484100 280856 484152
rect 374460 484100 374512 484152
rect 281264 484032 281316 484084
rect 376576 484032 376628 484084
rect 268936 483964 268988 484016
rect 370964 483964 371016 484016
rect 268476 483896 268528 483948
rect 377312 483896 377364 483948
rect 260564 483828 260616 483880
rect 369400 483828 369452 483880
rect 243360 483760 243412 483812
rect 366548 483760 366600 483812
rect 205456 483692 205508 483744
rect 217324 483692 217376 483744
rect 231860 483692 231912 483744
rect 366456 483692 366508 483744
rect 58716 483624 58768 483676
rect 96252 483624 96304 483676
rect 184296 483624 184348 483676
rect 214840 483624 214892 483676
rect 238484 483624 238536 483676
rect 378784 483624 378836 483676
rect 57704 482944 57756 482996
rect 114284 482944 114336 482996
rect 59636 482876 59688 482928
rect 127992 482876 128044 482928
rect 58440 482808 58492 482860
rect 128820 482808 128872 482860
rect 50344 482740 50396 482792
rect 126244 482740 126296 482792
rect 43628 482672 43680 482724
rect 123576 482672 123628 482724
rect 43812 482604 43864 482656
rect 124404 482604 124456 482656
rect 43904 482536 43956 482588
rect 124864 482536 124916 482588
rect 43720 482468 43772 482520
rect 125784 482468 125836 482520
rect 40960 482400 41012 482452
rect 123116 482400 123168 482452
rect 253020 482400 253072 482452
rect 375012 482400 375064 482452
rect 48780 482332 48832 482384
rect 133696 482332 133748 482384
rect 245108 482332 245160 482384
rect 370596 482332 370648 482384
rect 43260 482264 43312 482316
rect 143816 482264 143868 482316
rect 171968 482264 172020 482316
rect 203524 482264 203576 482316
rect 239864 482264 239916 482316
rect 378876 482264 378928 482316
rect 292672 481448 292724 481500
rect 357992 481448 358044 481500
rect 291844 481380 291896 481432
rect 365628 481380 365680 481432
rect 289636 481312 289688 481364
rect 368388 481312 368440 481364
rect 279056 481244 279108 481296
rect 360844 481244 360896 481296
rect 279516 481176 279568 481228
rect 364156 481176 364208 481228
rect 279884 481108 279936 481160
rect 367008 481108 367060 481160
rect 274640 481040 274692 481092
rect 364892 481040 364944 481092
rect 177764 480972 177816 481024
rect 202328 480972 202380 481024
rect 275100 480972 275152 481024
rect 367652 480972 367704 481024
rect 162308 480904 162360 480956
rect 204904 480904 204956 480956
rect 258816 480904 258868 480956
rect 365444 480904 365496 480956
rect 254400 479680 254452 479732
rect 373632 479680 373684 479732
rect 176384 479612 176436 479664
rect 209504 479612 209556 479664
rect 238116 479612 238168 479664
rect 376116 479612 376168 479664
rect 166264 479544 166316 479596
rect 213368 479544 213420 479596
rect 227904 479544 227956 479596
rect 367744 479544 367796 479596
rect 3516 479476 3568 479528
rect 309784 479476 309836 479528
rect 291384 478796 291436 478848
rect 362684 478796 362736 478848
rect 289176 478728 289228 478780
rect 360752 478728 360804 478780
rect 278596 478660 278648 478712
rect 357164 478660 357216 478712
rect 278136 478592 278188 478644
rect 362776 478592 362828 478644
rect 273720 478524 273772 478576
rect 360660 478524 360712 478576
rect 273260 478456 273312 478508
rect 364248 478456 364300 478508
rect 256148 478388 256200 478440
rect 356888 478388 356940 478440
rect 256608 478320 256660 478372
rect 358452 478320 358504 478372
rect 260104 478252 260156 478304
rect 362500 478252 362552 478304
rect 159272 478184 159324 478236
rect 204996 478184 205048 478236
rect 246028 478184 246080 478236
rect 369216 478184 369268 478236
rect 3608 478116 3660 478168
rect 434812 478116 434864 478168
rect 178592 476892 178644 476944
rect 200856 476892 200908 476944
rect 259644 476892 259696 476944
rect 370872 476892 370924 476944
rect 163228 476824 163280 476876
rect 210608 476824 210660 476876
rect 244648 476824 244700 476876
rect 371884 476824 371936 476876
rect 62764 476756 62816 476808
rect 199108 476756 199160 476808
rect 232780 476756 232832 476808
rect 364984 476756 365036 476808
rect 290924 475804 290976 475856
rect 361396 475804 361448 475856
rect 285680 475736 285732 475788
rect 358084 475736 358136 475788
rect 277676 475668 277728 475720
rect 364800 475668 364852 475720
rect 266268 475600 266320 475652
rect 358544 475600 358596 475652
rect 272892 475532 272944 475584
rect 366272 475532 366324 475584
rect 170680 475464 170732 475516
rect 211896 475464 211948 475516
rect 253940 475464 253992 475516
rect 361212 475464 361264 475516
rect 148232 475396 148284 475448
rect 213184 475396 213236 475448
rect 265348 475396 265400 475448
rect 376300 475396 376352 475448
rect 61936 475328 61988 475380
rect 199200 475328 199252 475380
rect 245568 475328 245620 475380
rect 362316 475328 362368 475380
rect 43352 474648 43404 474700
rect 72516 474648 72568 474700
rect 51724 474580 51776 474632
rect 99748 474580 99800 474632
rect 50252 474512 50304 474564
rect 98920 474512 98972 474564
rect 51632 474444 51684 474496
rect 100668 474444 100720 474496
rect 45192 474376 45244 474428
rect 105084 474376 105136 474428
rect 45100 474308 45152 474360
rect 105912 474308 105964 474360
rect 43536 474240 43588 474292
rect 103704 474240 103756 474292
rect 193956 474240 194008 474292
rect 205732 474240 205784 474292
rect 45008 474172 45060 474224
rect 105544 474172 105596 474224
rect 186136 474172 186188 474224
rect 213552 474172 213604 474224
rect 287796 474172 287848 474224
rect 369032 474172 369084 474224
rect 45376 474104 45428 474156
rect 106372 474104 106424 474156
rect 139860 474104 139912 474156
rect 207296 474104 207348 474156
rect 259184 474104 259236 474156
rect 372068 474104 372120 474156
rect 45284 474036 45336 474088
rect 106832 474036 106884 474088
rect 127532 474036 127584 474088
rect 204352 474036 204404 474088
rect 237196 474036 237248 474088
rect 362408 474036 362460 474088
rect 61476 473968 61528 474020
rect 199476 473968 199528 474020
rect 248236 473968 248288 474020
rect 376208 473968 376260 474020
rect 43444 473900 43496 473952
rect 72424 473900 72476 473952
rect 264060 473220 264112 473272
rect 362592 473220 362644 473272
rect 264520 473152 264572 473204
rect 363972 473152 364024 473204
rect 265808 473084 265860 473136
rect 365536 473084 365588 473136
rect 267556 473016 267608 473068
rect 375196 473016 375248 473068
rect 264980 472948 265032 473000
rect 373724 472948 373776 473000
rect 261852 472880 261904 472932
rect 376392 472880 376444 472932
rect 187424 472812 187476 472864
rect 207756 472812 207808 472864
rect 241612 472812 241664 472864
rect 370688 472812 370740 472864
rect 176016 472744 176068 472796
rect 205088 472744 205140 472796
rect 205916 472744 205968 472796
rect 217692 472744 217744 472796
rect 227076 472744 227128 472796
rect 362224 472744 362276 472796
rect 176844 472676 176896 472728
rect 210700 472676 210752 472728
rect 222660 472676 222712 472728
rect 365076 472676 365128 472728
rect 57612 472608 57664 472660
rect 113916 472608 113968 472660
rect 161020 472608 161072 472660
rect 206284 472608 206336 472660
rect 227536 472608 227588 472660
rect 374736 472608 374788 472660
rect 50988 471928 51040 471980
rect 83004 471928 83056 471980
rect 193128 471928 193180 471980
rect 214932 471928 214984 471980
rect 53472 471860 53524 471912
rect 85672 471860 85724 471912
rect 190920 471860 190972 471912
rect 215852 471860 215904 471912
rect 299756 471860 299808 471912
rect 373080 471860 373132 471912
rect 56324 471792 56376 471844
rect 90088 471792 90140 471844
rect 183008 471792 183060 471844
rect 216128 471792 216180 471844
rect 294880 471792 294932 471844
rect 372436 471792 372488 471844
rect 49332 471724 49384 471776
rect 83464 471724 83516 471776
rect 175096 471724 175148 471776
rect 212080 471724 212132 471776
rect 286048 471724 286100 471776
rect 366180 471724 366232 471776
rect 58900 471656 58952 471708
rect 95792 471656 95844 471708
rect 179052 471656 179104 471708
rect 216772 471656 216824 471708
rect 293592 471656 293644 471708
rect 375932 471656 375984 471708
rect 56876 471588 56928 471640
rect 102876 471588 102928 471640
rect 140320 471588 140372 471640
rect 196900 471588 196952 471640
rect 287428 471588 287480 471640
rect 370412 471588 370464 471640
rect 54668 471520 54720 471572
rect 102416 471520 102468 471572
rect 141148 471520 141200 471572
rect 200396 471520 200448 471572
rect 286508 471520 286560 471572
rect 369768 471520 369820 471572
rect 53196 471452 53248 471504
rect 101128 471452 101180 471504
rect 141608 471452 141660 471504
rect 204628 471452 204680 471504
rect 286968 471452 287020 471504
rect 375288 471452 375340 471504
rect 52828 471384 52880 471436
rect 101496 471384 101548 471436
rect 142068 471384 142120 471436
rect 205824 471384 205876 471436
rect 282552 471384 282604 471436
rect 374552 471384 374604 471436
rect 56692 471316 56744 471368
rect 114744 471316 114796 471368
rect 127072 471316 127124 471368
rect 202880 471316 202932 471368
rect 271512 471316 271564 471368
rect 371792 471316 371844 471368
rect 42616 471248 42668 471300
rect 104164 471248 104216 471300
rect 109500 471248 109552 471300
rect 202972 471248 203024 471300
rect 271144 471248 271196 471300
rect 373172 471248 373224 471300
rect 52092 471180 52144 471232
rect 83924 471180 83976 471232
rect 191380 471180 191432 471232
rect 210240 471180 210292 471232
rect 44732 471112 44784 471164
rect 65432 471112 65484 471164
rect 188712 471112 188764 471164
rect 200764 471112 200816 471164
rect 47676 471044 47728 471096
rect 64972 471044 65024 471096
rect 193864 470568 193916 470620
rect 201868 470568 201920 470620
rect 283472 470500 283524 470552
rect 360016 470500 360068 470552
rect 283012 470432 283064 470484
rect 359924 470432 359976 470484
rect 281632 470364 281684 470416
rect 359648 470364 359700 470416
rect 298008 470296 298060 470348
rect 378232 470296 378284 470348
rect 293132 470228 293184 470280
rect 376760 470228 376812 470280
rect 293960 470160 294012 470212
rect 379244 470160 379296 470212
rect 284760 470092 284812 470144
rect 377404 470092 377456 470144
rect 175556 470024 175608 470076
rect 210792 470024 210844 470076
rect 282092 470024 282144 470076
rect 379980 470024 380032 470076
rect 173808 469956 173860 470008
rect 209412 469956 209464 470008
rect 250812 469956 250864 470008
rect 365260 469956 365312 470008
rect 178132 469888 178184 469940
rect 215208 469888 215260 469940
rect 251272 469888 251324 469940
rect 373356 469888 373408 469940
rect 57520 469820 57572 469872
rect 112996 469820 113048 469872
rect 161480 469820 161532 469872
rect 207664 469820 207716 469872
rect 240232 469820 240284 469872
rect 366640 469820 366692 469872
rect 295800 469752 295852 469804
rect 357256 469752 357308 469804
rect 56048 469140 56100 469192
rect 81716 469140 81768 469192
rect 186504 469140 186556 469192
rect 206468 469140 206520 469192
rect 269304 469140 269356 469192
rect 359464 469140 359516 469192
rect 56140 469072 56192 469124
rect 87880 469072 87932 469124
rect 181720 469072 181772 469124
rect 203800 469072 203852 469124
rect 277308 469072 277360 469124
rect 367560 469072 367612 469124
rect 55036 469004 55088 469056
rect 87052 469004 87104 469056
rect 192668 469004 192720 469056
rect 217968 469004 218020 469056
rect 266728 469004 266780 469056
rect 358636 469004 358688 469056
rect 55956 468936 56008 468988
rect 88800 468936 88852 468988
rect 190460 468936 190512 468988
rect 217508 468936 217560 468988
rect 267096 468936 267148 468988
rect 359556 468936 359608 468988
rect 55864 468868 55916 468920
rect 89628 468868 89680 468920
rect 189632 468868 189684 468920
rect 217600 468868 217652 468920
rect 285220 468868 285272 468920
rect 377772 468868 377824 468920
rect 54944 468800 54996 468852
rect 88340 468800 88392 468852
rect 168472 468800 168524 468852
rect 209320 468800 209372 468852
rect 275468 468800 275520 468852
rect 370320 468800 370372 468852
rect 52000 468732 52052 468784
rect 86592 468732 86644 468784
rect 169392 468732 169444 468784
rect 211988 468732 212040 468784
rect 272432 468732 272484 468784
rect 368848 468732 368900 468784
rect 57336 468664 57388 468716
rect 113456 468664 113508 468716
rect 170220 468664 170272 468716
rect 213460 468664 213512 468716
rect 271972 468664 272024 468716
rect 372252 468664 372304 468716
rect 53380 468596 53432 468648
rect 87420 468596 87472 468648
rect 109868 468596 109920 468648
rect 197452 468596 197504 468648
rect 268016 468596 268068 468648
rect 377220 468596 377272 468648
rect 53288 468528 53340 468580
rect 94044 468528 94096 468580
rect 108120 468528 108172 468580
rect 200120 468528 200172 468580
rect 255228 468528 255280 468580
rect 366824 468528 366876 468580
rect 49240 468460 49292 468512
rect 94504 468460 94556 468512
rect 108580 468460 108632 468512
rect 201684 468460 201736 468512
rect 254768 468460 254820 468512
rect 375104 468460 375156 468512
rect 49976 468392 50028 468444
rect 68376 468392 68428 468444
rect 193588 468392 193640 468444
rect 213092 468392 213144 468444
rect 298836 468392 298888 468444
rect 378140 468392 378192 468444
rect 46112 468324 46164 468376
rect 64512 468324 64564 468376
rect 183928 468324 183980 468376
rect 200948 468324 201000 468376
rect 290464 468324 290516 468376
rect 363512 468324 363564 468376
rect 60004 468256 60056 468308
rect 67732 468256 67784 468308
rect 197268 468256 197320 468308
rect 209780 468256 209832 468308
rect 133144 467780 133196 467832
rect 178040 467780 178092 467832
rect 296628 467780 296680 467832
rect 360568 467780 360620 467832
rect 160744 467712 160796 467764
rect 179420 467712 179472 467764
rect 299296 467712 299348 467764
rect 371240 467712 371292 467764
rect 288256 467644 288308 467696
rect 375840 467644 375892 467696
rect 262312 467576 262364 467628
rect 364064 467576 364116 467628
rect 42524 467508 42576 467560
rect 61016 467508 61068 467560
rect 270684 467508 270736 467560
rect 377128 467508 377180 467560
rect 40868 467440 40920 467492
rect 62304 467440 62356 467492
rect 190092 467440 190144 467492
rect 208032 467440 208084 467492
rect 252192 467440 252244 467492
rect 361304 467440 361356 467492
rect 41144 467372 41196 467424
rect 68284 467372 68336 467424
rect 185216 467372 185268 467424
rect 212172 467372 212224 467424
rect 251732 467372 251784 467424
rect 365352 467372 365404 467424
rect 41236 467304 41288 467356
rect 72884 467304 72936 467356
rect 182180 467304 182232 467356
rect 209596 467304 209648 467356
rect 249524 467304 249576 467356
rect 367836 467304 367888 467356
rect 42708 467236 42760 467288
rect 94964 467236 95016 467288
rect 188344 467236 188396 467288
rect 216220 467236 216272 467288
rect 249984 467236 250036 467288
rect 369308 467236 369360 467288
rect 57428 467168 57480 467220
rect 112536 467168 112588 467220
rect 171600 467168 171652 467220
rect 214748 467168 214800 467220
rect 250444 467168 250496 467220
rect 371976 467168 372028 467220
rect 44916 467100 44968 467152
rect 107292 467100 107344 467152
rect 165436 467100 165488 467152
rect 218888 467100 218940 467152
rect 249064 467100 249116 467152
rect 370780 467100 370832 467152
rect 59268 467032 59320 467084
rect 67180 467032 67232 467084
rect 178040 466556 178092 466608
rect 204536 466556 204588 466608
rect 338488 466556 338540 466608
rect 361580 466556 361632 466608
rect 498476 466624 498528 466676
rect 499488 466624 499540 466676
rect 179420 466488 179472 466540
rect 201776 466488 201828 466540
rect 339776 466488 339828 466540
rect 362960 466488 363012 466540
rect 190920 466420 190972 466472
rect 210424 466420 210476 466472
rect 351000 466420 351052 466472
rect 358820 466420 358872 466472
rect 499764 466556 499816 466608
rect 517888 466556 517940 466608
rect 499488 466488 499540 466540
rect 510896 466488 510948 466540
rect 517520 466488 517572 466540
rect 517796 466420 517848 466472
rect 50712 466352 50764 466404
rect 79508 466352 79560 466404
rect 194048 466352 194100 466404
rect 212908 466352 212960 466404
rect 213828 466352 213880 466404
rect 221372 466352 221424 466404
rect 280344 466352 280396 466404
rect 368940 466352 368992 466404
rect 180340 466284 180392 466336
rect 207848 466284 207900 466336
rect 275928 466284 275980 466336
rect 372988 466284 373040 466336
rect 174176 466216 174228 466268
rect 203892 466216 203944 466268
rect 263140 466216 263192 466268
rect 369492 466216 369544 466268
rect 54392 466148 54444 466200
rect 63224 466148 63276 466200
rect 168012 466148 168064 466200
rect 203616 466148 203668 466200
rect 263600 466148 263652 466200
rect 372160 466148 372212 466200
rect 59176 466080 59228 466132
rect 67640 466080 67692 466132
rect 179512 466080 179564 466132
rect 216312 466080 216364 466132
rect 257436 466080 257488 466132
rect 366916 466080 366968 466132
rect 54300 466012 54352 466064
rect 63684 466012 63736 466064
rect 166724 466012 166776 466064
rect 206376 466012 206428 466064
rect 258356 466012 258408 466064
rect 368112 466012 368164 466064
rect 51540 465944 51592 465996
rect 66720 465944 66772 465996
rect 174636 465944 174688 465996
rect 219164 465944 219216 465996
rect 243820 465944 243872 465996
rect 358360 465944 358412 465996
rect 55588 465876 55640 465928
rect 75552 465876 75604 465928
rect 164976 465876 165028 465928
rect 214656 465876 214708 465928
rect 262772 465876 262824 465928
rect 379060 465876 379112 465928
rect 49516 465808 49568 465860
rect 71136 465808 71188 465860
rect 143356 465808 143408 465860
rect 200488 465808 200540 465860
rect 244280 465808 244332 465860
rect 373448 465808 373500 465860
rect 50804 465740 50856 465792
rect 50988 465740 51040 465792
rect 50620 465672 50672 465724
rect 93584 465740 93636 465792
rect 142528 465740 142580 465792
rect 207112 465740 207164 465792
rect 212448 465740 212500 465792
rect 221740 465740 221792 465792
rect 246396 465740 246448 465792
rect 378968 465740 379020 465792
rect 49608 465604 49660 465656
rect 71780 465672 71832 465724
rect 86224 465672 86276 465724
rect 198740 465672 198792 465724
rect 205548 465672 205600 465724
rect 220912 465672 220964 465724
rect 241152 465672 241204 465724
rect 374920 465672 374972 465724
rect 59820 465604 59872 465656
rect 62856 465604 62908 465656
rect 187884 465604 187936 465656
rect 202512 465604 202564 465656
rect 274180 465604 274232 465656
rect 362132 465604 362184 465656
rect 189172 465536 189224 465588
rect 202144 465536 202196 465588
rect 297088 465536 297140 465588
rect 362868 465536 362920 465588
rect 195796 465468 195848 465520
rect 206744 465468 206796 465520
rect 198740 465060 198792 465112
rect 358912 465060 358964 465112
rect 518900 465060 518952 465112
rect 196992 464992 197044 465044
rect 200580 464992 200632 465044
rect 58992 464720 59044 464772
rect 93216 464720 93268 464772
rect 192300 464720 192352 464772
rect 208952 464720 209004 464772
rect 49976 464652 50028 464704
rect 50712 464652 50764 464704
rect 53012 464652 53064 464704
rect 101956 464652 102008 464704
rect 191840 464652 191892 464704
rect 211620 464652 211672 464704
rect 55772 464584 55824 464636
rect 122656 464584 122708 464636
rect 194508 464584 194560 464636
rect 214472 464584 214524 464636
rect 54576 464516 54628 464568
rect 121828 464516 121880 464568
rect 180800 464516 180852 464568
rect 210884 464516 210936 464568
rect 57060 464448 57112 464500
rect 134984 464448 135036 464500
rect 142896 464448 142948 464500
rect 197820 464448 197872 464500
rect 52184 464380 52236 464432
rect 134156 464380 134208 464432
rect 137192 464380 137244 464432
rect 199016 464380 199068 464432
rect 47584 464312 47636 464364
rect 207388 464448 207440 464500
rect 208216 464448 208268 464500
rect 294420 464448 294472 464500
rect 370228 464448 370280 464500
rect 288716 464380 288768 464432
rect 367468 464380 367520 464432
rect 207480 464312 207532 464364
rect 208124 464312 208176 464364
rect 276848 464312 276900 464364
rect 357900 464312 357952 464364
rect 46020 464244 46072 464296
rect 208216 418752 208268 418804
rect 216864 418752 216916 418804
rect 46020 418072 46072 418124
rect 57796 418072 57848 418124
rect 47584 418004 47636 418056
rect 57244 418004 57296 418056
rect 203064 418004 203116 418056
rect 208216 418004 208268 418056
rect 208124 417392 208176 417444
rect 216772 417392 216824 417444
rect 358084 417392 358136 417444
rect 377036 417392 377088 417444
rect 377588 417392 377640 417444
rect 206836 416712 206888 416764
rect 207204 416712 207256 416764
rect 198188 416032 198240 416084
rect 203064 416032 203116 416084
rect 207204 414808 207256 414860
rect 216864 414808 216916 414860
rect 206192 414672 206244 414724
rect 216956 414672 217008 414724
rect 47492 413992 47544 414044
rect 57796 413992 57848 414044
rect 206008 413244 206060 413296
rect 216680 413244 216732 413296
rect 359832 413244 359884 413296
rect 377680 413244 377732 413296
rect 47400 412632 47452 412684
rect 57796 412632 57848 412684
rect 359740 411884 359792 411936
rect 377036 411884 377088 411936
rect 204444 411476 204496 411528
rect 206836 411476 206888 411528
rect 47584 411272 47636 411324
rect 57796 411272 57848 411324
rect 2964 411204 3016 411256
rect 15844 411204 15896 411256
rect 51632 410592 51684 410644
rect 52920 410592 52972 410644
rect 198096 410524 198148 410576
rect 204444 410524 204496 410576
rect 360016 410524 360068 410576
rect 377404 410524 377456 410576
rect 377864 410524 377916 410576
rect 51632 409844 51684 409896
rect 57796 409844 57848 409896
rect 217968 409844 218020 409896
rect 218612 409844 218664 409896
rect 206836 409096 206888 409148
rect 216772 409096 216824 409148
rect 216956 409096 217008 409148
rect 359924 409096 359976 409148
rect 377404 409096 377456 409148
rect 52368 408484 52420 408536
rect 57796 408484 57848 408536
rect 216680 407600 216732 407652
rect 216772 407396 216824 407448
rect 520924 405628 520976 405680
rect 580172 405628 580224 405680
rect 199016 400528 199068 400580
rect 199108 400528 199160 400580
rect 199844 400528 199896 400580
rect 199016 400324 199068 400376
rect 198924 400188 198976 400240
rect 208492 400188 208544 400240
rect 378140 398080 378192 398132
rect 378324 398080 378376 398132
rect 198096 397400 198148 397452
rect 199108 397400 199160 397452
rect 56508 391960 56560 392012
rect 57060 391960 57112 392012
rect 43260 391892 43312 391944
rect 57704 391892 57756 391944
rect 208216 391892 208268 391944
rect 216956 391892 217008 391944
rect 359648 391892 359700 391944
rect 376852 391892 376904 391944
rect 57152 390532 57204 390584
rect 58440 390532 58492 390584
rect 358820 390464 358872 390516
rect 376944 390464 376996 390516
rect 210424 389308 210476 389360
rect 216680 389308 216732 389360
rect 52460 389172 52512 389224
rect 53748 389172 53800 389224
rect 57428 389172 57480 389224
rect 358084 389172 358136 389224
rect 358820 389172 358872 389224
rect 47768 389104 47820 389156
rect 57244 389104 57296 389156
rect 202144 389104 202196 389156
rect 216956 389104 217008 389156
rect 359556 389104 359608 389156
rect 376944 389104 376996 389156
rect 56784 388492 56836 388544
rect 58532 388492 58584 388544
rect 45468 388424 45520 388476
rect 52460 388424 52512 388476
rect 57060 388424 57112 388476
rect 58440 388424 58492 388476
rect 57152 387948 57204 388000
rect 57796 387948 57848 388000
rect 378140 383936 378192 383988
rect 378324 383936 378376 383988
rect 199292 382916 199344 382968
rect 219808 382916 219860 382968
rect 57796 382032 57848 382084
rect 59360 382032 59412 382084
rect 195060 380944 195112 380996
rect 200580 380944 200632 380996
rect 55772 380876 55824 380928
rect 57060 380876 57112 380928
rect 58348 380876 58400 380928
rect 60740 380876 60792 380928
rect 194600 380876 194652 380928
rect 197728 380876 197780 380928
rect 217600 380876 217652 380928
rect 248236 380876 248288 380928
rect 358728 380876 358780 380928
rect 421104 380876 421156 380928
rect 47400 380808 47452 380860
rect 216772 380808 216824 380860
rect 47492 380740 47544 380792
rect 216680 380740 216732 380792
rect 356980 380740 357032 380792
rect 380992 380740 381044 380792
rect 51632 380672 51684 380724
rect 217140 380672 217192 380724
rect 377312 380672 377364 380724
rect 413560 380672 413612 380724
rect 52368 380604 52420 380656
rect 216864 380604 216916 380656
rect 357992 380604 358044 380656
rect 376484 380604 376536 380656
rect 377128 380604 377180 380656
rect 425980 380604 426032 380656
rect 155960 380536 156012 380588
rect 204628 380536 204680 380588
rect 360568 380536 360620 380588
rect 369584 380536 369636 380588
rect 372252 380536 372304 380588
rect 433616 380536 433668 380588
rect 143632 380468 143684 380520
rect 205732 380468 205784 380520
rect 368848 380468 368900 380520
rect 436008 380468 436060 380520
rect 56508 380400 56560 380452
rect 118332 380400 118384 380452
rect 121000 380400 121052 380452
rect 203064 380400 203116 380452
rect 366272 380400 366324 380452
rect 438492 380400 438544 380452
rect 52184 380332 52236 380384
rect 113548 380332 113600 380384
rect 163504 380332 163556 380384
rect 197820 380332 197872 380384
rect 201592 380332 201644 380384
rect 291844 380332 291896 380384
rect 364248 380332 364300 380384
rect 440884 380332 440936 380384
rect 48780 380264 48832 380316
rect 110972 380264 111024 380316
rect 148600 380264 148652 380316
rect 196900 380264 196952 380316
rect 199752 380264 199804 380316
rect 298008 380264 298060 380316
rect 364892 380264 364944 380316
rect 448244 380264 448296 380316
rect 57888 380196 57940 380248
rect 123484 380196 123536 380248
rect 135904 380196 135956 380248
rect 200304 380196 200356 380248
rect 201040 380196 201092 380248
rect 313464 380196 313516 380248
rect 360660 380196 360712 380248
rect 443460 380196 443512 380248
rect 48872 380128 48924 380180
rect 115940 380128 115992 380180
rect 128360 380128 128412 380180
rect 197636 380128 197688 380180
rect 201500 380128 201552 380180
rect 315856 380128 315908 380180
rect 362132 380128 362184 380180
rect 445944 380128 445996 380180
rect 158536 380060 158588 380112
rect 205824 380060 205876 380112
rect 160928 379992 160980 380044
rect 207112 379992 207164 380044
rect 213736 379992 213788 380044
rect 236000 379992 236052 380044
rect 166080 379924 166132 379976
rect 200488 379924 200540 379976
rect 215300 379924 215352 379976
rect 216404 379924 216456 379976
rect 243084 379924 243136 379976
rect 208308 379856 208360 379908
rect 237104 379856 237156 379908
rect 239772 379856 239824 379908
rect 261760 379856 261812 379908
rect 213644 379788 213696 379840
rect 214104 379788 214156 379840
rect 244280 379788 244332 379840
rect 375288 379788 375340 379840
rect 405464 379788 405516 379840
rect 212632 379720 212684 379772
rect 219716 379720 219768 379772
rect 254492 379720 254544 379772
rect 380992 379720 381044 379772
rect 413468 379720 413520 379772
rect 215668 379652 215720 379704
rect 216036 379652 216088 379704
rect 217324 379652 217376 379704
rect 216680 379584 216732 379636
rect 217600 379584 217652 379636
rect 204168 379516 204220 379568
rect 213736 379516 213788 379568
rect 216864 379516 216916 379568
rect 217324 379516 217376 379568
rect 217968 379652 218020 379704
rect 255872 379652 255924 379704
rect 369768 379652 369820 379704
rect 371148 379652 371200 379704
rect 404176 379652 404228 379704
rect 219256 379584 219308 379636
rect 219440 379584 219492 379636
rect 258080 379584 258132 379636
rect 369584 379584 369636 379636
rect 263876 379516 263928 379568
rect 54484 379448 54536 379500
rect 88340 379448 88392 379500
rect 92388 379448 92440 379500
rect 86592 379380 86644 379432
rect 210056 379380 210108 379432
rect 211528 379380 211580 379432
rect 85488 379312 85540 379364
rect 208768 379312 208820 379364
rect 88800 379244 88852 379296
rect 210332 379244 210384 379296
rect 210976 379244 211028 379296
rect 213736 379380 213788 379432
rect 219532 379448 219584 379500
rect 273260 379448 273312 379500
rect 291844 379448 291896 379500
rect 320916 379448 320968 379500
rect 369676 379516 369728 379568
rect 371240 379516 371292 379568
rect 376484 379584 376536 379636
rect 376668 379584 376720 379636
rect 420644 379584 420696 379636
rect 369768 379448 369820 379500
rect 431132 379516 431184 379568
rect 437940 379448 437992 379500
rect 218244 379380 218296 379432
rect 269764 379380 269816 379432
rect 298008 379380 298060 379432
rect 305828 379380 305880 379432
rect 378232 379380 378284 379432
rect 434260 379380 434312 379432
rect 220452 379312 220504 379364
rect 271052 379312 271104 379364
rect 375196 379312 375248 379364
rect 408316 379312 408368 379364
rect 218152 379244 218204 379296
rect 221004 379244 221056 379296
rect 222016 379244 222068 379296
rect 91376 379176 91428 379228
rect 44640 379108 44692 379160
rect 90732 379108 90784 379160
rect 90824 379108 90876 379160
rect 195980 379108 196032 379160
rect 211160 379108 211212 379160
rect 221464 379108 221516 379160
rect 44824 379040 44876 379092
rect 93492 379040 93544 379092
rect 93584 379040 93636 379092
rect 198648 379040 198700 379092
rect 220820 379040 220872 379092
rect 222108 379040 222160 379092
rect 46204 378972 46256 379024
rect 108212 378972 108264 379024
rect 115848 378972 115900 379024
rect 219900 378972 219952 379024
rect 220728 378972 220780 379024
rect 58624 378904 58676 378956
rect 105360 378904 105412 378956
rect 112352 378904 112404 378956
rect 204076 378904 204128 378956
rect 211712 378904 211764 378956
rect 368388 378904 368440 378956
rect 379612 378904 379664 378956
rect 379980 378904 380032 378956
rect 396080 378904 396132 378956
rect 58440 378836 58492 378888
rect 103520 378836 103572 378888
rect 117136 378836 117188 378888
rect 205548 378836 205600 378888
rect 213828 378836 213880 378888
rect 214104 378836 214156 378888
rect 266452 378836 266504 378888
rect 268292 378836 268344 378888
rect 360752 378836 360804 378888
rect 379520 378836 379572 378888
rect 56416 378768 56468 378820
rect 101036 378768 101088 378820
rect 195980 378768 196032 378820
rect 197268 378768 197320 378820
rect 77208 378700 77260 378752
rect 99380 378700 99432 378752
rect 211528 378700 211580 378752
rect 218336 378700 218388 378752
rect 220636 378768 220688 378820
rect 248604 378768 248656 378820
rect 374552 378768 374604 378820
rect 396356 378768 396408 378820
rect 219532 378700 219584 378752
rect 250076 378700 250128 378752
rect 343548 378700 343600 378752
rect 503628 378700 503680 378752
rect 50160 378632 50212 378684
rect 98460 378632 98512 378684
rect 210976 378632 211028 378684
rect 219992 378632 220044 378684
rect 220636 378632 220688 378684
rect 221096 378632 221148 378684
rect 221464 378632 221516 378684
rect 251180 378632 251232 378684
rect 369584 378632 369636 378684
rect 398196 378632 398248 378684
rect 47860 378564 47912 378616
rect 96068 378564 96120 378616
rect 205640 378564 205692 378616
rect 206836 378564 206888 378616
rect 219624 378564 219676 378616
rect 220452 378564 220504 378616
rect 222016 378564 222068 378616
rect 252284 378564 252336 378616
rect 342904 378564 342956 378616
rect 343456 378564 343508 378616
rect 358820 378564 358872 378616
rect 359280 378564 359332 378616
rect 370412 378564 370464 378616
rect 376484 378564 376536 378616
rect 405832 378564 405884 378616
rect 113456 378496 113508 378548
rect 213000 378496 213052 378548
rect 213736 378496 213788 378548
rect 222108 378496 222160 378548
rect 253388 378496 253440 378548
rect 262220 378496 262272 378548
rect 266360 378496 266412 378548
rect 280068 378496 280120 378548
rect 360016 378496 360068 378548
rect 208768 378428 208820 378480
rect 212356 378428 212408 378480
rect 244924 378428 244976 378480
rect 276020 378428 276072 378480
rect 277032 378428 277084 378480
rect 356980 378428 357032 378480
rect 114468 378360 114520 378412
rect 207020 378360 207072 378412
rect 207572 378360 207624 378412
rect 210332 378360 210384 378412
rect 239588 378360 239640 378412
rect 368296 378496 368348 378548
rect 399484 378496 399536 378548
rect 379612 378428 379664 378480
rect 412364 378428 412416 378480
rect 369032 378360 369084 378412
rect 373816 378360 373868 378412
rect 111248 378292 111300 378344
rect 205640 378292 205692 378344
rect 205732 378292 205784 378344
rect 206928 378292 206980 378344
rect 238208 378292 238260 378344
rect 369584 378292 369636 378344
rect 379520 378360 379572 378412
rect 411260 378360 411312 378412
rect 511908 378360 511960 378412
rect 517520 378360 517572 378412
rect 407580 378292 407632 378344
rect 204812 378224 204864 378276
rect 210976 378224 211028 378276
rect 44732 378156 44784 378208
rect 47768 378156 47820 378208
rect 80428 378156 80480 378208
rect 109776 378156 109828 378208
rect 218244 378224 218296 378276
rect 218336 378224 218388 378276
rect 246212 378224 246264 378276
rect 263876 378224 263928 378276
rect 267556 378224 267608 378276
rect 274640 378224 274692 378276
rect 275744 378224 275796 378276
rect 356612 378224 356664 378276
rect 359280 378224 359332 378276
rect 40868 378020 40920 378072
rect 198924 378088 198976 378140
rect 199660 378088 199712 378140
rect 211712 378156 211764 378208
rect 272156 378156 272208 378208
rect 273260 378156 273312 378208
rect 285956 378156 286008 378208
rect 503628 378224 503680 378276
rect 517612 378224 517664 378276
rect 580264 378224 580316 378276
rect 503352 378156 503404 378208
rect 517704 378156 517756 378208
rect 580172 378156 580224 378208
rect 217416 378088 217468 378140
rect 310980 378088 311032 378140
rect 360844 378088 360896 378140
rect 473452 378088 473504 378140
rect 205364 378020 205416 378072
rect 206192 378020 206244 378072
rect 210976 378020 211028 378072
rect 212264 378020 212316 378072
rect 325884 378020 325936 378072
rect 368940 378020 368992 378072
rect 480628 378020 480680 378072
rect 54300 377952 54352 378004
rect 182364 377952 182416 378004
rect 182916 377952 182968 378004
rect 205456 377952 205508 378004
rect 206560 377952 206612 378004
rect 206652 377952 206704 378004
rect 317788 377952 317840 378004
rect 376576 377952 376628 378004
rect 485964 377952 486016 378004
rect 54392 377884 54444 377936
rect 182272 377884 182324 377936
rect 200212 377884 200264 377936
rect 307852 377884 307904 377936
rect 357900 377884 357952 377936
rect 460940 377884 460992 377936
rect 196624 377816 196676 377868
rect 273260 377816 273312 377868
rect 367560 377816 367612 377868
rect 463516 377816 463568 377868
rect 150992 377748 151044 377800
rect 198096 377748 198148 377800
rect 198464 377748 198516 377800
rect 298100 377748 298152 377800
rect 372988 377748 373040 377800
rect 455604 377748 455656 377800
rect 198004 377680 198056 377732
rect 295892 377680 295944 377732
rect 370320 377680 370372 377732
rect 453028 377680 453080 377732
rect 197544 377612 197596 377664
rect 293316 377612 293368 377664
rect 367652 377612 367704 377664
rect 451004 377612 451056 377664
rect 197084 377544 197136 377596
rect 290188 377544 290240 377596
rect 373172 377544 373224 377596
rect 428188 377544 428240 377596
rect 196716 377476 196768 377528
rect 287704 377476 287756 377528
rect 377220 377476 377272 377528
rect 410340 377476 410392 377528
rect 199384 377408 199436 377460
rect 280804 377408 280856 377460
rect 363512 377408 363564 377460
rect 379888 377408 379940 377460
rect 414572 377408 414624 377460
rect 196808 377340 196860 377392
rect 278412 377340 278464 377392
rect 366180 377340 366232 377392
rect 372252 377340 372304 377392
rect 402980 377340 403032 377392
rect 146024 377272 146076 377324
rect 207296 377272 207348 377324
rect 213092 377272 213144 377324
rect 270960 377272 271012 377324
rect 104256 377204 104308 377256
rect 215668 377204 215720 377256
rect 217048 377204 217100 377256
rect 217692 377204 217744 377256
rect 141056 377136 141108 377188
rect 201868 377136 201920 377188
rect 219256 377136 219308 377188
rect 264980 377204 265032 377256
rect 153568 377068 153620 377120
rect 200396 377068 200448 377120
rect 42524 377000 42576 377052
rect 199752 377000 199804 377052
rect 369768 377000 369820 377052
rect 47584 376932 47636 376984
rect 217048 376932 217100 376984
rect 369584 376796 369636 376848
rect 368388 376728 368440 376780
rect 378140 376728 378192 376780
rect 378600 376728 378652 376780
rect 198832 376660 198884 376712
rect 300860 376660 300912 376712
rect 357164 376660 357216 376712
rect 470876 376660 470928 376712
rect 99472 376592 99524 376644
rect 214380 376592 214432 376644
rect 219808 376592 219860 376644
rect 302516 376592 302568 376644
rect 364156 376592 364208 376644
rect 474740 376592 474792 376644
rect 101864 376524 101916 376576
rect 214012 376524 214064 376576
rect 214472 376524 214524 376576
rect 276112 376524 276164 376576
rect 367008 376524 367060 376576
rect 477500 376524 477552 376576
rect 97080 376456 97132 376508
rect 205916 376456 205968 376508
rect 206744 376456 206796 376508
rect 283104 376456 283156 376508
rect 374460 376456 374512 376508
rect 483388 376456 483440 376508
rect 107568 376388 107620 376440
rect 207296 376388 207348 376440
rect 207940 376388 207992 376440
rect 212908 376388 212960 376440
rect 273444 376388 273496 376440
rect 362776 376388 362828 376440
rect 467932 376388 467984 376440
rect 125968 376320 126020 376372
rect 204444 376320 204496 376372
rect 208952 376320 209004 376372
rect 263600 376320 263652 376372
rect 364800 376320 364852 376372
rect 465080 376320 465132 376372
rect 131028 376252 131080 376304
rect 199016 376252 199068 376304
rect 214932 376252 214984 376304
rect 268016 376252 268068 376304
rect 357072 376252 357124 376304
rect 422852 376252 422904 376304
rect 133512 376184 133564 376236
rect 194600 376184 194652 376236
rect 211620 376184 211672 376236
rect 260932 376184 260984 376236
rect 371792 376184 371844 376236
rect 430672 376184 430724 376236
rect 138480 376116 138532 376168
rect 195060 376116 195112 376168
rect 210240 376116 210292 376168
rect 258356 376116 258408 376168
rect 359464 376116 359516 376168
rect 418436 376116 418488 376168
rect 77116 376048 77168 376100
rect 204168 376048 204220 376100
rect 218612 376048 218664 376100
rect 265900 376048 265952 376100
rect 378600 376048 378652 376100
rect 436192 376048 436244 376100
rect 98552 375980 98604 376032
rect 213092 375980 213144 376032
rect 219440 375980 219492 376032
rect 359924 375980 359976 376032
rect 519084 375980 519136 376032
rect 208032 375912 208084 375964
rect 250628 375912 250680 375964
rect 370964 375912 371016 375964
rect 416044 375912 416096 375964
rect 217508 375844 217560 375896
rect 253388 375844 253440 375896
rect 375840 375844 375892 375896
rect 379336 375844 379388 375896
rect 408684 375844 408736 375896
rect 214012 375776 214064 375828
rect 217416 375776 217468 375828
rect 239772 375776 239824 375828
rect 215852 375708 215904 375760
rect 255964 375708 256016 375760
rect 219440 375640 219492 375692
rect 220084 375640 220136 375692
rect 100760 375300 100812 375352
rect 213920 375300 213972 375352
rect 214932 375300 214984 375352
rect 215576 375300 215628 375352
rect 262772 375300 262824 375352
rect 375932 375300 375984 375352
rect 376760 375300 376812 375352
rect 422576 375300 422628 375352
rect 199384 375232 199436 375284
rect 199568 375232 199620 375284
rect 216680 375232 216732 375284
rect 263876 375232 263928 375284
rect 372436 375232 372488 375284
rect 378140 375232 378192 375284
rect 379244 375232 379296 375284
rect 423956 375232 424008 375284
rect 367468 375164 367520 375216
rect 377220 375164 377272 375216
rect 409972 375164 410024 375216
rect 370228 375096 370280 375148
rect 377036 375096 377088 375148
rect 377128 375096 377180 375148
rect 415860 375096 415912 375148
rect 368204 375028 368256 375080
rect 378692 375028 378744 375080
rect 419356 375028 419408 375080
rect 365628 374960 365680 375012
rect 376576 374960 376628 375012
rect 418160 374960 418212 375012
rect 206560 374892 206612 374944
rect 219808 374892 219860 374944
rect 220636 374892 220688 374944
rect 215852 374824 215904 374876
rect 260564 374824 260616 374876
rect 362684 374824 362736 374876
rect 374460 374892 374512 374944
rect 416964 374892 417016 374944
rect 377036 374824 377088 374876
rect 425152 374824 425204 374876
rect 206192 374756 206244 374808
rect 216036 374756 216088 374808
rect 262220 374756 262272 374808
rect 357256 374756 357308 374808
rect 102968 374688 103020 374740
rect 214932 374688 214984 374740
rect 220636 374688 220688 374740
rect 266452 374688 266504 374740
rect 199384 374620 199436 374672
rect 359004 374688 359056 374740
rect 359648 374688 359700 374740
rect 361396 374756 361448 374808
rect 377128 374756 377180 374808
rect 378140 374756 378192 374808
rect 426440 374756 426492 374808
rect 367008 374688 367060 374740
rect 428280 374688 428332 374740
rect 362868 374620 362920 374672
rect 370964 374620 371016 374672
rect 432236 374620 432288 374672
rect 213920 374280 213972 374332
rect 215852 374280 215904 374332
rect 359832 373260 359884 373312
rect 519268 373260 519320 373312
rect 359464 372580 359516 372632
rect 359832 372580 359884 372632
rect 519268 372580 519320 372632
rect 519636 372580 519688 372632
rect 199568 371152 199620 371204
rect 199752 371152 199804 371204
rect 208492 371152 208544 371204
rect 359096 371152 359148 371204
rect 359740 370472 359792 370524
rect 519176 370472 519228 370524
rect 519544 370472 519596 370524
rect 359096 369180 359148 369232
rect 359556 369180 359608 369232
rect 519360 369180 519412 369232
rect 199476 369112 199528 369164
rect 358912 369112 358964 369164
rect 359740 369112 359792 369164
rect 182916 367752 182968 367804
rect 201592 367752 201644 367804
rect 342904 367752 342956 367804
rect 379244 365032 379296 365084
rect 379428 365032 379480 365084
rect 359648 364964 359700 365016
rect 518992 364964 519044 365016
rect 199660 363604 199712 363656
rect 359188 363468 359240 363520
rect 359924 363468 359976 363520
rect 199752 362176 199804 362228
rect 359464 362176 359516 362228
rect 359280 361564 359332 361616
rect 359464 361564 359516 361616
rect 202788 360816 202840 360868
rect 210424 360816 210476 360868
rect 197544 360136 197596 360188
rect 201776 360136 201828 360188
rect 500776 359660 500828 359712
rect 518072 359660 518124 359712
rect 498844 359592 498896 359644
rect 517980 359592 518032 359644
rect 197728 359524 197780 359576
rect 204536 359524 204588 359576
rect 277308 359524 277360 359576
rect 357440 359524 357492 359576
rect 438124 359524 438176 359576
rect 516600 359524 516652 359576
rect 190920 359456 190972 359508
rect 201500 359456 201552 359508
rect 202788 359456 202840 359508
rect 351736 359456 351788 359508
rect 358084 359456 358136 359508
rect 360292 359252 360344 359304
rect 361580 359252 361632 359304
rect 342260 358912 342312 358964
rect 343548 358912 343600 358964
rect 359096 358912 359148 358964
rect 179696 358844 179748 358896
rect 197544 358844 197596 358896
rect 339776 358844 339828 358896
rect 357348 358844 357400 358896
rect 362960 358844 363012 358896
rect 178592 358776 178644 358828
rect 197728 358776 197780 358828
rect 338488 358776 338540 358828
rect 360292 358776 360344 358828
rect 510896 358776 510948 358828
rect 511908 358776 511960 358828
rect 517520 358776 517572 358828
rect 3332 358708 3384 358760
rect 18604 358708 18656 358760
rect 218520 358708 218572 358760
rect 220820 358708 220872 358760
rect 379428 358708 379480 358760
rect 380900 358708 380952 358760
rect 218612 358436 218664 358488
rect 221096 358436 221148 358488
rect 375932 358368 375984 358420
rect 381268 358368 381320 358420
rect 217232 358232 217284 358284
rect 221004 358232 221056 358284
rect 373172 358096 373224 358148
rect 381176 358096 381228 358148
rect 182824 358028 182876 358080
rect 197728 358028 197780 358080
rect 342260 358028 342312 358080
rect 372436 358028 372488 358080
rect 381084 358028 381136 358080
rect 214472 357620 214524 357672
rect 220912 357620 220964 357672
rect 379336 357484 379388 357536
rect 380992 357484 381044 357536
rect 55772 357348 55824 357400
rect 60740 357348 60792 357400
rect 58624 355988 58676 356040
rect 59636 355988 59688 356040
rect 518164 353200 518216 353252
rect 580172 353200 580224 353252
rect 46296 300772 46348 300824
rect 56968 300772 57020 300824
rect 57060 300772 57112 300824
rect 58532 300772 58584 300824
rect 520188 288396 520240 288448
rect 580264 288396 580316 288448
rect 519176 287036 519228 287088
rect 519636 287036 519688 287088
rect 580356 287036 580408 287088
rect 200764 284248 200816 284300
rect 216680 284248 216732 284300
rect 358636 284248 358688 284300
rect 376944 284248 376996 284300
rect 201500 282820 201552 282872
rect 216680 282820 216732 282872
rect 361304 282820 361356 282872
rect 376760 282820 376812 282872
rect 203892 282752 203944 282804
rect 216772 282752 216824 282804
rect 200764 282412 200816 282464
rect 201500 282412 201552 282464
rect 54484 282140 54536 282192
rect 57980 282140 58032 282192
rect 376944 281528 376996 281580
rect 45468 281460 45520 281512
rect 57244 281460 57296 281512
rect 57520 281460 57572 281512
rect 358084 281460 358136 281512
rect 360200 281460 360252 281512
rect 45284 273640 45336 273692
rect 145932 273640 145984 273692
rect 42616 273572 42668 273624
rect 131028 273572 131080 273624
rect 372528 273572 372580 273624
rect 379244 273572 379296 273624
rect 43352 273504 43404 273556
rect 133420 273504 133472 273556
rect 369032 273504 369084 273556
rect 378140 273504 378192 273556
rect 378600 273504 378652 273556
rect 379428 273504 379480 273556
rect 379796 273504 379848 273556
rect 427636 273504 427688 273556
rect 45192 273436 45244 273488
rect 135904 273436 135956 273488
rect 212080 273436 212132 273488
rect 250720 273436 250772 273488
rect 361212 273436 361264 273488
rect 416044 273436 416096 273488
rect 45008 273368 45060 273420
rect 138480 273368 138532 273420
rect 211712 273368 211764 273420
rect 272248 273368 272300 273420
rect 373172 273368 373224 273420
rect 433340 273368 433392 273420
rect 45100 273300 45152 273352
rect 140872 273300 140924 273352
rect 212816 273300 212868 273352
rect 273260 273300 273312 273352
rect 368112 273300 368164 273352
rect 440884 273300 440936 273352
rect 52368 273232 52420 273284
rect 57980 273232 58032 273284
rect 58808 273232 58860 273284
rect 50528 272960 50580 273012
rect 53840 272960 53892 273012
rect 46480 272892 46532 272944
rect 50988 272892 51040 272944
rect 207848 273232 207900 273284
rect 280896 273232 280948 273284
rect 358452 273232 358504 273284
rect 430948 273232 431000 273284
rect 374460 273164 374512 273216
rect 396724 273164 396776 273216
rect 379244 273096 379296 273148
rect 423772 273096 423824 273148
rect 378600 273028 378652 273080
rect 426440 273028 426492 273080
rect 366824 272960 366876 273012
rect 423404 272960 423456 273012
rect 98092 272892 98144 272944
rect 356888 272892 356940 272944
rect 428188 272892 428240 272944
rect 54852 272824 54904 272876
rect 88340 272824 88392 272876
rect 210884 272824 210936 272876
rect 283380 272824 283432 272876
rect 369492 272824 369544 272876
rect 468484 272824 468536 272876
rect 58808 272756 58860 272808
rect 99380 272756 99432 272808
rect 216128 272756 216180 272808
rect 295892 272756 295944 272808
rect 372160 272756 372212 272808
rect 470876 272756 470928 272808
rect 49056 272688 49108 272740
rect 90732 272688 90784 272740
rect 209596 272688 209648 272740
rect 290924 272688 290976 272740
rect 373724 272688 373776 272740
rect 478420 272688 478472 272740
rect 50436 272620 50488 272672
rect 93676 272620 93728 272672
rect 203800 272620 203852 272672
rect 288164 272620 288216 272672
rect 376300 272620 376352 272672
rect 480812 272620 480864 272672
rect 51816 272552 51868 272604
rect 98460 272552 98512 272604
rect 205180 272552 205232 272604
rect 298468 272552 298520 272604
rect 363972 272552 364024 272604
rect 475844 272552 475896 272604
rect 47952 272484 48004 272536
rect 95884 272484 95936 272536
rect 200948 272484 201000 272536
rect 300860 272484 300912 272536
rect 362592 272484 362644 272536
rect 473452 272484 473504 272536
rect 55772 272416 55824 272468
rect 59636 272416 59688 272468
rect 59728 272416 59780 272468
rect 60832 272416 60884 272468
rect 48044 272348 48096 272400
rect 77116 272348 77168 272400
rect 377036 272348 377088 272400
rect 379704 272348 379756 272400
rect 48964 272280 49016 272332
rect 54300 272280 54352 272332
rect 83004 272280 83056 272332
rect 374460 272280 374512 272332
rect 375196 272280 375248 272332
rect 67548 272212 67600 272264
rect 95976 272212 96028 272264
rect 53840 272144 53892 272196
rect 54116 272144 54168 272196
rect 85396 272144 85448 272196
rect 46388 272076 46440 272128
rect 75920 272076 75972 272128
rect 60832 272008 60884 272060
rect 94228 272008 94280 272060
rect 379612 272008 379664 272060
rect 380072 272008 380124 272060
rect 54208 271940 54260 271992
rect 54760 271940 54812 271992
rect 88340 271940 88392 271992
rect 379704 271940 379756 271992
rect 425060 271940 425112 271992
rect 58532 271872 58584 271924
rect 102140 271872 102192 271924
rect 213644 271872 213696 271924
rect 215668 271872 215720 271924
rect 236000 271872 236052 271924
rect 45376 271804 45428 271856
rect 143540 271804 143592 271856
rect 154488 271804 154540 271856
rect 200120 271804 200172 271856
rect 212172 271804 212224 271856
rect 307760 271804 307812 271856
rect 43444 271668 43496 271720
rect 125600 271736 125652 271788
rect 157248 271736 157300 271788
rect 201684 271736 201736 271788
rect 219532 271736 219584 271788
rect 219808 271736 219860 271788
rect 223580 271736 223632 271788
rect 302240 271736 302292 271788
rect 47676 271668 47728 271720
rect 47952 271668 48004 271720
rect 41052 271600 41104 271652
rect 107660 271668 107712 271720
rect 158628 271668 158680 271720
rect 197360 271668 197412 271720
rect 200856 271668 200908 271720
rect 270500 271668 270552 271720
rect 54668 271600 54720 271652
rect 120080 271600 120132 271652
rect 202328 271600 202380 271652
rect 264980 271600 265032 271652
rect 46664 271532 46716 271584
rect 52460 271532 52512 271584
rect 56876 271532 56928 271584
rect 123116 271532 123168 271584
rect 164148 271532 164200 271584
rect 197452 271532 197504 271584
rect 203708 271532 203760 271584
rect 263600 271532 263652 271584
rect 343548 271532 343600 271584
rect 359096 271872 359148 271924
rect 370412 271872 370464 271924
rect 428004 271872 428056 271924
rect 440148 271872 440200 271924
rect 516600 271872 516652 271924
rect 368020 271804 368072 271856
rect 458180 271804 458232 271856
rect 366732 271736 366784 271788
rect 455788 271736 455840 271788
rect 362500 271668 362552 271720
rect 449900 271668 449952 271720
rect 367008 271600 367060 271652
rect 370412 271600 370464 271652
rect 376392 271600 376444 271652
rect 460940 271600 460992 271652
rect 357072 271532 357124 271584
rect 369400 271532 369452 271584
rect 452660 271532 452712 271584
rect 53012 271464 53064 271516
rect 117320 271464 117372 271516
rect 161388 271464 161440 271516
rect 202972 271464 203024 271516
rect 216312 271464 216364 271516
rect 276112 271464 276164 271516
rect 365444 271464 365496 271516
rect 443000 271464 443052 271516
rect 46112 271396 46164 271448
rect 46664 271396 46716 271448
rect 52828 271396 52880 271448
rect 115940 271396 115992 271448
rect 197360 271396 197412 271448
rect 197728 271396 197780 271448
rect 216496 271396 216548 271448
rect 273260 271396 273312 271448
rect 343456 271396 343508 271448
rect 358820 271396 358872 271448
rect 370872 271396 370924 271448
rect 447140 271396 447192 271448
rect 53196 271328 53248 271380
rect 113548 271328 113600 271380
rect 214840 271328 214892 271380
rect 223580 271328 223632 271380
rect 224224 271328 224276 271380
rect 268016 271328 268068 271380
rect 278688 271328 278740 271380
rect 357440 271328 357492 271380
rect 372068 271328 372120 271380
rect 445760 271328 445812 271380
rect 52920 271260 52972 271312
rect 110420 271260 110472 271312
rect 183468 271260 183520 271312
rect 197360 271260 197412 271312
rect 205088 271260 205140 271312
rect 255320 271260 255372 271312
rect 277216 271260 277268 271312
rect 357164 271260 357216 271312
rect 358820 271260 358872 271312
rect 360016 271260 360068 271312
rect 366916 271260 366968 271312
rect 434720 271260 434772 271312
rect 503628 271260 503680 271312
rect 517704 271260 517756 271312
rect 51724 271192 51776 271244
rect 104900 271192 104952 271244
rect 210700 271192 210752 271244
rect 260840 271192 260892 271244
rect 280068 271192 280120 271244
rect 367928 271192 367980 271244
rect 51908 271124 51960 271176
rect 103520 271124 103572 271176
rect 183468 271124 183520 271176
rect 201592 271124 201644 271176
rect 209504 271124 209556 271176
rect 258264 271124 258316 271176
rect 275928 271124 275980 271176
rect 356612 271124 356664 271176
rect 356888 271124 356940 271176
rect 373540 271124 373592 271176
rect 50252 271056 50304 271108
rect 100760 271056 100812 271108
rect 219532 271056 219584 271108
rect 268108 271056 268160 271108
rect 375104 271056 375156 271108
rect 420920 271056 420972 271108
rect 46664 270988 46716 271040
rect 77300 270988 77352 271040
rect 210792 270988 210844 271040
rect 252560 270988 252612 271040
rect 373632 270988 373684 271040
rect 418344 270988 418396 271040
rect 437480 271124 437532 271176
rect 503536 271124 503588 271176
rect 517612 271124 517664 271176
rect 433340 271056 433392 271108
rect 47952 270920 48004 270972
rect 78680 270920 78732 270972
rect 219164 270920 219216 270972
rect 247040 270920 247092 270972
rect 375012 270920 375064 270972
rect 409880 270920 409932 270972
rect 215208 270852 215260 270904
rect 224224 270852 224276 270904
rect 264244 270852 264296 270904
rect 266360 270852 266412 270904
rect 425704 270852 425756 270904
rect 429200 270852 429252 270904
rect 517612 270784 517664 270836
rect 517888 270784 517940 270836
rect 422944 270580 422996 270632
rect 437480 270580 437532 270632
rect 102784 270512 102836 270564
rect 113180 270512 113232 270564
rect 268844 270512 268896 270564
rect 273260 270512 273312 270564
rect 421564 270512 421616 270564
rect 436100 270512 436152 270564
rect 44916 270444 44968 270496
rect 147680 270444 147732 270496
rect 210332 270444 210384 270496
rect 210884 270444 210936 270496
rect 211528 270444 211580 270496
rect 216956 270444 217008 270496
rect 224224 270444 224276 270496
rect 262220 270444 262272 270496
rect 369768 270444 369820 270496
rect 371700 270444 371752 270496
rect 379336 270444 379388 270496
rect 379520 270444 379572 270496
rect 379980 270444 380032 270496
rect 396080 270444 396132 270496
rect 58716 270376 58768 270428
rect 115940 270376 115992 270428
rect 212356 270376 212408 270428
rect 244280 270376 244332 270428
rect 378600 270376 378652 270428
rect 379612 270376 379664 270428
rect 380072 270376 380124 270428
rect 411260 270376 411312 270428
rect 60740 270308 60792 270360
rect 91100 270308 91152 270360
rect 210976 270308 211028 270360
rect 214840 270308 214892 270360
rect 219624 270308 219676 270360
rect 220452 270308 220504 270360
rect 249800 270308 249852 270360
rect 368296 270308 368348 270360
rect 398840 270308 398892 270360
rect 79048 270240 79100 270292
rect 110420 270240 110472 270292
rect 220176 270240 220228 270292
rect 248512 270240 248564 270292
rect 377036 270240 377088 270292
rect 380072 270240 380124 270292
rect 58624 270172 58676 270224
rect 89720 270172 89772 270224
rect 217232 270172 217284 270224
rect 219900 270172 219952 270224
rect 251272 270172 251324 270224
rect 376484 270172 376536 270224
rect 405740 270240 405792 270292
rect 380256 270172 380308 270224
rect 404360 270172 404412 270224
rect 56508 270104 56560 270156
rect 86960 270104 87012 270156
rect 210884 270104 210936 270156
rect 239128 270104 239180 270156
rect 371700 270104 371752 270156
rect 397460 270104 397512 270156
rect 59360 270036 59412 270088
rect 92480 270036 92532 270088
rect 215208 270036 215260 270088
rect 219440 270036 219492 270088
rect 220544 270036 220596 270088
rect 220636 270036 220688 270088
rect 251180 270036 251232 270088
rect 371148 270036 371200 270088
rect 375748 270036 375800 270088
rect 403532 270036 403584 270088
rect 51724 269968 51776 270020
rect 84200 269968 84252 270020
rect 217140 269968 217192 270020
rect 217324 269968 217376 270020
rect 53104 269900 53156 269952
rect 85580 269900 85632 269952
rect 88248 269900 88300 269952
rect 106280 269900 106332 269952
rect 214288 269900 214340 269952
rect 214932 269900 214984 269952
rect 220728 269968 220780 270020
rect 252560 269968 252612 270020
rect 371056 269968 371108 270020
rect 372068 269968 372120 270020
rect 400220 269968 400272 270020
rect 263600 269900 263652 269952
rect 376668 269900 376720 269952
rect 389180 269900 389232 269952
rect 419540 269900 419592 269952
rect 57980 269832 58032 269884
rect 103704 269832 103756 269884
rect 115848 269832 115900 269884
rect 196716 269832 196768 269884
rect 204352 269832 204404 269884
rect 214840 269832 214892 269884
rect 269120 269832 269172 269884
rect 373816 269832 373868 269884
rect 375840 269832 375892 269884
rect 407120 269832 407172 269884
rect 56876 269764 56928 269816
rect 104900 269764 104952 269816
rect 114468 269764 114520 269816
rect 196624 269764 196676 269816
rect 202880 269764 202932 269816
rect 206836 269764 206888 269816
rect 213000 269764 213052 269816
rect 270500 269764 270552 269816
rect 379520 269764 379572 269816
rect 413008 269764 413060 269816
rect 62120 269696 62172 269748
rect 91192 269696 91244 269748
rect 216956 269696 217008 269748
rect 245660 269696 245712 269748
rect 372344 269696 372396 269748
rect 375288 269696 375340 269748
rect 401692 269696 401744 269748
rect 81440 269628 81492 269680
rect 107660 269628 107712 269680
rect 206928 269628 206980 269680
rect 210792 269628 210844 269680
rect 237380 269628 237432 269680
rect 391940 269628 391992 269680
rect 83464 269560 83516 269612
rect 106372 269560 106424 269612
rect 220544 269560 220596 269612
rect 247040 269560 247092 269612
rect 375104 269560 375156 269612
rect 376576 269560 376628 269612
rect 379612 269560 379664 269612
rect 411352 269560 411404 269612
rect 214932 269492 214984 269544
rect 224224 269492 224276 269544
rect 374552 269492 374604 269544
rect 379980 269492 380032 269544
rect 218520 269288 218572 269340
rect 219440 269288 219492 269340
rect 220728 269288 220780 269340
rect 218612 269220 218664 269272
rect 219808 269220 219860 269272
rect 220636 269220 220688 269272
rect 216496 269152 216548 269204
rect 220176 269152 220228 269204
rect 373632 269152 373684 269204
rect 376484 269152 376536 269204
rect 219164 269084 219216 269136
rect 220452 269084 220504 269136
rect 373724 269084 373776 269136
rect 375196 269084 375248 269136
rect 380256 269084 380308 269136
rect 48136 269016 48188 269068
rect 53104 269016 53156 269068
rect 205640 269016 205692 269068
rect 256700 269016 256752 269068
rect 370964 269016 371016 269068
rect 373540 269016 373592 269068
rect 376760 269016 376812 269068
rect 377128 269016 377180 269068
rect 377220 269016 377272 269068
rect 379060 269016 379112 269068
rect 379244 269016 379296 269068
rect 420920 269016 420972 269068
rect 46848 268948 46900 269000
rect 51724 268948 51776 269000
rect 217232 268948 217284 269000
rect 217968 268948 218020 269000
rect 255320 268948 255372 269000
rect 44088 268880 44140 268932
rect 59360 268880 59412 268932
rect 219716 268880 219768 268932
rect 253940 268880 253992 268932
rect 378692 268948 378744 269000
rect 418528 268948 418580 269000
rect 415400 268880 415452 268932
rect 43628 268812 43680 268864
rect 56876 268812 56928 268864
rect 213736 268812 213788 268864
rect 244372 268812 244424 268864
rect 376576 268812 376628 268864
rect 378692 268812 378744 268864
rect 48228 268744 48280 268796
rect 58624 268744 58676 268796
rect 216404 268744 216456 268796
rect 242900 268744 242952 268796
rect 374460 268744 374512 268796
rect 379244 268812 379296 268864
rect 379888 268812 379940 268864
rect 414020 268812 414072 268864
rect 379152 268744 379204 268796
rect 408500 268744 408552 268796
rect 46756 268676 46808 268728
rect 55772 268676 55824 268728
rect 56508 268676 56560 268728
rect 214472 268676 214524 268728
rect 236000 268676 236052 268728
rect 391940 268676 391992 268728
rect 418160 268676 418212 268728
rect 43996 268608 44048 268660
rect 48136 268608 48188 268660
rect 60740 268608 60792 268660
rect 213092 268608 213144 268660
rect 233240 268608 233292 268660
rect 258080 268608 258132 268660
rect 46572 268540 46624 268592
rect 48228 268540 48280 268592
rect 62120 268540 62172 268592
rect 214380 268540 214432 268592
rect 231860 268540 231912 268592
rect 259460 268540 259512 268592
rect 43720 268472 43772 268524
rect 47584 268472 47636 268524
rect 79048 268472 79100 268524
rect 215852 268472 215904 268524
rect 230480 268472 230532 268524
rect 259552 268472 259604 268524
rect 372252 268472 372304 268524
rect 379244 268472 379296 268524
rect 402980 268472 403032 268524
rect 43904 268404 43956 268456
rect 47768 268404 47820 268456
rect 81440 268404 81492 268456
rect 208308 268404 208360 268456
rect 214472 268404 214524 268456
rect 230388 268404 230440 268456
rect 260840 268404 260892 268456
rect 379060 268404 379112 268456
rect 409880 268404 409932 268456
rect 43812 268336 43864 268388
rect 47676 268336 47728 268388
rect 88248 268336 88300 268388
rect 207572 268336 207624 268388
rect 212172 268336 212224 268388
rect 268844 268336 268896 268388
rect 373540 268336 373592 268388
rect 431960 268336 432012 268388
rect 43536 268268 43588 268320
rect 128360 268268 128412 268320
rect 40960 268200 41012 268252
rect 57980 268200 58032 268252
rect 60740 268200 60792 268252
rect 60924 268200 60976 268252
rect 377956 268200 378008 268252
rect 379152 268200 379204 268252
rect 357532 253988 357584 254040
rect 360292 253988 360344 254040
rect 198648 253852 198700 253904
rect 200764 253852 200816 253904
rect 340788 253852 340840 253904
rect 357348 253920 357400 253972
rect 357624 253920 357676 253972
rect 180156 253308 180208 253360
rect 197452 253308 197504 253360
rect 500868 253308 500920 253360
rect 517704 253308 517756 253360
rect 339408 253240 339460 253292
rect 357532 253240 357584 253292
rect 357716 253240 357768 253292
rect 499212 253240 499264 253292
rect 517612 253240 517664 253292
rect 517980 253240 518032 253292
rect 179328 253172 179380 253224
rect 197636 253172 197688 253224
rect 351828 253172 351880 253224
rect 360200 253172 360252 253224
rect 517704 253172 517756 253224
rect 518072 253172 518124 253224
rect 191748 252560 191800 252612
rect 198648 252560 198700 252612
rect 510896 252560 510948 252612
rect 517520 252560 517572 252612
rect 217968 252492 218020 252544
rect 265624 252492 265676 252544
rect 218428 252424 218480 252476
rect 219256 252424 219308 252476
rect 264980 252424 265032 252476
rect 58716 252016 58768 252068
rect 60832 252016 60884 252068
rect 216128 252016 216180 252068
rect 229100 252016 229152 252068
rect 379152 252016 379204 252068
rect 396724 252016 396776 252068
rect 58532 251948 58584 252000
rect 83464 251948 83516 252000
rect 216220 251948 216272 252000
rect 230480 251948 230532 252000
rect 372436 251948 372488 252000
rect 376392 251948 376444 252000
rect 425704 251948 425756 252000
rect 68376 251880 68428 251932
rect 96620 251880 96672 251932
rect 218612 251880 218664 251932
rect 233240 251880 233292 251932
rect 368388 251880 368440 251932
rect 371148 251880 371200 251932
rect 421564 251880 421616 251932
rect 53840 251812 53892 251864
rect 102784 251812 102836 251864
rect 216036 251812 216088 251864
rect 218520 251812 218572 251864
rect 264244 251812 264296 251864
rect 343548 251812 343600 251864
rect 360292 251812 360344 251864
rect 369676 251812 369728 251864
rect 371056 251812 371108 251864
rect 422944 251812 422996 251864
rect 49148 250452 49200 250504
rect 54852 250452 54904 250504
rect 68376 250452 68428 250504
rect 519360 183540 519412 183592
rect 520188 183540 520240 183592
rect 580264 183540 580316 183592
rect 520096 183472 520148 183524
rect 580356 183472 580408 183524
rect 209412 177964 209464 178016
rect 216680 177964 216732 178016
rect 365352 177964 365404 178016
rect 377036 177964 377088 178016
rect 360200 176604 360252 176656
rect 376944 176604 376996 176656
rect 358728 176128 358780 176180
rect 360200 176128 360252 176180
rect 198004 175924 198056 175976
rect 198648 175924 198700 175976
rect 216680 175924 216732 175976
rect 204996 175176 205048 175228
rect 216680 175176 216732 175228
rect 362408 175176 362460 175228
rect 377220 175176 377272 175228
rect 52092 166948 52144 167000
rect 101036 166948 101088 167000
rect 366640 166948 366692 167000
rect 423404 166948 423456 167000
rect 49332 166880 49384 166932
rect 98460 166880 98512 166932
rect 358268 166880 358320 166932
rect 416044 166880 416096 166932
rect 52276 166812 52328 166864
rect 105820 166812 105872 166864
rect 202236 166812 202288 166864
rect 253572 166812 253624 166864
rect 356704 166812 356756 166864
rect 418436 166812 418488 166864
rect 50712 166744 50764 166796
rect 108212 166744 108264 166796
rect 209228 166744 209280 166796
rect 270868 166744 270920 166796
rect 356796 166744 356848 166796
rect 425980 166744 426032 166796
rect 56232 166676 56284 166728
rect 138480 166676 138532 166728
rect 202420 166676 202472 166728
rect 265900 166676 265952 166728
rect 370780 166676 370832 166728
rect 473452 166676 473504 166728
rect 59820 166608 59872 166660
rect 143540 166608 143592 166660
rect 206376 166608 206428 166660
rect 288256 166608 288308 166660
rect 367836 166608 367888 166660
rect 475844 166608 475896 166660
rect 59084 166540 59136 166592
rect 145932 166540 145984 166592
rect 209320 166540 209372 166592
rect 298468 166540 298520 166592
rect 369308 166540 369360 166592
rect 478420 166540 478472 166592
rect 59912 166472 59964 166524
rect 150900 166472 150952 166524
rect 211988 166472 212040 166524
rect 303528 166472 303580 166524
rect 371976 166472 372028 166524
rect 480904 166472 480956 166524
rect 58992 166404 59044 166456
rect 153292 166404 153344 166456
rect 203616 166404 203668 166456
rect 295892 166404 295944 166456
rect 361120 166404 361172 166456
rect 470968 166404 471020 166456
rect 42708 166336 42760 166388
rect 163320 166336 163372 166388
rect 213460 166336 213512 166388
rect 308496 166336 308548 166388
rect 373356 166336 373408 166388
rect 485964 166336 486016 166388
rect 41144 166268 41196 166320
rect 165896 166268 165948 166320
rect 214748 166268 214800 166320
rect 315856 166268 315908 166320
rect 365260 166268 365312 166320
rect 483388 166268 483440 166320
rect 50804 166200 50856 166252
rect 96068 166200 96120 166252
rect 374920 166200 374972 166252
rect 428188 166200 428240 166252
rect 365168 166132 365220 166184
rect 408132 166132 408184 166184
rect 370412 166064 370464 166116
rect 380900 166064 380952 166116
rect 54392 165588 54444 165640
rect 113272 165588 113324 165640
rect 55864 165520 55916 165572
rect 132500 165520 132552 165572
rect 211896 165520 211948 165572
rect 310980 165520 311032 165572
rect 343272 165520 343324 165572
rect 357072 165520 357124 165572
rect 357532 165520 357584 165572
rect 362316 165520 362368 165572
rect 452660 165520 452712 165572
rect 55128 165452 55180 165504
rect 129740 165452 129792 165504
rect 210516 165452 210568 165504
rect 293316 165452 293368 165504
rect 369216 165452 369268 165504
rect 455420 165452 455472 165504
rect 55956 165384 56008 165436
rect 128360 165384 128412 165436
rect 219072 165384 219124 165436
rect 300860 165384 300912 165436
rect 358360 165384 358412 165436
rect 443000 165384 443052 165436
rect 54944 165316 54996 165368
rect 125876 165316 125928 165368
rect 213368 165316 213420 165368
rect 285956 165316 286008 165368
rect 370596 165316 370648 165368
rect 449900 165316 449952 165368
rect 56140 165248 56192 165300
rect 123484 165248 123536 165300
rect 211804 165248 211856 165300
rect 276020 165248 276072 165300
rect 378968 165248 379020 165300
rect 458364 165248 458416 165300
rect 53380 165180 53432 165232
rect 120908 165180 120960 165232
rect 214656 165180 214708 165232
rect 278412 165180 278464 165232
rect 371884 165180 371936 165232
rect 447324 165180 447376 165232
rect 56876 165112 56928 165164
rect 57336 165112 57388 165164
rect 59820 165112 59872 165164
rect 115940 165112 115992 165164
rect 183192 165112 183244 165164
rect 197360 165112 197412 165164
rect 218888 165112 218940 165164
rect 280804 165112 280856 165164
rect 366548 165112 366600 165164
rect 440240 165112 440292 165164
rect 503628 165112 503680 165164
rect 517796 165112 517848 165164
rect 55036 165044 55088 165096
rect 118332 165044 118384 165096
rect 204904 165044 204956 165096
rect 263600 165044 263652 165096
rect 361028 165044 361080 165096
rect 422944 165044 422996 165096
rect 53564 164976 53616 165028
rect 113548 164976 113600 165028
rect 183468 164976 183520 165028
rect 201500 164976 201552 165028
rect 215944 164976 215996 165028
rect 273444 164976 273496 165028
rect 373448 164976 373500 165028
rect 445760 164976 445812 165028
rect 503260 164976 503312 165028
rect 517888 165044 517940 165096
rect 52000 164908 52052 164960
rect 59820 164908 59872 164960
rect 59912 164908 59964 164960
rect 103520 164908 103572 164960
rect 116032 164908 116084 164960
rect 196716 164908 196768 164960
rect 210608 164908 210660 164960
rect 267740 164908 267792 164960
rect 363880 164908 363932 164960
rect 434812 164908 434864 164960
rect 440240 164908 440292 164960
rect 516600 164976 516652 165028
rect 510528 164908 510580 164960
rect 517520 164908 517572 164960
rect 57336 164840 57388 164892
rect 104900 164840 104952 164892
rect 114560 164840 114612 164892
rect 196624 164840 196676 164892
rect 207664 164840 207716 164892
rect 258080 164840 258132 164892
rect 343548 164840 343600 164892
rect 360292 164840 360344 164892
rect 369124 164840 369176 164892
rect 437756 164840 437808 164892
rect 50896 164772 50948 164824
rect 59912 164772 59964 164824
rect 49424 164636 49476 164688
rect 89904 164772 89956 164824
rect 206284 164772 206336 164824
rect 255320 164772 255372 164824
rect 378876 164772 378928 164824
rect 420920 164772 420972 164824
rect 422944 164772 422996 164824
rect 433340 164772 433392 164824
rect 56048 164568 56100 164620
rect 88340 164704 88392 164756
rect 209136 164704 209188 164756
rect 249800 164704 249852 164756
rect 378784 164704 378836 164756
rect 413560 164704 413612 164756
rect 214564 164636 214616 164688
rect 247040 164636 247092 164688
rect 376116 164636 376168 164688
rect 410432 164636 410484 164688
rect 428832 164500 428884 164552
rect 433340 164500 433392 164552
rect 83464 164432 83516 164484
rect 107752 164432 107804 164484
rect 97264 164364 97316 164416
rect 100760 164364 100812 164416
rect 88984 164296 89036 164348
rect 106280 164296 106332 164348
rect 269764 164228 269816 164280
rect 273812 164228 273864 164280
rect 47584 164160 47636 164212
rect 52276 164160 52328 164212
rect 54576 164160 54628 164212
rect 57520 164160 57572 164212
rect 116400 164160 116452 164212
rect 214288 164160 214340 164212
rect 215760 164160 215812 164212
rect 219532 164160 219584 164212
rect 219992 164160 220044 164212
rect 267740 164160 267792 164212
rect 377312 164160 377364 164212
rect 437848 164160 437900 164212
rect 55680 164092 55732 164144
rect 59636 164092 59688 164144
rect 117872 164092 117924 164144
rect 370688 164092 370740 164144
rect 430580 164092 430632 164144
rect 53472 164024 53524 164076
rect 110880 164024 110932 164076
rect 376392 164024 376444 164076
rect 429292 164024 429344 164076
rect 53012 163956 53064 164008
rect 109684 163956 109736 164008
rect 379796 163956 379848 164008
rect 426440 163956 426492 164008
rect 379704 163888 379756 163940
rect 425060 163888 425112 163940
rect 379152 163820 379204 163872
rect 416872 163820 416924 163872
rect 59084 163752 59136 163804
rect 95240 163752 95292 163804
rect 374552 163752 374604 163804
rect 396080 163752 396132 163804
rect 50988 163684 51040 163736
rect 55036 163684 55088 163736
rect 98000 163684 98052 163736
rect 217140 163684 217192 163736
rect 219072 163684 219124 163736
rect 263784 163684 263836 163736
rect 374368 163684 374420 163736
rect 396172 163684 396224 163736
rect 52276 163616 52328 163668
rect 111156 163616 111208 163668
rect 215760 163616 215812 163668
rect 262220 163616 262272 163668
rect 50344 163548 50396 163600
rect 53564 163548 53616 163600
rect 111892 163548 111944 163600
rect 220728 163548 220780 163600
rect 266452 163548 266504 163600
rect 375196 163548 375248 163600
rect 430672 163548 430724 163600
rect 52736 163480 52788 163532
rect 59084 163480 59136 163532
rect 59452 163480 59504 163532
rect 118884 163480 118936 163532
rect 218888 163480 218940 163532
rect 219256 163480 219308 163532
rect 266544 163480 266596 163532
rect 371148 163480 371200 163532
rect 375840 163480 375892 163532
rect 436100 163480 436152 163532
rect 372160 163140 372212 163192
rect 374276 163140 374328 163192
rect 375196 163140 375248 163192
rect 218520 162936 218572 162988
rect 219532 162936 219584 162988
rect 220728 162936 220780 162988
rect 217232 162800 217284 162852
rect 217968 162800 218020 162852
rect 216128 162732 216180 162784
rect 260840 162800 260892 162852
rect 375104 162800 375156 162852
rect 379612 162800 379664 162852
rect 214656 162528 214708 162580
rect 216220 162528 216272 162580
rect 259552 162732 259604 162784
rect 375012 162732 375064 162784
rect 434812 162800 434864 162852
rect 379888 162732 379940 162784
rect 428832 162732 428884 162784
rect 218888 162664 218940 162716
rect 259460 162664 259512 162716
rect 374460 162664 374512 162716
rect 420920 162664 420972 162716
rect 218612 162596 218664 162648
rect 258172 162596 258224 162648
rect 376760 162460 376812 162512
rect 378048 162460 378100 162512
rect 378140 162460 378192 162512
rect 419540 162596 419592 162648
rect 376484 162392 376536 162444
rect 379888 162392 379940 162444
rect 379612 162188 379664 162240
rect 418252 162188 418304 162240
rect 220176 162120 220228 162172
rect 256700 162120 256752 162172
rect 373540 162120 373592 162172
rect 375196 162120 375248 162172
rect 431960 162120 432012 162172
rect 214748 161848 214800 161900
rect 216680 161848 216732 161900
rect 378048 161508 378100 161560
rect 395344 161508 395396 161560
rect 217968 161440 218020 161492
rect 235264 161440 235316 161492
rect 376668 161440 376720 161492
rect 396724 161440 396776 161492
rect 205548 161372 205600 161424
rect 220176 161372 220228 161424
rect 219808 156612 219860 156664
rect 220084 156612 220136 156664
rect 219440 156476 219492 156528
rect 219808 156476 219860 156528
rect 219440 156340 219492 156392
rect 220176 156340 220228 156392
rect 57980 148996 58032 149048
rect 103612 148996 103664 149048
rect 212816 148996 212868 149048
rect 274640 148996 274692 149048
rect 274732 148996 274784 149048
rect 275284 148996 275336 149048
rect 356888 148996 356940 149048
rect 379520 148996 379572 149048
rect 412732 148996 412784 149048
rect 58808 148928 58860 148980
rect 102140 148928 102192 148980
rect 212172 148928 212224 148980
rect 269764 148928 269816 148980
rect 375288 148928 375340 148980
rect 401600 148928 401652 148980
rect 213644 148860 213696 148912
rect 240140 148860 240192 148912
rect 47768 148792 47820 148844
rect 59912 148792 59964 148844
rect 83464 148792 83516 148844
rect 47952 148724 48004 148776
rect 52092 148724 52144 148776
rect 78680 148724 78732 148776
rect 47860 148656 47912 148708
rect 52000 148656 52052 148708
rect 80060 148656 80112 148708
rect 49056 148588 49108 148640
rect 53380 148588 53432 148640
rect 81440 148588 81492 148640
rect 374920 148588 374972 148640
rect 375288 148588 375340 148640
rect 56048 148520 56100 148572
rect 58808 148520 58860 148572
rect 58992 148520 59044 148572
rect 88984 148520 89036 148572
rect 212908 148520 212960 148572
rect 213644 148520 213696 148572
rect 58532 148452 58584 148504
rect 59820 148452 59872 148504
rect 107660 148452 107712 148504
rect 210884 148452 210936 148504
rect 213460 148452 213512 148504
rect 238760 148452 238812 148504
rect 375288 148452 375340 148504
rect 398840 148452 398892 148504
rect 54944 148384 54996 148436
rect 116032 148384 116084 148436
rect 213736 148384 213788 148436
rect 241520 148384 241572 148436
rect 372068 148384 372120 148436
rect 373356 148384 373408 148436
rect 400220 148384 400272 148436
rect 53196 148316 53248 148368
rect 114560 148316 114612 148368
rect 213092 148316 213144 148368
rect 274732 148316 274784 148368
rect 373172 148316 373224 148368
rect 374552 148316 374604 148368
rect 434720 148316 434772 148368
rect 47676 148248 47728 148300
rect 58532 148248 58584 148300
rect 58992 148248 59044 148300
rect 56140 147636 56192 147688
rect 57980 147636 58032 147688
rect 212816 147636 212868 147688
rect 208124 147568 208176 147620
rect 213368 147568 213420 147620
rect 213736 147568 213788 147620
rect 379336 147636 379388 147688
rect 379520 147636 379572 147688
rect 368296 147500 368348 147552
rect 374828 147500 374880 147552
rect 375288 147500 375340 147552
rect 213736 147432 213788 147484
rect 60096 146276 60148 146328
rect 215852 146276 215904 146328
rect 277400 146276 277452 146328
rect 46664 146208 46716 146260
rect 51908 146208 51960 146260
rect 55772 146208 55824 146260
rect 56232 146208 56284 146260
rect 58624 146208 58676 146260
rect 58900 146208 58952 146260
rect 58992 146208 59044 146260
rect 59360 146208 59412 146260
rect 92480 146208 92532 146260
rect 179052 146208 179104 146260
rect 197544 146208 197596 146260
rect 219716 146208 219768 146260
rect 253940 146208 253992 146260
rect 357440 146208 357492 146260
rect 358728 146208 358780 146260
rect 510620 146208 510672 146260
rect 54208 146140 54260 146192
rect 56324 146140 56376 146192
rect 58716 146140 58768 146192
rect 59636 146140 59688 146192
rect 53288 146004 53340 146056
rect 85580 146140 85632 146192
rect 179696 146140 179748 146192
rect 197452 146140 197504 146192
rect 219808 146140 219860 146192
rect 60924 146072 60976 146124
rect 86960 146072 87012 146124
rect 235264 146140 235316 146192
rect 255412 146140 255464 146192
rect 338488 146140 338540 146192
rect 357716 146140 357768 146192
rect 374460 146140 374512 146192
rect 375748 146140 375800 146192
rect 375932 146140 375984 146192
rect 376300 146140 376352 146192
rect 378876 146140 378928 146192
rect 379244 146140 379296 146192
rect 396724 146140 396776 146192
rect 418160 146140 418212 146192
rect 498660 146140 498712 146192
rect 517612 146140 517664 146192
rect 518440 146140 518492 146192
rect 252560 146072 252612 146124
rect 340236 146072 340288 146124
rect 357624 146072 357676 146124
rect 379980 146072 380032 146124
rect 414020 146072 414072 146124
rect 499856 146072 499908 146124
rect 517520 146072 517572 146124
rect 517704 146072 517756 146124
rect 60096 146004 60148 146056
rect 89812 146004 89864 146056
rect 216496 146004 216548 146056
rect 248420 146004 248472 146056
rect 375932 146004 375984 146056
rect 377956 146004 378008 146056
rect 378968 146004 379020 146056
rect 411260 146004 411312 146056
rect 54116 145936 54168 145988
rect 54760 145936 54812 145988
rect 84292 145936 84344 145988
rect 220084 145936 220136 145988
rect 251180 145936 251232 145988
rect 376300 145936 376352 145988
rect 407120 145936 407172 145988
rect 54300 145868 54352 145920
rect 54484 145868 54536 145920
rect 82820 145868 82872 145920
rect 219900 145868 219952 145920
rect 251272 145868 251324 145920
rect 377312 145868 377364 145920
rect 379060 145868 379112 145920
rect 409972 145868 410024 145920
rect 56416 145800 56468 145852
rect 84200 145800 84252 145852
rect 214380 145800 214432 145852
rect 215208 145800 215260 145852
rect 219164 145800 219216 145852
rect 249892 145800 249944 145852
rect 377956 145800 378008 145852
rect 408500 145800 408552 145852
rect 56324 145732 56376 145784
rect 88432 145732 88484 145784
rect 217232 145732 217284 145784
rect 245660 145732 245712 145784
rect 375748 145732 375800 145784
rect 402980 145732 403032 145784
rect 57520 145664 57572 145716
rect 91192 145664 91244 145716
rect 216220 145664 216272 145716
rect 242900 145664 242952 145716
rect 343548 145664 343600 145716
rect 356612 145664 356664 145716
rect 378876 145664 378928 145716
rect 403072 145664 403124 145716
rect 503628 145664 503680 145716
rect 517796 145664 517848 145716
rect 59636 145596 59688 145648
rect 93860 145596 93912 145648
rect 183468 145596 183520 145648
rect 197452 145596 197504 145648
rect 218520 145596 218572 145648
rect 244372 145596 244424 145648
rect 280068 145596 280120 145648
rect 356704 145596 356756 145648
rect 358820 145596 358872 145648
rect 378784 145596 378836 145648
rect 405740 145596 405792 145648
rect 517520 145596 517572 145648
rect 580264 145596 580316 145648
rect 58624 145528 58676 145580
rect 100760 145528 100812 145580
rect 191748 145528 191800 145580
rect 198004 145528 198056 145580
rect 214564 145528 214616 145580
rect 216496 145528 216548 145580
rect 244280 145528 244332 145580
rect 351644 145528 351696 145580
rect 358728 145528 358780 145580
rect 376576 145528 376628 145580
rect 404360 145528 404412 145580
rect 518440 145528 518492 145580
rect 580356 145528 580408 145580
rect 51908 145460 51960 145512
rect 77300 145460 77352 145512
rect 214288 145460 214340 145512
rect 236000 145460 236052 145512
rect 371700 145460 371752 145512
rect 373448 145460 373500 145512
rect 397460 145460 397512 145512
rect 48044 145392 48096 145444
rect 54668 145392 54720 145444
rect 76012 145392 76064 145444
rect 215668 145392 215720 145444
rect 236092 145392 236144 145444
rect 378600 145392 378652 145444
rect 396172 145392 396224 145444
rect 46480 145324 46532 145376
rect 54852 145324 54904 145376
rect 75920 145324 75972 145376
rect 215208 145324 215260 145376
rect 247132 145324 247184 145376
rect 378692 145324 378744 145376
rect 396080 145324 396132 145376
rect 56232 145256 56284 145308
rect 60924 145256 60976 145308
rect 377036 145256 377088 145308
rect 411352 145256 411404 145308
rect 217140 145052 217192 145104
rect 220084 145052 220136 145104
rect 218612 144984 218664 145036
rect 219808 144984 219860 145036
rect 218888 144916 218940 144968
rect 219900 144916 219952 144968
rect 51724 144848 51776 144900
rect 55956 144848 56008 144900
rect 56416 144848 56468 144900
rect 210792 144848 210844 144900
rect 211804 144848 211856 144900
rect 213552 144848 213604 144900
rect 218520 144848 218572 144900
rect 373632 144848 373684 144900
rect 378784 144848 378836 144900
rect 50528 144780 50580 144832
rect 55864 144780 55916 144832
rect 56508 144780 56560 144832
rect 213000 144780 213052 144832
rect 215944 144780 215996 144832
rect 216404 144780 216456 144832
rect 373724 144780 373776 144832
rect 376116 144780 376168 144832
rect 376576 144780 376628 144832
rect 51632 144712 51684 144764
rect 58624 144712 58676 144764
rect 212264 144712 212316 144764
rect 216036 144712 216088 144764
rect 216496 144712 216548 144764
rect 48136 144644 48188 144696
rect 56968 144644 57020 144696
rect 57520 144644 57572 144696
rect 48228 144576 48280 144628
rect 58716 144576 58768 144628
rect 215668 143692 215720 143744
rect 216496 143692 216548 143744
rect 55680 96568 55732 96620
rect 57060 96568 57112 96620
rect 215852 96568 215904 96620
rect 217508 96568 217560 96620
rect 520188 79976 520240 80028
rect 580448 79976 580500 80028
rect 41328 70320 41380 70372
rect 57520 70320 57572 70372
rect 370504 70320 370556 70372
rect 376944 70320 376996 70372
rect 214564 68960 214616 69012
rect 215208 68960 215260 69012
rect 213276 68892 213328 68944
rect 216772 68892 216824 68944
rect 215208 68348 215260 68400
rect 216680 68348 216732 68400
rect 358728 68280 358780 68332
rect 376944 68280 376996 68332
rect 358084 68144 358136 68196
rect 358728 68144 358780 68196
rect 214748 61956 214800 62008
rect 214932 61956 214984 62008
rect 378968 60664 379020 60716
rect 379244 60664 379296 60716
rect 54668 59780 54720 59832
rect 77116 59780 77168 59832
rect 55956 59712 56008 59764
rect 84200 59712 84252 59764
rect 378692 59712 378744 59764
rect 396080 59712 396132 59764
rect 55864 59644 55916 59696
rect 100760 59644 100812 59696
rect 217968 59644 218020 59696
rect 255872 59644 255924 59696
rect 378600 59644 378652 59696
rect 397092 59644 397144 59696
rect 54484 59576 54536 59628
rect 83096 59576 83148 59628
rect 219072 59576 219124 59628
rect 263876 59576 263928 59628
rect 378876 59576 378928 59628
rect 403072 59576 403124 59628
rect 54576 59508 54628 59560
rect 99472 59508 99524 59560
rect 216128 59508 216180 59560
rect 261760 59508 261812 59560
rect 378048 59508 378100 59560
rect 415860 59508 415912 59560
rect 56048 59440 56100 59492
rect 102784 59440 102836 59492
rect 214656 59440 214708 59492
rect 260656 59440 260708 59492
rect 376668 59440 376720 59492
rect 419448 59440 419500 59492
rect 58808 59372 58860 59424
rect 107568 59372 107620 59424
rect 215760 59372 215812 59424
rect 262864 59372 262916 59424
rect 360936 59372 360988 59424
rect 413560 59372 413612 59424
rect 54760 59304 54812 59356
rect 85396 59304 85448 59356
rect 214748 59304 214800 59356
rect 215208 59304 215260 59356
rect 358084 59304 358136 59356
rect 373448 59304 373500 59356
rect 398196 59304 398248 59356
rect 59084 59236 59136 59288
rect 95884 59236 95936 59288
rect 374644 59236 374696 59288
rect 410708 59236 410760 59288
rect 55036 59168 55088 59220
rect 98092 59168 98144 59220
rect 219440 59168 219492 59220
rect 256976 59168 257028 59220
rect 379152 59168 379204 59220
rect 416964 59168 417016 59220
rect 59820 59100 59872 59152
rect 106372 59100 106424 59152
rect 214932 59100 214984 59152
rect 259460 59100 259512 59152
rect 379612 59100 379664 59152
rect 418160 59100 418212 59152
rect 56140 59032 56192 59084
rect 103888 59032 103940 59084
rect 213828 59032 213880 59084
rect 298468 59032 298520 59084
rect 379704 59032 379756 59084
rect 425244 59032 425296 59084
rect 57336 58964 57388 59016
rect 105268 58964 105320 59016
rect 198556 58964 198608 59016
rect 295892 58964 295944 59016
rect 374368 58964 374420 59016
rect 421748 58964 421800 59016
rect 53196 58896 53248 58948
rect 114376 58896 114428 58948
rect 209044 58896 209096 58948
rect 308496 58896 308548 58948
rect 358176 58896 358228 58948
rect 423496 58896 423548 58948
rect 55588 58828 55640 58880
rect 138388 58828 138440 58880
rect 201408 58828 201460 58880
rect 303436 58828 303488 58880
rect 363696 58828 363748 58880
rect 468484 58828 468536 58880
rect 52184 58760 52236 58812
rect 143540 58760 143592 58812
rect 219348 58760 219400 58812
rect 425980 58760 426032 58812
rect 55496 58692 55548 58744
rect 150900 58692 150952 58744
rect 219624 58692 219676 58744
rect 421012 58692 421064 58744
rect 50068 58624 50120 58676
rect 148508 58624 148560 58676
rect 219072 58624 219124 58676
rect 428188 58624 428240 58676
rect 219348 57944 219400 57996
rect 430948 57944 431000 57996
rect 57244 57876 57296 57928
rect 57888 57876 57940 57928
rect 214748 57876 214800 57928
rect 343180 57876 343232 57928
rect 357532 57876 357584 57928
rect 361488 57876 361540 57928
rect 475844 57876 475896 57928
rect 503352 57876 503404 57928
rect 517796 57876 517848 57928
rect 53748 57808 53800 57860
rect 145564 57808 145616 57860
rect 183468 57808 183520 57860
rect 197452 57808 197504 57860
rect 209688 57808 209740 57860
rect 325884 57808 325936 57860
rect 343456 57808 343508 57860
rect 356612 57808 356664 57860
rect 373908 57808 373960 57860
rect 480628 57808 480680 57860
rect 503260 57808 503312 57860
rect 517888 57808 517940 57860
rect 53656 57740 53708 57792
rect 130844 57740 130896 57792
rect 183192 57740 183244 57792
rect 197360 57740 197412 57792
rect 215024 57740 215076 57792
rect 313372 57740 313424 57792
rect 378968 57740 379020 57792
rect 483388 57740 483440 57792
rect 49608 57672 49660 57724
rect 120724 57672 120776 57724
rect 212448 57672 212500 57724
rect 310980 57672 311032 57724
rect 364984 57672 365036 57724
rect 465908 57672 465960 57724
rect 49516 57604 49568 57656
rect 113548 57604 113600 57656
rect 218980 57604 219032 57656
rect 305828 57604 305880 57656
rect 366456 57604 366508 57656
rect 460940 57604 460992 57656
rect 57060 57536 57112 57588
rect 117964 57536 118016 57588
rect 216588 57536 216640 57588
rect 300860 57536 300912 57588
rect 379428 57536 379480 57588
rect 470876 57536 470928 57588
rect 59912 57468 59964 57520
rect 108580 57468 108632 57520
rect 211068 57468 211120 57520
rect 293316 57468 293368 57520
rect 362224 57468 362276 57520
rect 433524 57468 433576 57520
rect 60004 57400 60056 57452
rect 98460 57400 98512 57452
rect 213184 57400 213236 57452
rect 268200 57400 268252 57452
rect 279056 57400 279108 57452
rect 356704 57400 356756 57452
rect 367744 57400 367796 57452
rect 438492 57400 438544 57452
rect 51540 57332 51592 57384
rect 88432 57332 88484 57384
rect 215116 57332 215168 57384
rect 287612 57332 287664 57384
rect 374736 57332 374788 57384
rect 435916 57332 435968 57384
rect 59176 57264 59228 57316
rect 93676 57264 93728 57316
rect 218796 57264 218848 57316
rect 263600 57264 263652 57316
rect 373264 57264 373316 57316
rect 418436 57264 418488 57316
rect 59268 57196 59320 57248
rect 90732 57196 90784 57248
rect 218704 57196 218756 57248
rect 248144 57196 248196 57248
rect 365076 57196 365128 57248
rect 408316 57196 408368 57248
rect 54852 57128 54904 57180
rect 76012 57128 76064 57180
rect 214104 57128 214156 57180
rect 318248 57128 318300 57180
rect 41236 56516 41288 56568
rect 123484 56516 123536 56568
rect 213092 56516 213144 56568
rect 275652 56516 275704 56568
rect 375012 56516 375064 56568
rect 435088 56516 435140 56568
rect 52276 56448 52328 56500
rect 111156 56448 111208 56500
rect 217508 56448 217560 56500
rect 278044 56448 278096 56500
rect 374552 56448 374604 56500
rect 433340 56448 433392 56500
rect 53012 56380 53064 56432
rect 109500 56380 109552 56432
rect 213736 56380 213788 56432
rect 273260 56380 273312 56432
rect 374276 56380 374328 56432
rect 430580 56380 430632 56432
rect 58624 56312 58676 56364
rect 101772 56312 101824 56364
rect 215944 56312 215996 56364
rect 271236 56312 271288 56364
rect 376392 56312 376444 56364
rect 429660 56312 429712 56364
rect 59728 56244 59780 56296
rect 94412 56244 94464 56296
rect 219992 56244 220044 56296
rect 268660 56244 268712 56296
rect 379796 56244 379848 56296
rect 427636 56244 427688 56296
rect 58716 56176 58768 56228
rect 92204 56176 92256 56228
rect 219532 56176 219584 56228
rect 266360 56176 266412 56228
rect 376208 56176 376260 56228
rect 422852 56176 422904 56228
rect 53288 56108 53340 56160
rect 86500 56108 86552 56160
rect 217140 56108 217192 56160
rect 251180 56108 251232 56160
rect 379980 56108 380032 56160
rect 414572 56108 414624 56160
rect 58900 56040 58952 56092
rect 89996 56040 90048 56092
rect 218612 56040 218664 56092
rect 253388 56040 253440 56092
rect 379336 56040 379388 56092
rect 413468 56040 413520 56092
rect 52000 55972 52052 56024
rect 80428 55972 80480 56024
rect 214380 55972 214432 56024
rect 247684 55972 247736 56024
rect 375932 55972 375984 56024
rect 408684 55972 408736 56024
rect 51908 55904 51960 55956
rect 78220 55904 78272 55956
rect 216036 55904 216088 55956
rect 245292 55904 245344 55956
rect 379244 55904 379296 55956
rect 411260 55904 411312 55956
rect 211804 55836 211856 55888
rect 238116 55836 238168 55888
rect 374460 55836 374512 55888
rect 404084 55836 404136 55888
rect 213644 55768 213696 55820
rect 240508 55768 240560 55820
rect 373356 55768 373408 55820
rect 400404 55768 400456 55820
rect 54944 55156 54996 55208
rect 114560 55156 114612 55208
rect 218520 55156 218572 55208
rect 244372 55156 244424 55208
rect 375840 55156 375892 55208
rect 436100 55156 436152 55208
rect 53564 55088 53616 55140
rect 111800 55088 111852 55140
rect 214288 55088 214340 55140
rect 236000 55088 236052 55140
rect 376484 55088 376536 55140
rect 433708 55088 433760 55140
rect 54392 55020 54444 55072
rect 113180 55020 113232 55072
rect 219256 55020 219308 55072
rect 266452 55020 266504 55072
rect 375196 55020 375248 55072
rect 431960 55020 432012 55072
rect 56968 54952 57020 55004
rect 91192 54952 91244 55004
rect 219716 54952 219768 55004
rect 253940 54952 253992 55004
rect 379060 54952 379112 55004
rect 426532 54952 426584 55004
rect 58992 54884 59044 54936
rect 92480 54884 92532 54936
rect 218888 54884 218940 54936
rect 251364 54884 251416 54936
rect 378416 54884 378468 54936
rect 423680 54884 423732 54936
rect 56324 54816 56376 54868
rect 88340 54816 88392 54868
rect 216404 54816 216456 54868
rect 248420 54816 248472 54868
rect 377220 54816 377272 54868
rect 411352 54816 411404 54868
rect 56232 54748 56284 54800
rect 86960 54748 87012 54800
rect 219164 54748 219216 54800
rect 249800 54748 249852 54800
rect 377312 54748 377364 54800
rect 409880 54748 409932 54800
rect 53380 54680 53432 54732
rect 81440 54680 81492 54732
rect 217232 54680 217284 54732
rect 245660 54680 245712 54732
rect 376300 54680 376352 54732
rect 407120 54680 407172 54732
rect 52092 54612 52144 54664
rect 78680 54612 78732 54664
rect 213368 54612 213420 54664
rect 241520 54612 241572 54664
rect 376116 54612 376168 54664
rect 404360 54612 404412 54664
rect 216312 54544 216364 54596
rect 242900 54544 242952 54596
rect 378784 54544 378836 54596
rect 405832 54544 405884 54596
rect 214840 54476 214892 54528
rect 271880 54476 271932 54528
rect 374920 54476 374972 54528
rect 401600 54476 401652 54528
rect 214196 54408 214248 54460
rect 269120 54408 269172 54460
rect 374828 54408 374880 54460
rect 398840 54408 398892 54460
rect 213460 54340 213512 54392
rect 238760 54340 238812 54392
rect 216496 54272 216548 54324
rect 236092 54272 236144 54324
rect 2780 20340 2832 20392
rect 4804 20340 4856 20392
rect 147128 3476 147180 3528
rect 363604 3476 363656 3528
rect 572 3408 624 3460
rect 57244 3408 57296 3460
rect 125876 3408 125928 3460
rect 366364 3408 366416 3460
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 643754 3464 684247
rect 18604 645992 18656 645998
rect 18604 645934 18656 645940
rect 3424 643748 3476 643754
rect 3424 643690 3476 643696
rect 3422 632088 3478 632097
rect 3422 632023 3478 632032
rect 3148 580984 3200 580990
rect 3148 580926 3200 580932
rect 3160 580009 3188 580926
rect 3146 580000 3202 580009
rect 3146 579935 3202 579944
rect 3436 576162 3464 632023
rect 3424 576156 3476 576162
rect 3424 576098 3476 576104
rect 4804 574796 4856 574802
rect 4804 574738 4856 574744
rect 3424 567248 3476 567254
rect 3424 567190 3476 567196
rect 2964 411256 3016 411262
rect 2964 411198 3016 411204
rect 2976 410553 3004 411198
rect 2962 410544 3018 410553
rect 2962 410479 3018 410488
rect 3332 358760 3384 358766
rect 3332 358702 3384 358708
rect 3344 358465 3372 358702
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3436 97617 3464 567190
rect 3516 553104 3568 553110
rect 3516 553046 3568 553052
rect 3528 514865 3556 553046
rect 3514 514856 3570 514865
rect 3514 514791 3570 514800
rect 3516 479528 3568 479534
rect 3516 479470 3568 479476
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 3528 58585 3556 479470
rect 3608 478168 3660 478174
rect 3608 478110 3660 478116
rect 3620 462641 3648 478110
rect 3606 462632 3662 462641
rect 3606 462567 3662 462576
rect 3514 58576 3570 58585
rect 3514 58511 3570 58520
rect 4816 20398 4844 574738
rect 15844 491972 15896 491978
rect 15844 491914 15896 491920
rect 15856 411262 15884 491914
rect 15844 411256 15896 411262
rect 15844 411198 15896 411204
rect 18616 358766 18644 645934
rect 40052 563038 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 59176 654832 59228 654838
rect 59176 654774 59228 654780
rect 55128 644700 55180 644706
rect 55128 644642 55180 644648
rect 54944 644632 54996 644638
rect 54944 644574 54996 644580
rect 54852 642388 54904 642394
rect 54852 642330 54904 642336
rect 40040 563032 40092 563038
rect 40040 562974 40092 562980
rect 54864 555966 54892 642330
rect 54956 556102 54984 644574
rect 55036 644564 55088 644570
rect 55036 644506 55088 644512
rect 54944 556096 54996 556102
rect 54944 556038 54996 556044
rect 55048 556034 55076 644506
rect 55036 556028 55088 556034
rect 55036 555970 55088 555976
rect 54852 555960 54904 555966
rect 54852 555902 54904 555908
rect 55140 555762 55168 644642
rect 56324 643408 56376 643414
rect 56324 643350 56376 643356
rect 55128 555756 55180 555762
rect 55128 555698 55180 555704
rect 56336 555422 56364 643350
rect 56508 643340 56560 643346
rect 56508 643282 56560 643288
rect 56416 643204 56468 643210
rect 56416 643146 56468 643152
rect 56428 555830 56456 643146
rect 56416 555824 56468 555830
rect 56416 555766 56468 555772
rect 56520 555626 56548 643282
rect 57888 641776 57940 641782
rect 57888 641718 57940 641724
rect 57702 640656 57758 640665
rect 57702 640591 57758 640600
rect 57610 631816 57666 631825
rect 57610 631751 57666 631760
rect 57518 613456 57574 613465
rect 57518 613391 57574 613400
rect 57426 607336 57482 607345
rect 57426 607271 57482 607280
rect 57334 601216 57390 601225
rect 57334 601151 57390 601160
rect 57242 591696 57298 591705
rect 57242 591631 57298 591640
rect 57150 585576 57206 585585
rect 57150 585511 57206 585520
rect 57058 582856 57114 582865
rect 57058 582791 57114 582800
rect 57072 567866 57100 582791
rect 57164 569226 57192 585511
rect 57256 576298 57284 591631
rect 57348 580650 57376 601151
rect 57440 581262 57468 607271
rect 57428 581256 57480 581262
rect 57428 581198 57480 581204
rect 57336 580644 57388 580650
rect 57336 580586 57388 580592
rect 57244 576292 57296 576298
rect 57244 576234 57296 576240
rect 57532 570722 57560 613391
rect 57624 579086 57652 631751
rect 57716 579154 57744 640591
rect 57794 634536 57850 634545
rect 57794 634471 57850 634480
rect 57704 579148 57756 579154
rect 57704 579090 57756 579096
rect 57612 579080 57664 579086
rect 57612 579022 57664 579028
rect 57520 570716 57572 570722
rect 57520 570658 57572 570664
rect 57152 569220 57204 569226
rect 57152 569162 57204 569168
rect 57060 567860 57112 567866
rect 57060 567802 57112 567808
rect 57808 562358 57836 634471
rect 57900 616185 57928 641718
rect 59082 637936 59138 637945
rect 59082 637871 59138 637880
rect 58898 628416 58954 628425
rect 58898 628351 58954 628360
rect 58530 625696 58586 625705
rect 58530 625631 58586 625640
rect 57886 616176 57942 616185
rect 57886 616111 57942 616120
rect 57796 562352 57848 562358
rect 57796 562294 57848 562300
rect 56508 555620 56560 555626
rect 56508 555562 56560 555568
rect 56324 555416 56376 555422
rect 56324 555358 56376 555364
rect 57900 523025 57928 616111
rect 58438 597816 58494 597825
rect 58438 597751 58494 597760
rect 58452 579222 58480 597751
rect 58440 579216 58492 579222
rect 58440 579158 58492 579164
rect 58544 558210 58572 625631
rect 58806 610056 58862 610065
rect 58806 609991 58862 610000
rect 58622 603936 58678 603945
rect 58622 603871 58678 603880
rect 58636 574938 58664 603871
rect 58714 588976 58770 588985
rect 58714 588911 58770 588920
rect 58624 574932 58676 574938
rect 58624 574874 58676 574880
rect 58728 559570 58756 588911
rect 58820 580718 58848 609991
rect 58808 580712 58860 580718
rect 58808 580654 58860 580660
rect 58912 577658 58940 628351
rect 58990 622296 59046 622305
rect 58990 622231 59046 622240
rect 58900 577652 58952 577658
rect 58900 577594 58952 577600
rect 59004 566506 59032 622231
rect 59096 573510 59124 637871
rect 59188 619585 59216 654774
rect 104912 653410 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 170324 700330 170352 703520
rect 235184 700398 235212 703520
rect 235172 700392 235224 700398
rect 235172 700334 235224 700340
rect 170312 700324 170364 700330
rect 170312 700266 170364 700272
rect 147312 683188 147364 683194
rect 147312 683130 147364 683136
rect 104900 653404 104952 653410
rect 104900 653346 104952 653352
rect 145472 645312 145524 645318
rect 145472 645254 145524 645260
rect 144920 645176 144972 645182
rect 144920 645118 144972 645124
rect 142804 645108 142856 645114
rect 142804 645050 142856 645056
rect 115388 645040 115440 645046
rect 115388 644982 115440 644988
rect 124588 645040 124640 645046
rect 124588 644982 124640 644988
rect 86408 644972 86460 644978
rect 86408 644914 86460 644920
rect 80612 644700 80664 644706
rect 80612 644642 80664 644648
rect 59360 644496 59412 644502
rect 59360 644438 59412 644444
rect 59268 643272 59320 643278
rect 59268 643214 59320 643220
rect 59174 619576 59230 619585
rect 59174 619511 59230 619520
rect 59174 595096 59230 595105
rect 59174 595031 59230 595040
rect 59188 579630 59216 595031
rect 59176 579624 59228 579630
rect 59176 579566 59228 579572
rect 59084 573504 59136 573510
rect 59084 573446 59136 573452
rect 58992 566500 59044 566506
rect 58992 566442 59044 566448
rect 58716 559564 58768 559570
rect 58716 559506 58768 559512
rect 58532 558204 58584 558210
rect 58532 558146 58584 558152
rect 59280 555694 59308 643214
rect 59372 557534 59400 644438
rect 71596 643408 71648 643414
rect 71596 643350 71648 643356
rect 65800 643340 65852 643346
rect 65800 643282 65852 643288
rect 65812 643076 65840 643282
rect 69296 643136 69348 643142
rect 69046 643084 69296 643090
rect 69046 643078 69348 643084
rect 69046 643062 69336 643078
rect 71608 643076 71636 643350
rect 74816 643272 74868 643278
rect 74816 643214 74868 643220
rect 74828 643076 74856 643214
rect 77392 643204 77444 643210
rect 77392 643146 77444 643152
rect 77404 643076 77432 643146
rect 80624 643076 80652 644642
rect 83188 643204 83240 643210
rect 83188 643146 83240 643152
rect 83200 643076 83228 643146
rect 86420 643076 86448 644914
rect 94780 644904 94832 644910
rect 94780 644846 94832 644852
rect 92204 644632 92256 644638
rect 92204 644574 92256 644580
rect 88984 644564 89036 644570
rect 88984 644506 89036 644512
rect 88996 643076 89024 644506
rect 92216 643076 92244 644574
rect 94792 643076 94820 644846
rect 106372 644836 106424 644842
rect 106372 644778 106424 644784
rect 103796 644700 103848 644706
rect 103796 644642 103848 644648
rect 100576 644632 100628 644638
rect 100576 644574 100628 644580
rect 98000 644496 98052 644502
rect 98000 644438 98052 644444
rect 98012 643076 98040 644438
rect 100588 643076 100616 644574
rect 103808 643076 103836 644642
rect 106384 643076 106412 644778
rect 109592 644768 109644 644774
rect 109592 644710 109644 644716
rect 109604 643076 109632 644710
rect 112168 644564 112220 644570
rect 112168 644506 112220 644512
rect 112180 643076 112208 644506
rect 115400 643076 115428 644982
rect 124220 644972 124272 644978
rect 124220 644914 124272 644920
rect 120908 644904 120960 644910
rect 120908 644846 120960 644852
rect 117964 644496 118016 644502
rect 117964 644438 118016 644444
rect 117976 643076 118004 644438
rect 59464 642382 60030 642410
rect 62960 642394 63250 642410
rect 62948 642388 63250 642394
rect 59464 573442 59492 642382
rect 63000 642382 63250 642388
rect 120566 642382 120764 642410
rect 62948 642330 63000 642336
rect 120736 581806 120764 642382
rect 120814 618352 120870 618361
rect 120814 618287 120870 618296
rect 120724 581800 120776 581806
rect 120724 581742 120776 581748
rect 120722 581632 120778 581641
rect 120722 581567 120778 581576
rect 59912 581256 59964 581262
rect 59912 581198 59964 581204
rect 59924 576854 59952 581198
rect 60924 580712 60976 580718
rect 60924 580654 60976 580660
rect 119344 580712 119396 580718
rect 119344 580654 119396 580660
rect 60030 580094 60320 580122
rect 60292 577726 60320 580094
rect 60280 577720 60332 577726
rect 60280 577662 60332 577668
rect 59924 576826 60412 576854
rect 59452 573436 59504 573442
rect 59452 573378 59504 573384
rect 59372 557506 60320 557534
rect 59268 555688 59320 555694
rect 59268 555630 59320 555636
rect 60292 552976 60320 557506
rect 60384 555898 60412 576826
rect 60372 555892 60424 555898
rect 60372 555834 60424 555840
rect 60936 552976 60964 580654
rect 61384 580644 61436 580650
rect 61384 580586 61436 580592
rect 61396 555354 61424 580586
rect 112536 580304 112588 580310
rect 112536 580246 112588 580252
rect 62224 580094 62606 580122
rect 64984 580094 65182 580122
rect 68402 580094 68784 580122
rect 70978 580094 71360 580122
rect 62224 563786 62252 580094
rect 62396 579624 62448 579630
rect 62396 579566 62448 579572
rect 62212 563780 62264 563786
rect 62212 563722 62264 563728
rect 61660 555552 61712 555558
rect 61660 555494 61712 555500
rect 61384 555348 61436 555354
rect 61384 555290 61436 555296
rect 61672 552976 61700 555494
rect 62408 552976 62436 579566
rect 63776 578944 63828 578950
rect 63776 578886 63828 578892
rect 63132 560992 63184 560998
rect 63132 560934 63184 560940
rect 63144 552976 63172 560934
rect 63788 552976 63816 578886
rect 64984 576910 65012 580094
rect 66720 579012 66772 579018
rect 66720 578954 66772 578960
rect 64144 576904 64196 576910
rect 64144 576846 64196 576852
rect 64972 576904 65024 576910
rect 64972 576846 65024 576852
rect 64156 555558 64184 576846
rect 65248 576224 65300 576230
rect 65248 576166 65300 576172
rect 64512 573368 64564 573374
rect 64512 573310 64564 573316
rect 64144 555552 64196 555558
rect 64144 555494 64196 555500
rect 64524 552976 64552 573310
rect 65260 552976 65288 576166
rect 65984 572008 66036 572014
rect 65984 571950 66036 571956
rect 65996 552976 66024 571950
rect 66732 552976 66760 578954
rect 68756 577590 68784 580094
rect 68836 579216 68888 579222
rect 68836 579158 68888 579164
rect 68744 577584 68796 577590
rect 68744 577526 68796 577532
rect 68100 572280 68152 572286
rect 68100 572222 68152 572228
rect 67364 556096 67416 556102
rect 67364 556038 67416 556044
rect 67376 552976 67404 556038
rect 68112 552976 68140 572222
rect 68848 552976 68876 579158
rect 71044 579148 71096 579154
rect 71044 579090 71096 579096
rect 70308 574864 70360 574870
rect 70308 574806 70360 574812
rect 69572 559632 69624 559638
rect 69572 559574 69624 559580
rect 69584 552976 69612 559574
rect 70320 552976 70348 574806
rect 70952 572076 71004 572082
rect 70952 572018 71004 572024
rect 70964 552976 70992 572018
rect 71056 556102 71084 579090
rect 71136 577720 71188 577726
rect 71136 577662 71188 577668
rect 71148 565146 71176 577662
rect 71332 577522 71360 580094
rect 73172 580094 74198 580122
rect 76774 580094 77064 580122
rect 71320 577516 71372 577522
rect 71320 577458 71372 577464
rect 71136 565140 71188 565146
rect 71136 565082 71188 565088
rect 71688 563712 71740 563718
rect 71688 563654 71740 563660
rect 71044 556096 71096 556102
rect 71044 556038 71096 556044
rect 71700 552976 71728 563654
rect 73172 555422 73200 580094
rect 77036 577794 77064 580094
rect 78692 580094 79994 580122
rect 81452 580094 82570 580122
rect 85790 580094 86080 580122
rect 88366 580094 88472 580122
rect 77024 577788 77076 577794
rect 77024 577730 77076 577736
rect 75276 577720 75328 577726
rect 75276 577662 75328 577668
rect 74540 577652 74592 577658
rect 74540 577594 74592 577600
rect 73252 559700 73304 559706
rect 73252 559642 73304 559648
rect 72424 555416 72476 555422
rect 72424 555358 72476 555364
rect 73160 555416 73212 555422
rect 73160 555358 73212 555364
rect 72436 552976 72464 555358
rect 73264 553194 73292 559642
rect 73804 555552 73856 555558
rect 73804 555494 73856 555500
rect 73188 553166 73292 553194
rect 73188 552976 73216 553166
rect 73816 552976 73844 555494
rect 74552 552976 74580 577594
rect 75288 552976 75316 577662
rect 76012 573436 76064 573442
rect 76012 573378 76064 573384
rect 76024 552976 76052 573378
rect 78692 567934 78720 580094
rect 79324 576292 79376 576298
rect 79324 576234 79376 576240
rect 78864 570648 78916 570654
rect 78864 570590 78916 570596
rect 78680 567928 78732 567934
rect 78680 567870 78732 567876
rect 76748 561060 76800 561066
rect 76748 561002 76800 561008
rect 76760 552976 76788 561002
rect 77392 556096 77444 556102
rect 77392 556038 77444 556044
rect 77404 552976 77432 556038
rect 78128 555552 78180 555558
rect 78128 555494 78180 555500
rect 78140 552976 78168 555494
rect 78876 552976 78904 570590
rect 79336 555286 79364 576234
rect 80336 573436 80388 573442
rect 80336 573378 80388 573384
rect 79600 556028 79652 556034
rect 79600 555970 79652 555976
rect 79324 555280 79376 555286
rect 79324 555222 79376 555228
rect 79612 552976 79640 555970
rect 80348 552976 80376 573378
rect 81452 569362 81480 580094
rect 83188 579080 83240 579086
rect 83188 579022 83240 579028
rect 84568 579080 84620 579086
rect 84568 579022 84620 579028
rect 81440 569356 81492 569362
rect 81440 569298 81492 569304
rect 80980 569288 81032 569294
rect 80980 569230 81032 569236
rect 80992 552976 81020 569230
rect 82452 563848 82504 563854
rect 82452 563790 82504 563796
rect 81716 555280 81768 555286
rect 81716 555222 81768 555228
rect 81728 552976 81756 555222
rect 82464 552976 82492 563790
rect 83200 552976 83228 579022
rect 83924 555824 83976 555830
rect 83924 555766 83976 555772
rect 83936 552976 83964 555766
rect 84580 552976 84608 579022
rect 86052 577658 86080 580094
rect 87420 579216 87472 579222
rect 87420 579158 87472 579164
rect 86776 577788 86828 577794
rect 86776 577730 86828 577736
rect 86040 577652 86092 577658
rect 86040 577594 86092 577600
rect 86040 566568 86092 566574
rect 86040 566510 86092 566516
rect 85304 555824 85356 555830
rect 85304 555766 85356 555772
rect 85316 552976 85344 555766
rect 86052 552976 86080 566510
rect 86788 552976 86816 577730
rect 87432 552976 87460 579158
rect 88156 579148 88208 579154
rect 88156 579090 88208 579096
rect 87604 570716 87656 570722
rect 87604 570658 87656 570664
rect 87616 555286 87644 570658
rect 87604 555280 87656 555286
rect 87604 555222 87656 555228
rect 88168 552976 88196 579090
rect 88444 567194 88472 580094
rect 91112 580094 91586 580122
rect 94162 580094 94544 580122
rect 91112 576298 91140 580094
rect 93952 579284 94004 579290
rect 93952 579226 94004 579232
rect 91100 576292 91152 576298
rect 91100 576234 91152 576240
rect 91008 574932 91060 574938
rect 91008 574874 91060 574880
rect 89628 570716 89680 570722
rect 89628 570658 89680 570664
rect 88352 567166 88472 567194
rect 88352 562426 88380 567166
rect 88340 562420 88392 562426
rect 88340 562362 88392 562368
rect 88892 555960 88944 555966
rect 88892 555902 88944 555908
rect 88904 552976 88932 555902
rect 89640 552976 89668 570658
rect 90364 569356 90416 569362
rect 90364 569298 90416 569304
rect 90376 552976 90404 569298
rect 91020 552976 91048 574874
rect 92480 573504 92532 573510
rect 92480 573446 92532 573452
rect 91744 555280 91796 555286
rect 91744 555222 91796 555228
rect 91756 552976 91784 555222
rect 92492 552976 92520 573446
rect 93216 555756 93268 555762
rect 93216 555698 93268 555704
rect 93228 552976 93256 555698
rect 93964 552976 93992 579226
rect 94516 577794 94544 580094
rect 97000 580094 97382 580122
rect 99958 580094 100248 580122
rect 94504 577788 94556 577794
rect 94504 577730 94556 577736
rect 97000 577726 97028 580094
rect 97448 579420 97500 579426
rect 97448 579362 97500 579368
rect 96988 577720 97040 577726
rect 96988 577662 97040 577668
rect 96804 576292 96856 576298
rect 96804 576234 96856 576240
rect 94596 556844 94648 556850
rect 94596 556786 94648 556792
rect 94608 552976 94636 556786
rect 95332 555892 95384 555898
rect 95332 555834 95384 555840
rect 95344 552976 95372 555834
rect 96068 555280 96120 555286
rect 96068 555222 96120 555228
rect 96080 552976 96108 555222
rect 96816 552976 96844 576234
rect 97460 552976 97488 579362
rect 98184 579352 98236 579358
rect 98184 579294 98236 579300
rect 98196 552976 98224 579294
rect 100220 577726 100248 580094
rect 102152 580094 103178 580122
rect 104912 580094 105754 580122
rect 108592 580094 108974 580122
rect 110524 580094 111550 580122
rect 100208 577720 100260 577726
rect 100208 577662 100260 577668
rect 100392 576292 100444 576298
rect 100392 576234 100444 576240
rect 98644 569356 98696 569362
rect 98644 569298 98696 569304
rect 98656 555286 98684 569298
rect 99656 555688 99708 555694
rect 99656 555630 99708 555636
rect 98920 555620 98972 555626
rect 98920 555562 98972 555568
rect 98644 555280 98696 555286
rect 98644 555222 98696 555228
rect 98932 552976 98960 555562
rect 99668 552976 99696 555630
rect 100404 552976 100432 576234
rect 101036 567860 101088 567866
rect 101036 567802 101088 567808
rect 101048 552976 101076 567802
rect 102152 555234 102180 580094
rect 104164 577788 104216 577794
rect 104164 577730 104216 577736
rect 103244 569220 103296 569226
rect 103244 569162 103296 569168
rect 102508 566500 102560 566506
rect 102508 566442 102560 566448
rect 102060 555206 102180 555234
rect 102060 553194 102088 555206
rect 101800 553166 102088 553194
rect 101800 552976 101828 553166
rect 102520 552976 102548 566442
rect 103256 552976 103284 569162
rect 103980 555620 104032 555626
rect 103980 555562 104032 555568
rect 103992 552976 104020 555562
rect 104176 555286 104204 577730
rect 104912 570722 104940 580094
rect 107568 579488 107620 579494
rect 107568 579430 107620 579436
rect 106924 578196 106976 578202
rect 106924 578138 106976 578144
rect 105544 577584 105596 577590
rect 105544 577526 105596 577532
rect 104900 570716 104952 570722
rect 104900 570658 104952 570664
rect 105360 565140 105412 565146
rect 105360 565082 105412 565088
rect 104624 562420 104676 562426
rect 104624 562362 104676 562368
rect 104164 555280 104216 555286
rect 104164 555222 104216 555228
rect 104636 552976 104664 562362
rect 105372 552976 105400 565082
rect 105556 555218 105584 577526
rect 106936 559706 106964 578138
rect 106924 559700 106976 559706
rect 106924 559642 106976 559648
rect 106832 555688 106884 555694
rect 106832 555630 106884 555636
rect 106096 555280 106148 555286
rect 106096 555222 106148 555228
rect 105544 555212 105596 555218
rect 105544 555154 105596 555160
rect 106108 552976 106136 555222
rect 106844 552976 106872 555630
rect 107580 552976 107608 579430
rect 108592 578202 108620 580094
rect 108580 578196 108632 578202
rect 108580 578138 108632 578144
rect 108304 577652 108356 577658
rect 108304 577594 108356 577600
rect 108212 558204 108264 558210
rect 108212 558146 108264 558152
rect 108224 552976 108252 558146
rect 108316 555286 108344 577594
rect 108396 577516 108448 577522
rect 108396 577458 108448 577464
rect 110420 577516 110472 577522
rect 110420 577458 110472 577464
rect 108408 556102 108436 577458
rect 109684 563780 109736 563786
rect 109684 563722 109736 563728
rect 108396 556096 108448 556102
rect 108396 556038 108448 556044
rect 108304 555280 108356 555286
rect 108304 555222 108356 555228
rect 108948 555212 109000 555218
rect 108948 555154 109000 555160
rect 108960 552976 108988 555154
rect 109696 552976 109724 563722
rect 110432 552976 110460 577458
rect 110524 560998 110552 580094
rect 110512 560992 110564 560998
rect 110512 560934 110564 560940
rect 111064 559564 111116 559570
rect 111064 559506 111116 559512
rect 111076 552976 111104 559506
rect 111800 555280 111852 555286
rect 111800 555222 111852 555228
rect 111812 552976 111840 555222
rect 112548 552976 112576 580246
rect 114572 580094 114770 580122
rect 117346 580094 117452 580122
rect 114572 559638 114600 580094
rect 117424 578202 117452 580094
rect 116584 578196 116636 578202
rect 116584 578138 116636 578144
rect 117412 578196 117464 578202
rect 117412 578138 117464 578144
rect 115204 577720 115256 577726
rect 115204 577662 115256 577668
rect 114560 559632 114612 559638
rect 114560 559574 114612 559580
rect 114652 556096 114704 556102
rect 114652 556038 114704 556044
rect 114008 555756 114060 555762
rect 114008 555698 114060 555704
rect 113272 555416 113324 555422
rect 113272 555358 113324 555364
rect 113284 552976 113312 555358
rect 114020 552976 114048 555698
rect 114664 552976 114692 556038
rect 115216 555286 115244 577662
rect 115388 567928 115440 567934
rect 115388 567870 115440 567876
rect 115204 555280 115256 555286
rect 115204 555222 115256 555228
rect 115400 552976 115428 567870
rect 116596 561066 116624 578138
rect 116676 577652 116728 577658
rect 116676 577594 116728 577600
rect 116688 563854 116716 577594
rect 116676 563848 116728 563854
rect 116676 563790 116728 563796
rect 116676 562352 116728 562358
rect 116676 562294 116728 562300
rect 116584 561060 116636 561066
rect 116584 561002 116636 561008
rect 116688 555286 116716 562294
rect 118240 555892 118292 555898
rect 118240 555834 118292 555840
rect 116860 555484 116912 555490
rect 116860 555426 116912 555432
rect 116124 555280 116176 555286
rect 116124 555222 116176 555228
rect 116676 555280 116728 555286
rect 116676 555222 116728 555228
rect 116136 552976 116164 555222
rect 116872 552976 116900 555426
rect 117596 555280 117648 555286
rect 117596 555222 117648 555228
rect 117608 552976 117636 555222
rect 118252 552976 118280 555834
rect 118976 555484 119028 555490
rect 118976 555426 119028 555432
rect 118988 552976 119016 555426
rect 119356 555422 119384 580654
rect 120184 580094 120566 580122
rect 120184 577658 120212 580094
rect 120736 579018 120764 581567
rect 120724 579012 120776 579018
rect 120724 578954 120776 578960
rect 120172 577652 120224 577658
rect 120172 577594 120224 577600
rect 120828 573442 120856 618287
rect 120816 573436 120868 573442
rect 120816 573378 120868 573384
rect 119712 570716 119764 570722
rect 119712 570658 119764 570664
rect 119344 555416 119396 555422
rect 119344 555358 119396 555364
rect 119724 552976 119752 570658
rect 120448 559632 120500 559638
rect 120448 559574 120500 559580
rect 120460 552976 120488 559574
rect 120920 555830 120948 644846
rect 121644 644836 121696 644842
rect 121644 644778 121696 644784
rect 121460 644700 121512 644706
rect 121460 644642 121512 644648
rect 121000 644564 121052 644570
rect 121000 644506 121052 644512
rect 121012 579426 121040 644506
rect 121090 603256 121146 603265
rect 121090 603191 121146 603200
rect 121000 579420 121052 579426
rect 121000 579362 121052 579368
rect 121104 569294 121132 603191
rect 121184 581800 121236 581806
rect 121184 581742 121236 581748
rect 121196 577522 121224 581742
rect 121184 577516 121236 577522
rect 121184 577458 121236 577464
rect 121092 569288 121144 569294
rect 121092 569230 121144 569236
rect 121092 561128 121144 561134
rect 121092 561070 121144 561076
rect 120908 555824 120960 555830
rect 120908 555766 120960 555772
rect 121104 552976 121132 561070
rect 121472 555558 121500 644642
rect 121550 633856 121606 633865
rect 121550 633791 121606 633800
rect 121564 566574 121592 633791
rect 121656 579222 121684 644778
rect 122840 643136 122892 643142
rect 122840 643078 122892 643084
rect 121826 631136 121882 631145
rect 121826 631071 121882 631080
rect 121734 627736 121790 627745
rect 121734 627671 121790 627680
rect 121644 579216 121696 579222
rect 121644 579158 121696 579164
rect 121552 566568 121604 566574
rect 121552 566510 121604 566516
rect 121748 563718 121776 627671
rect 121840 572286 121868 631071
rect 121918 621616 121974 621625
rect 121918 621551 121974 621560
rect 121828 572280 121880 572286
rect 121828 572222 121880 572228
rect 121828 572144 121880 572150
rect 121828 572086 121880 572092
rect 121736 563712 121788 563718
rect 121736 563654 121788 563660
rect 121460 555552 121512 555558
rect 121460 555494 121512 555500
rect 121840 552976 121868 572086
rect 121932 572082 121960 621551
rect 122010 606656 122066 606665
rect 122010 606591 122066 606600
rect 122024 576230 122052 606591
rect 122102 600536 122158 600545
rect 122102 600471 122158 600480
rect 122116 579086 122144 600471
rect 122194 597136 122250 597145
rect 122194 597071 122250 597080
rect 122104 579080 122156 579086
rect 122104 579022 122156 579028
rect 122012 576224 122064 576230
rect 122012 576166 122064 576172
rect 122208 574870 122236 597071
rect 122286 588296 122342 588305
rect 122286 588231 122342 588240
rect 122300 578950 122328 588231
rect 122288 578944 122340 578950
rect 122288 578886 122340 578892
rect 122564 576360 122616 576366
rect 122564 576302 122616 576308
rect 122196 574864 122248 574870
rect 122196 574806 122248 574812
rect 121920 572076 121972 572082
rect 121920 572018 121972 572024
rect 122576 552976 122604 576302
rect 122852 555762 122880 643078
rect 122930 639976 122986 639985
rect 122930 639911 122986 639920
rect 122944 573374 122972 639911
rect 123114 637256 123170 637265
rect 123114 637191 123170 637200
rect 123022 612776 123078 612785
rect 123022 612711 123078 612720
rect 122932 573368 122984 573374
rect 122932 573310 122984 573316
rect 123036 556850 123064 612711
rect 123128 585002 123156 637191
rect 123206 625016 123262 625025
rect 123206 624951 123262 624960
rect 123116 584996 123168 585002
rect 123116 584938 123168 584944
rect 123114 584896 123170 584905
rect 123114 584831 123170 584840
rect 123128 580718 123156 584831
rect 123116 580712 123168 580718
rect 123116 580654 123168 580660
rect 123116 579216 123168 579222
rect 123116 579158 123168 579164
rect 123128 567194 123156 579158
rect 123220 572014 123248 624951
rect 123390 615496 123446 615505
rect 123390 615431 123446 615440
rect 123298 594416 123354 594425
rect 123298 594351 123354 594360
rect 123312 576298 123340 594351
rect 123300 576292 123352 576298
rect 123300 576234 123352 576240
rect 123208 572008 123260 572014
rect 123208 571950 123260 571956
rect 123404 569362 123432 615431
rect 124034 609376 124090 609385
rect 124034 609311 124090 609320
rect 124048 608666 124076 609311
rect 124036 608660 124088 608666
rect 124036 608602 124088 608608
rect 123482 591016 123538 591025
rect 123482 590951 123538 590960
rect 123496 570654 123524 590951
rect 123576 584996 123628 585002
rect 123576 584938 123628 584944
rect 123588 580310 123616 584938
rect 123576 580304 123628 580310
rect 123576 580246 123628 580252
rect 123484 570648 123536 570654
rect 123484 570590 123536 570596
rect 123392 569356 123444 569362
rect 123392 569298 123444 569304
rect 124036 569220 124088 569226
rect 124036 569162 124088 569168
rect 123128 567166 123340 567194
rect 123024 556844 123076 556850
rect 123024 556786 123076 556792
rect 122840 555756 122892 555762
rect 122840 555698 122892 555704
rect 123312 552976 123340 567166
rect 124048 552976 124076 569162
rect 124232 555626 124260 644914
rect 124404 644632 124456 644638
rect 124404 644574 124456 644580
rect 124312 643204 124364 643210
rect 124312 643146 124364 643152
rect 124324 555694 124352 643146
rect 124416 579290 124444 644574
rect 124496 644496 124548 644502
rect 124496 644438 124548 644444
rect 124404 579284 124456 579290
rect 124404 579226 124456 579232
rect 124508 579154 124536 644438
rect 124600 579494 124628 644982
rect 126980 644768 127032 644774
rect 126980 644710 127032 644716
rect 126244 643544 126296 643550
rect 126244 643486 126296 643492
rect 125416 643204 125468 643210
rect 125416 643146 125468 643152
rect 124588 579488 124640 579494
rect 124588 579430 124640 579436
rect 124496 579148 124548 579154
rect 124496 579090 124548 579096
rect 124680 565208 124732 565214
rect 124680 565150 124732 565156
rect 124312 555688 124364 555694
rect 124312 555630 124364 555636
rect 124220 555620 124272 555626
rect 124220 555562 124272 555568
rect 124692 552976 124720 565150
rect 125428 552976 125456 643146
rect 126152 573436 126204 573442
rect 126152 573378 126204 573384
rect 126164 552976 126192 573378
rect 126256 555898 126284 643486
rect 126888 597576 126940 597582
rect 126888 597518 126940 597524
rect 126244 555892 126296 555898
rect 126244 555834 126296 555840
rect 126900 552976 126928 597518
rect 126992 579358 127020 644710
rect 134064 644496 134116 644502
rect 134064 644438 134116 644444
rect 132592 627972 132644 627978
rect 132592 627914 132644 627920
rect 129096 610020 129148 610026
rect 129096 609962 129148 609968
rect 126980 579352 127032 579358
rect 126980 579294 127032 579300
rect 128268 575000 128320 575006
rect 128268 574942 128320 574948
rect 127624 556844 127676 556850
rect 127624 556786 127676 556792
rect 127636 552976 127664 556786
rect 128280 552976 128308 574942
rect 129004 566636 129056 566642
rect 129004 566578 129056 566584
rect 129016 552976 129044 566578
rect 129108 555490 129136 609962
rect 130476 577652 130528 577658
rect 130476 577594 130528 577600
rect 129740 561060 129792 561066
rect 129740 561002 129792 561008
rect 129096 555484 129148 555490
rect 129096 555426 129148 555432
rect 129752 552976 129780 561002
rect 130488 552976 130516 577594
rect 131212 563780 131264 563786
rect 131212 563722 131264 563728
rect 131224 552976 131252 563722
rect 131856 558204 131908 558210
rect 131856 558146 131908 558152
rect 131868 552976 131896 558146
rect 132604 552976 132632 627914
rect 133328 577584 133380 577590
rect 133328 577526 133380 577532
rect 133340 552976 133368 577526
rect 134076 552976 134104 644438
rect 141884 643408 141936 643414
rect 141884 643350 141936 643356
rect 137652 643340 137704 643346
rect 137652 643282 137704 643288
rect 134708 577516 134760 577522
rect 134708 577458 134760 577464
rect 134720 552976 134748 577458
rect 136916 570784 136968 570790
rect 136916 570726 136968 570732
rect 135444 556232 135496 556238
rect 135444 556174 135496 556180
rect 135456 552976 135484 556174
rect 136180 556164 136232 556170
rect 136180 556106 136232 556112
rect 136192 552976 136220 556106
rect 136928 552976 136956 570726
rect 137664 552976 137692 643282
rect 140044 640348 140096 640354
rect 140044 640290 140096 640296
rect 139768 590708 139820 590714
rect 139768 590650 139820 590656
rect 139032 572212 139084 572218
rect 139032 572154 139084 572160
rect 138296 555552 138348 555558
rect 138296 555494 138348 555500
rect 138308 552976 138336 555494
rect 139044 552976 139072 572154
rect 139780 552976 139808 590650
rect 140056 556238 140084 640290
rect 141240 630692 141292 630698
rect 141240 630634 141292 630640
rect 140504 559564 140556 559570
rect 140504 559506 140556 559512
rect 140044 556232 140096 556238
rect 140044 556174 140096 556180
rect 140516 552976 140544 559506
rect 141252 552976 141280 630634
rect 141896 552976 141924 643350
rect 142620 563848 142672 563854
rect 142620 563790 142672 563796
rect 142632 552976 142660 563790
rect 142816 558210 142844 645050
rect 143356 644836 143408 644842
rect 143356 644778 143408 644784
rect 142804 558204 142856 558210
rect 142804 558146 142856 558152
rect 143368 552976 143396 644778
rect 144184 643272 144236 643278
rect 144184 643214 144236 643220
rect 144196 556170 144224 643214
rect 144276 594856 144328 594862
rect 144276 594798 144328 594804
rect 144288 559638 144316 594798
rect 144276 559632 144328 559638
rect 144276 559574 144328 559580
rect 144736 558204 144788 558210
rect 144736 558146 144788 558152
rect 144184 556164 144236 556170
rect 144184 556106 144236 556112
rect 144092 555484 144144 555490
rect 144092 555426 144144 555432
rect 144104 552976 144132 555426
rect 144748 552976 144776 558146
rect 144932 555286 144960 645118
rect 144920 555280 144972 555286
rect 144920 555222 144972 555228
rect 145484 552976 145512 645254
rect 146116 643136 146168 643142
rect 146116 643078 146168 643084
rect 145564 608660 145616 608666
rect 145564 608602 145616 608608
rect 145576 580922 145604 608602
rect 145564 580916 145616 580922
rect 145564 580858 145616 580864
rect 146128 555762 146156 643078
rect 146208 641776 146260 641782
rect 146208 641718 146260 641724
rect 146220 616185 146248 641718
rect 146298 640656 146354 640665
rect 146298 640591 146354 640600
rect 146312 640354 146340 640591
rect 146300 640348 146352 640354
rect 146300 640290 146352 640296
rect 146298 631816 146354 631825
rect 146298 631751 146354 631760
rect 146312 630698 146340 631751
rect 146300 630692 146352 630698
rect 146300 630634 146352 630640
rect 146298 628416 146354 628425
rect 146298 628351 146354 628360
rect 146312 627978 146340 628351
rect 146300 627972 146352 627978
rect 146300 627914 146352 627920
rect 147218 625696 147274 625705
rect 147218 625631 147274 625640
rect 146206 616176 146262 616185
rect 146206 616111 146262 616120
rect 146298 610056 146354 610065
rect 146298 609991 146300 610000
rect 146352 609991 146354 610000
rect 146300 609962 146352 609968
rect 147126 607336 147182 607345
rect 147126 607271 147182 607280
rect 146298 597816 146354 597825
rect 146298 597751 146354 597760
rect 146312 597582 146340 597751
rect 146300 597576 146352 597582
rect 146300 597518 146352 597524
rect 146942 595096 146998 595105
rect 146942 595031 146998 595040
rect 146956 594862 146984 595031
rect 146944 594856 146996 594862
rect 146944 594798 146996 594804
rect 146298 591696 146354 591705
rect 146298 591631 146354 591640
rect 146312 590714 146340 591631
rect 146300 590708 146352 590714
rect 146300 590650 146352 590656
rect 147034 588976 147090 588985
rect 147034 588911 147090 588920
rect 147048 572014 147076 588911
rect 147140 580718 147168 607271
rect 147128 580712 147180 580718
rect 147128 580654 147180 580660
rect 147232 578882 147260 625631
rect 147324 619585 147352 683130
rect 299492 652050 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 307024 700392 307076 700398
rect 307024 700334 307076 700340
rect 299480 652044 299532 652050
rect 299480 651986 299532 651992
rect 235080 646536 235132 646542
rect 235080 646478 235132 646484
rect 234344 646264 234396 646270
rect 234344 646206 234396 646212
rect 147496 645380 147548 645386
rect 147496 645322 147548 645328
rect 164516 645380 164568 645386
rect 164516 645322 164568 645328
rect 147402 634536 147458 634545
rect 147402 634471 147458 634480
rect 147310 619576 147366 619585
rect 147310 619511 147366 619520
rect 147310 601216 147366 601225
rect 147310 601151 147366 601160
rect 147220 578876 147272 578882
rect 147220 578818 147272 578824
rect 147036 572008 147088 572014
rect 147036 571950 147088 571956
rect 147036 567928 147088 567934
rect 147036 567870 147088 567876
rect 146944 557184 146996 557190
rect 146944 557126 146996 557132
rect 146116 555756 146168 555762
rect 146116 555698 146168 555704
rect 146208 555280 146260 555286
rect 146208 555222 146260 555228
rect 146220 552976 146248 555222
rect 146956 552976 146984 557126
rect 147048 555558 147076 567870
rect 147324 562358 147352 601151
rect 147312 562352 147364 562358
rect 147312 562294 147364 562300
rect 147416 558278 147444 634471
rect 147404 558272 147456 558278
rect 147404 558214 147456 558220
rect 147508 555694 147536 645322
rect 156604 645176 156656 645182
rect 156656 645124 156736 645130
rect 156604 645118 156736 645124
rect 156616 645102 156736 645118
rect 156708 645046 156736 645102
rect 161480 645108 161532 645114
rect 161480 645050 161532 645056
rect 148784 645040 148836 645046
rect 156696 645040 156748 645046
rect 148784 644982 148836 644988
rect 147588 644904 147640 644910
rect 147588 644846 147640 644852
rect 147496 555688 147548 555694
rect 147496 555630 147548 555636
rect 147600 555558 147628 644846
rect 148416 644564 148468 644570
rect 148416 644506 148468 644512
rect 148230 603936 148286 603945
rect 148230 603871 148286 603880
rect 147680 557048 147732 557054
rect 147680 556990 147732 556996
rect 147036 555552 147088 555558
rect 147036 555494 147088 555500
rect 147588 555552 147640 555558
rect 147588 555494 147640 555500
rect 147692 552976 147720 556990
rect 148244 556238 148272 603871
rect 148324 583092 148376 583098
rect 148324 583034 148376 583040
rect 148336 579086 148364 583034
rect 148324 579080 148376 579086
rect 148324 579022 148376 579028
rect 148324 558340 148376 558346
rect 148324 558282 148376 558288
rect 148232 556232 148284 556238
rect 148232 556174 148284 556180
rect 148336 552976 148364 558282
rect 148428 557190 148456 644506
rect 148598 637936 148654 637945
rect 148598 637871 148654 637880
rect 148506 613456 148562 613465
rect 148506 613391 148562 613400
rect 148520 558890 148548 613391
rect 148612 579630 148640 637871
rect 148690 622296 148746 622305
rect 148690 622231 148746 622240
rect 148600 579624 148652 579630
rect 148600 579566 148652 579572
rect 148704 559638 148732 622231
rect 148796 583098 148824 644982
rect 156432 644978 156644 644994
rect 156696 644982 156748 644988
rect 148968 644972 149020 644978
rect 148968 644914 149020 644920
rect 156420 644972 156656 644978
rect 156472 644966 156604 644972
rect 156420 644914 156472 644920
rect 156604 644914 156656 644920
rect 148876 644632 148928 644638
rect 148876 644574 148928 644580
rect 148784 583092 148836 583098
rect 148784 583034 148836 583040
rect 148784 582956 148836 582962
rect 148784 582898 148836 582904
rect 148796 579018 148824 582898
rect 148888 579358 148916 644574
rect 148980 582962 149008 644914
rect 155224 644904 155276 644910
rect 155224 644846 155276 644852
rect 149704 644768 149756 644774
rect 149704 644710 149756 644716
rect 149058 585576 149114 585585
rect 149058 585511 149114 585520
rect 148968 582956 149020 582962
rect 148968 582898 149020 582904
rect 148966 582856 149022 582865
rect 148966 582791 149022 582800
rect 148876 579352 148928 579358
rect 148876 579294 148928 579300
rect 148980 579154 149008 582791
rect 148968 579148 149020 579154
rect 148968 579090 149020 579096
rect 148784 579012 148836 579018
rect 148784 578954 148836 578960
rect 149072 565146 149100 585511
rect 149716 578950 149744 644710
rect 149796 644700 149848 644706
rect 149796 644642 149848 644648
rect 149808 579290 149836 644642
rect 155236 644570 155264 644846
rect 153200 644564 153252 644570
rect 153200 644506 153252 644512
rect 155224 644564 155276 644570
rect 155224 644506 155276 644512
rect 158720 644564 158772 644570
rect 158720 644506 158772 644512
rect 149980 644496 150032 644502
rect 149980 644438 150032 644444
rect 149888 643476 149940 643482
rect 149888 643418 149940 643424
rect 149796 579284 149848 579290
rect 149796 579226 149848 579232
rect 149704 578944 149756 578950
rect 149704 578886 149756 578892
rect 149060 565140 149112 565146
rect 149060 565082 149112 565088
rect 148692 559632 148744 559638
rect 148692 559574 148744 559580
rect 148508 558884 148560 558890
rect 148508 558826 148560 558832
rect 149796 558884 149848 558890
rect 149796 558826 149848 558832
rect 148416 557184 148468 557190
rect 148416 557126 148468 557132
rect 149060 556232 149112 556238
rect 149060 556174 149112 556180
rect 149072 552976 149100 556174
rect 149808 552976 149836 558826
rect 149900 555286 149928 643418
rect 149992 643090 150020 644438
rect 153212 643090 153240 644506
rect 155500 643136 155552 643142
rect 149992 643062 150052 643090
rect 153212 643062 153272 643090
rect 158732 643090 158760 644506
rect 161492 643090 161520 645050
rect 164528 643090 164556 645322
rect 196072 645176 196124 645182
rect 196072 645118 196124 645124
rect 172888 644972 172940 644978
rect 172888 644914 172940 644920
rect 170312 643476 170364 643482
rect 170312 643418 170364 643424
rect 167092 643408 167144 643414
rect 167092 643350 167144 643356
rect 167104 643090 167132 643350
rect 170324 643090 170352 643418
rect 172900 643090 172928 644914
rect 176108 644904 176160 644910
rect 176108 644846 176160 644852
rect 176120 643090 176148 644846
rect 184480 644836 184532 644842
rect 184480 644778 184532 644784
rect 179006 643340 179058 643346
rect 179006 643282 179058 643288
rect 155552 643084 155848 643090
rect 155500 643078 155848 643084
rect 155512 643062 155848 643078
rect 158732 643062 159068 643090
rect 161492 643062 161644 643090
rect 164528 643062 164864 643090
rect 167104 643062 167440 643090
rect 170324 643062 170660 643090
rect 172900 643062 173236 643090
rect 176120 643062 176456 643090
rect 179018 643076 179046 643282
rect 182226 643204 182278 643210
rect 182226 643146 182278 643152
rect 182238 643076 182266 643146
rect 184492 643090 184520 644778
rect 190460 644768 190512 644774
rect 190460 644710 190512 644716
rect 187700 643544 187752 643550
rect 187700 643486 187752 643492
rect 187712 643090 187740 643486
rect 190472 643090 190500 644710
rect 193818 643272 193870 643278
rect 193818 643214 193870 643220
rect 184492 643062 184828 643090
rect 187712 643062 188048 643090
rect 190472 643062 190624 643090
rect 193830 643076 193858 643214
rect 196084 643090 196112 645118
rect 215024 645108 215076 645114
rect 215024 645050 215076 645056
rect 207664 645040 207716 645046
rect 207664 644982 207716 644988
rect 199292 644700 199344 644706
rect 199292 644642 199344 644648
rect 199304 643090 199332 644642
rect 201868 644564 201920 644570
rect 201868 644506 201920 644512
rect 201880 643090 201908 644506
rect 205548 644496 205600 644502
rect 205548 644438 205600 644444
rect 205560 643090 205588 644438
rect 196084 643062 196420 643090
rect 199304 643062 199640 643090
rect 201880 643062 202216 643090
rect 205436 643062 205588 643090
rect 207676 643090 207704 644982
rect 214288 644972 214340 644978
rect 214288 644914 214340 644920
rect 211160 644496 211212 644502
rect 211160 644438 211212 644444
rect 207676 643062 208012 643090
rect 210588 642382 210740 642410
rect 151084 580712 151136 580718
rect 151084 580654 151136 580660
rect 150052 580094 150388 580122
rect 150360 577794 150388 580094
rect 150532 579624 150584 579630
rect 150532 579566 150584 579572
rect 150348 577788 150400 577794
rect 150348 577730 150400 577736
rect 149888 555280 149940 555286
rect 149888 555222 149940 555228
rect 150544 552976 150572 579566
rect 151096 556102 151124 580654
rect 199384 580304 199436 580310
rect 199384 580246 199436 580252
rect 151924 580094 152628 580122
rect 154684 580094 155204 580122
rect 157352 580094 158424 580122
rect 160112 580094 161000 580122
rect 163884 580094 164220 580122
rect 165724 580094 166796 580122
rect 169772 580094 170016 580122
rect 172532 580094 172592 580122
rect 175476 580094 175812 580122
rect 178052 580094 178388 580122
rect 181272 580094 181608 580122
rect 183848 580094 184184 580122
rect 187068 580094 187404 580122
rect 189644 580094 189980 580122
rect 192864 580094 193200 580122
rect 195440 580094 195776 580122
rect 198752 580094 198996 580122
rect 151820 578944 151872 578950
rect 151820 578886 151872 578892
rect 151176 577788 151228 577794
rect 151176 577730 151228 577736
rect 151188 566574 151216 577730
rect 151176 566568 151228 566574
rect 151176 566510 151228 566516
rect 151832 557534 151860 578886
rect 151924 576854 151952 580094
rect 151924 576826 152044 576854
rect 151832 557506 151952 557534
rect 151084 556096 151136 556102
rect 151084 556038 151136 556044
rect 151268 555280 151320 555286
rect 151268 555222 151320 555228
rect 151280 552976 151308 555222
rect 151924 552976 151952 557506
rect 152016 555626 152044 576826
rect 154684 570722 154712 580094
rect 155500 579352 155552 579358
rect 155500 579294 155552 579300
rect 154856 577788 154908 577794
rect 154856 577730 154908 577736
rect 154672 570716 154724 570722
rect 154672 570658 154724 570664
rect 152648 565276 152700 565282
rect 152648 565218 152700 565224
rect 152004 555620 152056 555626
rect 152004 555562 152056 555568
rect 152660 552976 152688 565218
rect 153384 556096 153436 556102
rect 153384 556038 153436 556044
rect 153396 552976 153424 556038
rect 154120 555280 154172 555286
rect 154120 555222 154172 555228
rect 154132 552976 154160 555222
rect 154868 552976 154896 577730
rect 155512 552976 155540 579294
rect 156236 579284 156288 579290
rect 156236 579226 156288 579232
rect 156248 552976 156276 579226
rect 157352 555830 157380 580094
rect 159088 579148 159140 579154
rect 159088 579090 159140 579096
rect 158352 562420 158404 562426
rect 158352 562362 158404 562368
rect 157340 555824 157392 555830
rect 157340 555766 157392 555772
rect 156972 555756 157024 555762
rect 156972 555698 157024 555704
rect 156984 552976 157012 555698
rect 157708 555688 157760 555694
rect 157708 555630 157760 555636
rect 157720 552976 157748 555630
rect 158364 552976 158392 562362
rect 159100 552976 159128 579090
rect 159824 577720 159876 577726
rect 159824 577662 159876 577668
rect 159836 552976 159864 577662
rect 160112 566506 160140 580094
rect 161940 579080 161992 579086
rect 161940 579022 161992 579028
rect 160744 576428 160796 576434
rect 160744 576370 160796 576376
rect 160100 566500 160152 566506
rect 160100 566442 160152 566448
rect 160560 559632 160612 559638
rect 160560 559574 160612 559580
rect 160572 552976 160600 559574
rect 160756 555286 160784 576370
rect 161296 565140 161348 565146
rect 161296 565082 161348 565088
rect 160744 555280 160796 555286
rect 160744 555222 160796 555228
rect 161308 552976 161336 565082
rect 161952 552976 161980 579022
rect 162676 577924 162728 577930
rect 162676 577866 162728 577872
rect 162688 552976 162716 577866
rect 163884 577658 163912 580094
rect 165528 579284 165580 579290
rect 165528 579226 165580 579232
rect 164884 579012 164936 579018
rect 164884 578954 164936 578960
rect 164148 577856 164200 577862
rect 164148 577798 164200 577804
rect 163872 577652 163924 577658
rect 163872 577594 163924 577600
rect 163412 566568 163464 566574
rect 163412 566510 163464 566516
rect 163424 552976 163452 566510
rect 164160 552976 164188 577798
rect 164896 552976 164924 578954
rect 165540 552976 165568 579226
rect 165724 558210 165752 580094
rect 166264 578876 166316 578882
rect 166264 578818 166316 578824
rect 165712 558204 165764 558210
rect 165712 558146 165764 558152
rect 166276 552976 166304 578818
rect 169116 572008 169168 572014
rect 169116 571950 169168 571956
rect 168380 558204 168432 558210
rect 168380 558146 168432 558152
rect 167000 555824 167052 555830
rect 167000 555766 167052 555772
rect 167012 552976 167040 555766
rect 167736 555620 167788 555626
rect 167736 555562 167788 555568
rect 167748 552976 167776 555562
rect 168392 552976 168420 558146
rect 169128 552976 169156 571950
rect 169772 562306 169800 580094
rect 169852 577652 169904 577658
rect 169852 577594 169904 577600
rect 169864 562442 169892 577594
rect 169864 562414 170076 562442
rect 169772 562278 169984 562306
rect 169852 562216 169904 562222
rect 169852 562158 169904 562164
rect 169760 558272 169812 558278
rect 169760 558214 169812 558220
rect 169772 555694 169800 558214
rect 169760 555688 169812 555694
rect 169760 555630 169812 555636
rect 169864 552976 169892 562158
rect 169956 556170 169984 562278
rect 170048 562222 170076 562414
rect 170036 562216 170088 562222
rect 170036 562158 170088 562164
rect 172532 558346 172560 580094
rect 174176 577992 174228 577998
rect 174176 577934 174228 577940
rect 172704 566500 172756 566506
rect 172704 566442 172756 566448
rect 172520 558340 172572 558346
rect 172520 558282 172572 558288
rect 171324 558272 171376 558278
rect 171324 558214 171376 558220
rect 169944 556164 169996 556170
rect 169944 556106 169996 556112
rect 170588 555620 170640 555626
rect 170588 555562 170640 555568
rect 170600 552976 170628 555562
rect 171336 552976 171364 558214
rect 171968 555552 172020 555558
rect 171968 555494 172020 555500
rect 171980 552976 172008 555494
rect 172716 552976 172744 566442
rect 173440 556164 173492 556170
rect 173440 556106 173492 556112
rect 173452 552976 173480 556106
rect 174188 552976 174216 577934
rect 175476 577658 175504 580094
rect 178052 577930 178080 580094
rect 179880 578944 179932 578950
rect 179880 578886 179932 578892
rect 178040 577924 178092 577930
rect 178040 577866 178092 577872
rect 175464 577652 175516 577658
rect 175464 577594 175516 577600
rect 177028 573504 177080 573510
rect 177028 573446 177080 573452
rect 174912 562352 174964 562358
rect 174912 562294 174964 562300
rect 174924 552976 174952 562294
rect 176292 556980 176344 556986
rect 176292 556922 176344 556928
rect 175556 555688 175608 555694
rect 175556 555630 175608 555636
rect 175568 552976 175596 555630
rect 176304 552976 176332 556922
rect 177040 552976 177068 573446
rect 178500 569288 178552 569294
rect 178500 569230 178552 569236
rect 177764 566704 177816 566710
rect 177764 566646 177816 566652
rect 177776 552976 177804 566646
rect 178512 552976 178540 569230
rect 179144 565140 179196 565146
rect 179144 565082 179196 565088
rect 179156 552976 179184 565082
rect 179892 552976 179920 578886
rect 181272 577794 181300 580094
rect 183848 577862 183876 580094
rect 184204 579012 184256 579018
rect 184204 578954 184256 578960
rect 183836 577856 183888 577862
rect 183836 577798 183888 577804
rect 181260 577788 181312 577794
rect 181260 577730 181312 577736
rect 183468 577652 183520 577658
rect 183468 577594 183520 577600
rect 180616 576224 180668 576230
rect 180616 576166 180668 576172
rect 180628 552976 180656 576166
rect 181352 574864 181404 574870
rect 181352 574806 181404 574812
rect 181364 552976 181392 574806
rect 181996 573368 182048 573374
rect 181996 573310 182048 573316
rect 182008 552976 182036 573310
rect 182732 560992 182784 560998
rect 182732 560934 182784 560940
rect 182744 552976 182772 560934
rect 183480 552976 183508 577594
rect 184216 552976 184244 578954
rect 187068 577590 187096 580094
rect 189644 577998 189672 580094
rect 191104 578196 191156 578202
rect 191104 578138 191156 578144
rect 189632 577992 189684 577998
rect 189632 577934 189684 577940
rect 187056 577584 187108 577590
rect 187056 577526 187108 577532
rect 187792 574932 187844 574938
rect 187792 574874 187844 574880
rect 185584 570648 185636 570654
rect 185584 570590 185636 570596
rect 184940 559632 184992 559638
rect 184940 559574 184992 559580
rect 184952 552976 184980 559574
rect 185596 552976 185624 570590
rect 187056 563712 187108 563718
rect 187056 563654 187108 563660
rect 186320 555824 186372 555830
rect 186320 555766 186372 555772
rect 186332 552976 186360 555766
rect 187068 552976 187096 563654
rect 187804 552976 187832 574874
rect 189908 572280 189960 572286
rect 189908 572222 189960 572228
rect 189172 562352 189224 562358
rect 189172 562294 189224 562300
rect 188528 556912 188580 556918
rect 188528 556854 188580 556860
rect 188540 552976 188568 556854
rect 189184 552976 189212 562294
rect 189920 552976 189948 572222
rect 190644 558340 190696 558346
rect 190644 558282 190696 558288
rect 190656 552976 190684 558282
rect 191116 557054 191144 578138
rect 192484 578128 192536 578134
rect 192484 578070 192536 578076
rect 192116 570852 192168 570858
rect 192116 570794 192168 570800
rect 191380 566568 191432 566574
rect 191380 566510 191432 566516
rect 191104 557048 191156 557054
rect 191104 556990 191156 556996
rect 191392 552976 191420 566510
rect 192128 552976 192156 570794
rect 192496 563786 192524 578070
rect 192864 577726 192892 580094
rect 195440 578202 195468 580094
rect 196348 579080 196400 579086
rect 196348 579022 196400 579028
rect 195428 578196 195480 578202
rect 195428 578138 195480 578144
rect 192852 577720 192904 577726
rect 192852 577662 192904 577668
rect 195244 577584 195296 577590
rect 195244 577526 195296 577532
rect 194968 572008 195020 572014
rect 194968 571950 195020 571956
rect 193496 563916 193548 563922
rect 193496 563858 193548 563864
rect 192484 563780 192536 563786
rect 192484 563722 192536 563728
rect 192760 563780 192812 563786
rect 192760 563722 192812 563728
rect 192772 552976 192800 563722
rect 193508 552976 193536 563858
rect 194232 555688 194284 555694
rect 194232 555630 194284 555636
rect 194244 552976 194272 555630
rect 194980 552976 195008 571950
rect 195256 555490 195284 577526
rect 195612 555552 195664 555558
rect 195612 555494 195664 555500
rect 195244 555484 195296 555490
rect 195244 555426 195296 555432
rect 195624 552976 195652 555494
rect 196360 552976 196388 579022
rect 198752 578134 198780 580094
rect 198740 578128 198792 578134
rect 198740 578070 198792 578076
rect 198004 577720 198056 577726
rect 198004 577662 198056 577668
rect 197084 570716 197136 570722
rect 197084 570658 197136 570664
rect 197096 552976 197124 570658
rect 197820 559700 197872 559706
rect 197820 559642 197872 559648
rect 197832 552976 197860 559642
rect 198016 559570 198044 577662
rect 199200 567996 199252 568002
rect 199200 567938 199252 567944
rect 198556 566500 198608 566506
rect 198556 566442 198608 566448
rect 198004 559564 198056 559570
rect 198004 559506 198056 559512
rect 198568 552976 198596 566442
rect 199212 552976 199240 567938
rect 199396 555626 199424 580246
rect 201512 580094 201572 580122
rect 204456 580094 204792 580122
rect 207032 580094 207368 580122
rect 210252 580094 210588 580122
rect 200672 579148 200724 579154
rect 200672 579090 200724 579096
rect 199476 576904 199528 576910
rect 199476 576846 199528 576852
rect 199488 561134 199516 576846
rect 199476 561128 199528 561134
rect 199476 561070 199528 561076
rect 199936 555756 199988 555762
rect 199936 555698 199988 555704
rect 199384 555620 199436 555626
rect 199384 555562 199436 555568
rect 199948 552976 199976 555698
rect 200684 552976 200712 579090
rect 201512 576910 201540 580094
rect 204456 577250 204484 580094
rect 207032 577522 207060 580094
rect 210252 577726 210280 580094
rect 210240 577720 210292 577726
rect 210240 577662 210292 577668
rect 207020 577516 207072 577522
rect 207020 577458 207072 577464
rect 202236 577244 202288 577250
rect 202236 577186 202288 577192
rect 204444 577244 204496 577250
rect 204444 577186 204496 577192
rect 201500 576904 201552 576910
rect 201500 576846 201552 576852
rect 202144 559564 202196 559570
rect 202144 559506 202196 559512
rect 201408 555892 201460 555898
rect 201408 555834 201460 555840
rect 201420 552976 201448 555834
rect 202156 552976 202184 559506
rect 202248 556850 202276 577186
rect 206284 576292 206336 576298
rect 206284 576234 206336 576240
rect 204260 573572 204312 573578
rect 204260 573514 204312 573520
rect 202788 565344 202840 565350
rect 202788 565286 202840 565292
rect 202236 556844 202288 556850
rect 202236 556786 202288 556792
rect 202800 552976 202828 565286
rect 203524 555960 203576 555966
rect 203524 555902 203576 555908
rect 203536 552976 203564 555902
rect 204272 552976 204300 573514
rect 204996 569356 205048 569362
rect 204996 569298 205048 569304
rect 205008 552976 205036 569298
rect 205640 567860 205692 567866
rect 205640 567802 205692 567808
rect 205652 552976 205680 567802
rect 206296 555830 206324 576234
rect 209780 572076 209832 572082
rect 209780 572018 209832 572024
rect 207112 562488 207164 562494
rect 207112 562430 207164 562436
rect 206376 561128 206428 561134
rect 206376 561070 206428 561076
rect 206284 555824 206336 555830
rect 206284 555766 206336 555772
rect 206388 552976 206416 561070
rect 207124 552976 207152 562430
rect 208584 558408 208636 558414
rect 208584 558350 208636 558356
rect 207848 556844 207900 556850
rect 207848 556786 207900 556792
rect 207860 552976 207888 556786
rect 208596 552976 208624 558350
rect 209792 557534 209820 572018
rect 210712 558210 210740 642382
rect 210790 584352 210846 584361
rect 210790 584287 210846 584296
rect 210804 558278 210832 584287
rect 210882 581632 210938 581641
rect 210882 581567 210938 581576
rect 210896 565214 210924 581567
rect 211172 579290 211200 644438
rect 211250 639432 211306 639441
rect 211250 639367 211306 639376
rect 211160 579284 211212 579290
rect 211160 579226 211212 579232
rect 211264 576366 211292 639367
rect 212630 636712 212686 636721
rect 212630 636647 212686 636656
rect 211342 630728 211398 630737
rect 211342 630663 211398 630672
rect 211252 576360 211304 576366
rect 211252 576302 211304 576308
rect 211356 573442 211384 630663
rect 212538 627192 212594 627201
rect 212538 627127 212594 627136
rect 211526 624472 211582 624481
rect 211526 624407 211582 624416
rect 211434 621072 211490 621081
rect 211434 621007 211490 621016
rect 211344 573436 211396 573442
rect 211344 573378 211396 573384
rect 211448 566642 211476 621007
rect 211540 569226 211568 624407
rect 211710 606248 211766 606257
rect 211710 606183 211766 606192
rect 211618 600672 211674 600681
rect 211618 600607 211674 600616
rect 211528 569220 211580 569226
rect 211528 569162 211580 569168
rect 211436 566636 211488 566642
rect 211436 566578 211488 566584
rect 210884 565208 210936 565214
rect 210884 565150 210936 565156
rect 211632 563854 211660 600607
rect 211724 579222 211752 606183
rect 211802 596728 211858 596737
rect 211802 596663 211858 596672
rect 211712 579216 211764 579222
rect 211712 579158 211764 579164
rect 211816 575006 211844 596663
rect 211894 588024 211950 588033
rect 211894 587959 211950 587968
rect 211804 575000 211856 575006
rect 211804 574942 211856 574948
rect 211908 572150 211936 587959
rect 211896 572144 211948 572150
rect 211896 572086 211948 572092
rect 211620 563848 211672 563854
rect 211620 563790 211672 563796
rect 212552 561066 212580 627127
rect 212644 580310 212672 636647
rect 212722 633448 212778 633457
rect 212722 633383 212778 633392
rect 212632 580304 212684 580310
rect 212632 580246 212684 580252
rect 212736 577590 212764 633383
rect 212814 618352 212870 618361
rect 212814 618287 212870 618296
rect 212724 577584 212776 577590
rect 212724 577526 212776 577532
rect 212828 567934 212856 618287
rect 212998 614952 213054 614961
rect 212998 614887 213054 614896
rect 212906 612912 212962 612921
rect 212906 612847 212962 612856
rect 212816 567928 212868 567934
rect 212816 567870 212868 567876
rect 212920 565282 212948 612847
rect 213012 576434 213040 614887
rect 213826 608832 213882 608841
rect 213882 608790 213960 608818
rect 213826 608767 213882 608776
rect 213090 603392 213146 603401
rect 213090 603327 213146 603336
rect 213000 576428 213052 576434
rect 213000 576370 213052 576376
rect 213104 572218 213132 603327
rect 213274 593872 213330 593881
rect 213274 593807 213330 593816
rect 213182 590744 213238 590753
rect 213182 590679 213238 590688
rect 213092 572212 213144 572218
rect 213092 572154 213144 572160
rect 213196 570790 213224 590679
rect 213184 570784 213236 570790
rect 213184 570726 213236 570732
rect 212908 565276 212960 565282
rect 212908 565218 212960 565224
rect 213288 562426 213316 593807
rect 213932 580922 213960 608790
rect 213920 580916 213972 580922
rect 213920 580858 213972 580864
rect 213276 562420 213328 562426
rect 213276 562362 213328 562368
rect 212540 561060 212592 561066
rect 212540 561002 212592 561008
rect 210792 558272 210844 558278
rect 210792 558214 210844 558220
rect 212816 558272 212868 558278
rect 212816 558214 212868 558220
rect 210700 558204 210752 558210
rect 210700 558146 210752 558152
rect 212172 558204 212224 558210
rect 212172 558146 212224 558152
rect 209792 557506 210740 557534
rect 209228 555824 209280 555830
rect 209228 555766 209280 555772
rect 209240 552976 209268 555766
rect 209964 555620 210016 555626
rect 209964 555562 210016 555568
rect 209976 552976 210004 555562
rect 210712 552976 210740 557506
rect 211436 557048 211488 557054
rect 211436 556990 211488 556996
rect 211448 552976 211476 556990
rect 212184 552976 212212 558146
rect 212828 552976 212856 558214
rect 213552 555484 213604 555490
rect 213552 555426 213604 555432
rect 213564 552976 213592 555426
rect 214300 552976 214328 644914
rect 214564 641844 214616 641850
rect 214564 641786 214616 641792
rect 214576 555694 214604 641786
rect 214564 555688 214616 555694
rect 214564 555630 214616 555636
rect 215036 552976 215064 645050
rect 226432 645040 226484 645046
rect 226432 644982 226484 644988
rect 222936 644768 222988 644774
rect 222936 644710 222988 644716
rect 220084 643544 220136 643550
rect 220084 643486 220136 643492
rect 215944 643204 215996 643210
rect 215944 643146 215996 643152
rect 215760 638240 215812 638246
rect 215760 638182 215812 638188
rect 215772 552976 215800 638182
rect 215956 555898 215984 643146
rect 217324 643136 217376 643142
rect 217324 643078 217376 643084
rect 216036 594856 216088 594862
rect 216036 594798 216088 594804
rect 216048 569294 216076 594798
rect 217140 577516 217192 577522
rect 217140 577458 217192 577464
rect 216404 573436 216456 573442
rect 216404 573378 216456 573384
rect 216036 569288 216088 569294
rect 216036 569230 216088 569236
rect 215944 555892 215996 555898
rect 215944 555834 215996 555840
rect 216416 552976 216444 573378
rect 217152 552976 217180 577458
rect 217336 555966 217364 643078
rect 218612 621036 218664 621042
rect 218612 620978 218664 620984
rect 217416 610020 217468 610026
rect 217416 609962 217468 609968
rect 217428 573510 217456 609962
rect 217508 590708 217560 590714
rect 217508 590650 217560 590656
rect 217416 573504 217468 573510
rect 217416 573446 217468 573452
rect 217520 559706 217548 590650
rect 217876 559768 217928 559774
rect 217876 559710 217928 559716
rect 217508 559700 217560 559706
rect 217508 559642 217560 559648
rect 217324 555960 217376 555966
rect 217324 555902 217376 555908
rect 217888 552976 217916 559710
rect 218624 552976 218652 620978
rect 219256 585200 219308 585206
rect 219256 585142 219308 585148
rect 219268 552976 219296 585142
rect 220096 555762 220124 643486
rect 220176 643408 220228 643414
rect 220176 643350 220228 643356
rect 220188 555830 220216 643350
rect 222844 641912 222896 641918
rect 222844 641854 222896 641860
rect 220268 607232 220320 607238
rect 220268 607174 220320 607180
rect 220280 557054 220308 607174
rect 220728 577720 220780 577726
rect 220728 577662 220780 577668
rect 220268 557048 220320 557054
rect 220268 556990 220320 556996
rect 220176 555824 220228 555830
rect 220176 555766 220228 555772
rect 220084 555756 220136 555762
rect 220084 555698 220136 555704
rect 219992 555280 220044 555286
rect 219992 555222 220044 555228
rect 220004 552976 220032 555222
rect 220740 552976 220768 577662
rect 222200 577584 222252 577590
rect 222200 577526 222252 577532
rect 221464 555824 221516 555830
rect 221464 555766 221516 555772
rect 221476 552976 221504 555766
rect 222212 552976 222240 577526
rect 222856 552976 222884 641854
rect 222948 556986 222976 644710
rect 223580 642388 223632 642394
rect 223580 642330 223632 642336
rect 223488 582412 223540 582418
rect 223488 582354 223540 582360
rect 223500 577522 223528 582354
rect 223488 577516 223540 577522
rect 223488 577458 223540 577464
rect 222936 556980 222988 556986
rect 222936 556922 222988 556928
rect 223592 552976 223620 642330
rect 224316 625184 224368 625190
rect 224316 625126 224368 625132
rect 224328 552976 224356 625126
rect 225788 555892 225840 555898
rect 225788 555834 225840 555840
rect 225052 555688 225104 555694
rect 225052 555630 225104 555636
rect 225064 552976 225092 555630
rect 225800 552976 225828 555834
rect 226444 552976 226472 644982
rect 232504 644904 232556 644910
rect 232504 644846 232556 644852
rect 231124 644836 231176 644842
rect 231124 644778 231176 644784
rect 228364 643476 228416 643482
rect 228364 643418 228416 643424
rect 227168 587920 227220 587926
rect 227168 587862 227220 587868
rect 227180 552976 227208 587862
rect 227904 577856 227956 577862
rect 227904 577798 227956 577804
rect 227916 552976 227944 577798
rect 228376 555286 228404 643418
rect 229744 603152 229796 603158
rect 229744 603094 229796 603100
rect 228640 576360 228692 576366
rect 228640 576302 228692 576308
rect 228364 555280 228416 555286
rect 228364 555222 228416 555228
rect 228652 552976 228680 576302
rect 229284 569220 229336 569226
rect 229284 569162 229336 569168
rect 229296 552976 229324 569162
rect 229756 562494 229784 603094
rect 229744 562488 229796 562494
rect 229744 562430 229796 562436
rect 230756 555756 230808 555762
rect 230756 555698 230808 555704
rect 230020 555280 230072 555286
rect 230020 555222 230072 555228
rect 230032 552976 230060 555222
rect 230768 552976 230796 555698
rect 231136 555286 231164 644778
rect 231216 643340 231268 643346
rect 231216 643282 231268 643288
rect 231228 555626 231256 643282
rect 232228 577788 232280 577794
rect 232228 577730 232280 577736
rect 231308 577516 231360 577522
rect 231308 577458 231360 577464
rect 231320 555830 231348 577458
rect 231308 555824 231360 555830
rect 231308 555766 231360 555772
rect 231216 555620 231268 555626
rect 231216 555562 231268 555568
rect 231492 555620 231544 555626
rect 231492 555562 231544 555568
rect 231124 555280 231176 555286
rect 231124 555222 231176 555228
rect 231504 552976 231532 555562
rect 232240 552976 232268 577730
rect 232516 577658 232544 644846
rect 233608 633480 233660 633486
rect 233608 633422 233660 633428
rect 232596 630692 232648 630698
rect 232596 630634 232648 630640
rect 232504 577652 232556 577658
rect 232504 577594 232556 577600
rect 232608 568002 232636 630634
rect 232872 600364 232924 600370
rect 232872 600306 232924 600312
rect 232596 567996 232648 568002
rect 232596 567938 232648 567944
rect 232884 552976 232912 600306
rect 233620 552976 233648 633422
rect 233884 612808 233936 612814
rect 233884 612750 233936 612756
rect 233896 556850 233924 612750
rect 233884 556844 233936 556850
rect 233884 556786 233936 556792
rect 234356 552976 234384 646206
rect 235092 552976 235120 646478
rect 239404 646060 239456 646066
rect 239404 646002 239456 646008
rect 238024 645924 238076 645930
rect 238024 645866 238076 645872
rect 237472 644564 237524 644570
rect 237472 644506 237524 644512
rect 236644 643272 236696 643278
rect 236644 643214 236696 643220
rect 235264 640348 235316 640354
rect 235264 640290 235316 640296
rect 235276 563922 235304 640290
rect 235356 597576 235408 597582
rect 235356 597518 235408 597524
rect 235264 563916 235316 563922
rect 235264 563858 235316 563864
rect 235368 559638 235396 597518
rect 235448 577652 235500 577658
rect 235448 577594 235500 577600
rect 235356 559632 235408 559638
rect 235356 559574 235408 559580
rect 235460 555898 235488 577594
rect 235448 555892 235500 555898
rect 235448 555834 235500 555840
rect 236656 555490 236684 643214
rect 237378 640792 237434 640801
rect 237378 640727 237434 640736
rect 237392 640354 237420 640727
rect 237380 640348 237432 640354
rect 237380 640290 237432 640296
rect 237484 638246 237512 644506
rect 238036 641782 238064 645866
rect 238852 645176 238904 645182
rect 238852 645118 238904 645124
rect 238116 643612 238168 643618
rect 238116 643554 238168 643560
rect 238024 641776 238076 641782
rect 238024 641718 238076 641724
rect 237472 638240 237524 638246
rect 237472 638182 237524 638188
rect 237378 634400 237434 634409
rect 237378 634335 237434 634344
rect 237392 633486 237420 634335
rect 237380 633480 237432 633486
rect 237380 633422 237432 633428
rect 237378 631680 237434 631689
rect 237378 631615 237434 631624
rect 237392 630698 237420 631615
rect 237380 630692 237432 630698
rect 237380 630634 237432 630640
rect 237378 625560 237434 625569
rect 237378 625495 237434 625504
rect 237392 625190 237420 625495
rect 237380 625184 237432 625190
rect 237380 625126 237432 625132
rect 237378 622160 237434 622169
rect 237378 622095 237434 622104
rect 237392 621042 237420 622095
rect 237380 621036 237432 621042
rect 237380 620978 237432 620984
rect 238036 616185 238064 641718
rect 238022 616176 238078 616185
rect 238022 616111 238078 616120
rect 237378 613320 237434 613329
rect 237378 613255 237434 613264
rect 237392 612814 237420 613255
rect 237380 612808 237432 612814
rect 237380 612750 237432 612756
rect 237378 610056 237434 610065
rect 237378 609991 237380 610000
rect 237432 609991 237434 610000
rect 237380 609962 237432 609968
rect 237378 607336 237434 607345
rect 237378 607271 237434 607280
rect 237392 607238 237420 607271
rect 237380 607232 237432 607238
rect 237380 607174 237432 607180
rect 237378 603800 237434 603809
rect 237378 603735 237434 603744
rect 237392 603158 237420 603735
rect 237380 603152 237432 603158
rect 237380 603094 237432 603100
rect 237378 601080 237434 601089
rect 237378 601015 237434 601024
rect 237392 600370 237420 601015
rect 237380 600364 237432 600370
rect 237380 600306 237432 600312
rect 237378 597680 237434 597689
rect 237378 597615 237434 597624
rect 237392 597582 237420 597615
rect 237380 597576 237432 597582
rect 237380 597518 237432 597524
rect 237378 594960 237434 594969
rect 237378 594895 237434 594904
rect 237392 594862 237420 594895
rect 237380 594856 237432 594862
rect 237380 594798 237432 594804
rect 237378 591560 237434 591569
rect 237378 591495 237434 591504
rect 237392 590714 237420 591495
rect 237380 590708 237432 590714
rect 237380 590650 237432 590656
rect 237378 588840 237434 588849
rect 237378 588775 237434 588784
rect 237392 587926 237420 588775
rect 237380 587920 237432 587926
rect 237380 587862 237432 587868
rect 237378 585440 237434 585449
rect 237378 585375 237434 585384
rect 237392 585206 237420 585375
rect 237380 585200 237432 585206
rect 237380 585142 237432 585148
rect 237378 582720 237434 582729
rect 237378 582655 237434 582664
rect 237392 582418 237420 582655
rect 237380 582412 237432 582418
rect 237380 582354 237432 582360
rect 237932 557592 237984 557598
rect 237932 557534 237984 557540
rect 236644 555484 236696 555490
rect 236644 555426 236696 555432
rect 237196 555484 237248 555490
rect 237196 555426 237248 555432
rect 236460 554260 236512 554266
rect 236460 554202 236512 554208
rect 235816 554192 235868 554198
rect 235816 554134 235868 554140
rect 235828 552976 235856 554134
rect 236472 552976 236500 554202
rect 237208 552976 237236 555426
rect 237944 552976 237972 557534
rect 238128 555558 238156 643554
rect 238206 637800 238262 637809
rect 238206 637735 238262 637744
rect 238220 558414 238248 637735
rect 238298 628280 238354 628289
rect 238298 628215 238354 628224
rect 238208 558408 238260 558414
rect 238208 558350 238260 558356
rect 238312 558346 238340 628215
rect 238864 619585 238892 645118
rect 238944 638648 238996 638654
rect 238944 638590 238996 638596
rect 238850 619576 238906 619585
rect 238850 619511 238906 619520
rect 238956 570858 238984 638590
rect 238944 570852 238996 570858
rect 238944 570794 238996 570800
rect 238300 558340 238352 558346
rect 238300 558282 238352 558288
rect 238116 555552 238168 555558
rect 238116 555494 238168 555500
rect 238666 554976 238722 554985
rect 238666 554911 238722 554920
rect 238680 552976 238708 554911
rect 239416 552976 239444 646002
rect 245660 645108 245712 645114
rect 245660 645050 245712 645056
rect 239680 644700 239732 644706
rect 239680 644642 239732 644648
rect 239588 644632 239640 644638
rect 239588 644574 239640 644580
rect 239496 644496 239548 644502
rect 239496 644438 239548 644444
rect 239508 569362 239536 644438
rect 239600 572286 239628 644574
rect 239692 573578 239720 644642
rect 242900 644496 242952 644502
rect 242900 644438 242952 644444
rect 242912 643090 242940 644438
rect 245672 643090 245700 645050
rect 300308 645040 300360 645046
rect 300308 644982 300360 644988
rect 289268 644972 289320 644978
rect 289268 644914 289320 644920
rect 271972 644904 272024 644910
rect 271972 644846 272024 644852
rect 248788 644836 248840 644842
rect 248788 644778 248840 644784
rect 249156 644836 249208 644842
rect 249156 644778 249208 644784
rect 248800 643090 248828 644778
rect 242912 643062 243294 643090
rect 245672 643062 245870 643090
rect 248800 643062 249090 643090
rect 239784 642382 240074 642410
rect 249168 642394 249196 644778
rect 251364 644632 251416 644638
rect 251364 644574 251416 644580
rect 251376 643090 251404 644574
rect 254492 644564 254544 644570
rect 254492 644506 254544 644512
rect 254504 643090 254532 644506
rect 268660 643612 268712 643618
rect 268660 643554 268712 643560
rect 257068 643544 257120 643550
rect 257068 643486 257120 643492
rect 257080 643090 257108 643486
rect 266544 643476 266596 643482
rect 266544 643418 266596 643424
rect 260380 643408 260432 643414
rect 260380 643350 260432 643356
rect 260392 643090 260420 643350
rect 251376 643062 251666 643090
rect 254504 643062 254886 643090
rect 257080 643062 257462 643090
rect 260392 643062 260682 643090
rect 266556 642954 266584 643418
rect 268672 643090 268700 643554
rect 271984 643090 272012 644846
rect 277676 644768 277728 644774
rect 277676 644710 277728 644716
rect 274640 643204 274692 643210
rect 274640 643146 274692 643152
rect 274652 643090 274680 643146
rect 277688 643090 277716 644710
rect 280252 643340 280304 643346
rect 280252 643282 280304 643288
rect 280264 643090 280292 643282
rect 286140 643136 286192 643142
rect 268672 643062 269054 643090
rect 271984 643062 272274 643090
rect 274652 643062 274850 643090
rect 277688 643062 278070 643090
rect 280264 643062 280646 643090
rect 289280 643090 289308 644914
rect 295524 644836 295576 644842
rect 295524 644778 295576 644784
rect 291844 643272 291896 643278
rect 291844 643214 291896 643220
rect 291856 643090 291884 643214
rect 295536 643090 295564 644778
rect 297732 644700 297784 644706
rect 297732 644642 297784 644648
rect 286192 643084 286442 643090
rect 286140 643078 286442 643084
rect 286152 643062 286442 643078
rect 289280 643062 289662 643090
rect 291856 643062 292238 643090
rect 295458 643062 295564 643090
rect 297744 643090 297772 644642
rect 300320 643090 300348 644982
rect 304264 644904 304316 644910
rect 304264 644846 304316 644852
rect 297744 643062 298034 643090
rect 300320 643062 300610 643090
rect 266478 642926 266584 642954
rect 262968 642394 263258 642410
rect 283576 642394 283866 642410
rect 249156 642388 249208 642394
rect 239784 638654 239812 642382
rect 249156 642330 249208 642336
rect 262956 642388 263258 642394
rect 263008 642382 263258 642388
rect 283564 642388 283866 642394
rect 262956 642330 263008 642336
rect 283616 642382 283866 642388
rect 283564 642330 283616 642336
rect 300858 639432 300914 639441
rect 300858 639367 300914 639376
rect 239772 638648 239824 638654
rect 239772 638590 239824 638596
rect 300674 581632 300730 581641
rect 300674 581567 300730 581576
rect 239784 580094 240074 580122
rect 242360 580094 242650 580122
rect 244292 580094 245226 580122
rect 248446 580094 248552 580122
rect 239784 577522 239812 580094
rect 242360 577658 242388 580094
rect 242348 577652 242400 577658
rect 242348 577594 242400 577600
rect 239772 577516 239824 577522
rect 239772 577458 239824 577464
rect 242164 576972 242216 576978
rect 242164 576914 242216 576920
rect 239680 573572 239732 573578
rect 239680 573514 239732 573520
rect 240784 573504 240836 573510
rect 240784 573446 240836 573452
rect 239588 572280 239640 572286
rect 239588 572222 239640 572228
rect 239496 569356 239548 569362
rect 239496 569298 239548 569304
rect 240048 554328 240100 554334
rect 240048 554270 240100 554276
rect 240060 552976 240088 554270
rect 240796 552976 240824 573446
rect 242176 555694 242204 576914
rect 244292 566710 244320 580094
rect 245844 579216 245896 579222
rect 245844 579158 245896 579164
rect 244924 576904 244976 576910
rect 244924 576846 244976 576852
rect 244280 566704 244332 566710
rect 244280 566646 244332 566652
rect 242900 563848 242952 563854
rect 242900 563790 242952 563796
rect 242164 555688 242216 555694
rect 242164 555630 242216 555636
rect 242256 555416 242308 555422
rect 242256 555358 242308 555364
rect 241518 555112 241574 555121
rect 241518 555047 241574 555056
rect 241532 552976 241560 555047
rect 242268 552976 242296 555358
rect 242912 552976 242940 563790
rect 244936 555762 244964 576846
rect 245108 563916 245160 563922
rect 245108 563858 245160 563864
rect 244924 555756 244976 555762
rect 244924 555698 244976 555704
rect 243636 553784 243688 553790
rect 243636 553726 243688 553732
rect 243648 552976 243676 553726
rect 244372 553580 244424 553586
rect 244372 553522 244424 553528
rect 244384 552976 244412 553522
rect 245120 552976 245148 563858
rect 245856 552976 245884 579158
rect 248524 576978 248552 580094
rect 250640 580094 251022 580122
rect 253952 580094 254242 580122
rect 256818 580094 256924 580122
rect 249064 577652 249116 577658
rect 249064 577594 249116 577600
rect 248512 576972 248564 576978
rect 248512 576914 248564 576920
rect 247960 567928 248012 567934
rect 247960 567870 248012 567876
rect 246488 565208 246540 565214
rect 246488 565150 246540 565156
rect 246500 552976 246528 565150
rect 247224 553852 247276 553858
rect 247224 553794 247276 553800
rect 247236 552976 247264 553794
rect 247972 552976 248000 567870
rect 248696 557660 248748 557666
rect 248696 557602 248748 557608
rect 248708 552976 248736 557602
rect 249076 555626 249104 577594
rect 250640 576910 250668 580094
rect 250628 576904 250680 576910
rect 250628 576846 250680 576852
rect 253664 570784 253716 570790
rect 253664 570726 253716 570732
rect 250812 569288 250864 569294
rect 250812 569230 250864 569236
rect 250076 566636 250128 566642
rect 250076 566578 250128 566584
rect 249064 555620 249116 555626
rect 249064 555562 249116 555568
rect 249430 553888 249486 553897
rect 249430 553823 249486 553832
rect 249444 552976 249472 553823
rect 250088 552976 250116 566578
rect 250824 552976 250852 569230
rect 251548 561060 251600 561066
rect 251548 561002 251600 561008
rect 251560 552976 251588 561002
rect 252284 557728 252336 557734
rect 252284 557670 252336 557676
rect 252296 552976 252324 557670
rect 252928 555620 252980 555626
rect 252928 555562 252980 555568
rect 252940 552976 252968 555562
rect 253676 552976 253704 570726
rect 253952 556918 253980 580094
rect 256896 567194 256924 580094
rect 259656 580094 260038 580122
rect 262232 580094 262614 580122
rect 265544 580094 265834 580122
rect 268120 580094 268410 580122
rect 271248 580094 271630 580122
rect 273824 580094 274206 580122
rect 277426 580094 277532 580122
rect 258724 579284 258776 579290
rect 258724 579226 258776 579232
rect 257988 577516 258040 577522
rect 257988 577458 258040 577464
rect 256712 567166 256924 567194
rect 256712 565350 256740 567166
rect 256700 565344 256752 565350
rect 256700 565286 256752 565292
rect 256516 559700 256568 559706
rect 256516 559642 256568 559648
rect 253940 556912 253992 556918
rect 253940 556854 253992 556860
rect 255872 556572 255924 556578
rect 255872 556514 255924 556520
rect 254400 556232 254452 556238
rect 254400 556174 254452 556180
rect 254412 552976 254440 556174
rect 255134 555520 255190 555529
rect 255134 555455 255190 555464
rect 255148 552976 255176 555455
rect 255884 552976 255912 556514
rect 256528 552976 256556 559642
rect 257252 555008 257304 555014
rect 257252 554950 257304 554956
rect 257264 552976 257292 554950
rect 258000 552976 258028 577458
rect 258736 552976 258764 579226
rect 259656 577658 259684 580094
rect 259644 577652 259696 577658
rect 259644 577594 259696 577600
rect 259460 566704 259512 566710
rect 259460 566646 259512 566652
rect 259472 552976 259500 566646
rect 262232 561134 262260 580094
rect 265544 577862 265572 580094
rect 265532 577856 265584 577862
rect 265532 577798 265584 577804
rect 268120 577726 268148 580094
rect 268108 577720 268160 577726
rect 268108 577662 268160 577668
rect 271248 577250 271276 580094
rect 273824 577590 273852 580094
rect 273904 577720 273956 577726
rect 273904 577662 273956 577668
rect 273812 577584 273864 577590
rect 273812 577526 273864 577532
rect 269764 577244 269816 577250
rect 269764 577186 269816 577192
rect 271236 577244 271288 577250
rect 271236 577186 271288 577192
rect 266544 575000 266596 575006
rect 266544 574942 266596 574948
rect 263692 567996 263744 568002
rect 263692 567938 263744 567944
rect 262220 561128 262272 561134
rect 262220 561070 262272 561076
rect 260104 559632 260156 559638
rect 260104 559574 260156 559580
rect 260116 552976 260144 559574
rect 263048 556300 263100 556306
rect 263048 556242 263100 556248
rect 261576 555552 261628 555558
rect 261576 555494 261628 555500
rect 260840 553988 260892 553994
rect 260840 553930 260892 553936
rect 260852 552976 260880 553930
rect 261588 552976 261616 555494
rect 262312 553716 262364 553722
rect 262312 553658 262364 553664
rect 262324 552976 262352 553658
rect 263060 552976 263088 556242
rect 263704 552976 263732 567938
rect 264428 556436 264480 556442
rect 264428 556378 264480 556384
rect 264440 552976 264468 556378
rect 265900 556368 265952 556374
rect 265900 556310 265952 556316
rect 265164 554940 265216 554946
rect 265164 554882 265216 554888
rect 265176 552976 265204 554882
rect 265912 552976 265940 556310
rect 266556 552976 266584 574942
rect 267280 572144 267332 572150
rect 267280 572086 267332 572092
rect 267292 552976 267320 572086
rect 268016 571396 268068 571402
rect 268016 571338 268068 571344
rect 268028 552976 268056 571338
rect 269488 570852 269540 570858
rect 269488 570794 269540 570800
rect 268752 554124 268804 554130
rect 268752 554066 268804 554072
rect 268764 552976 268792 554066
rect 269500 552976 269528 570794
rect 269776 558278 269804 577186
rect 273916 559774 273944 577662
rect 274456 569356 274508 569362
rect 274456 569298 274508 569304
rect 273904 559768 273956 559774
rect 273904 559710 273956 559716
rect 269764 558272 269816 558278
rect 269764 558214 269816 558220
rect 271604 558272 271656 558278
rect 271604 558214 271656 558220
rect 270132 556844 270184 556850
rect 270132 556786 270184 556792
rect 270144 552976 270172 556786
rect 270868 555688 270920 555694
rect 270868 555630 270920 555636
rect 270880 552976 270908 555630
rect 271616 552976 271644 558214
rect 273720 556504 273772 556510
rect 273720 556446 273772 556452
rect 272340 553920 272392 553926
rect 272340 553862 272392 553868
rect 272352 552976 272380 553862
rect 273076 553444 273128 553450
rect 273076 553386 273128 553392
rect 273088 552976 273116 553386
rect 273732 552976 273760 556446
rect 274468 552976 274496 569298
rect 277504 567194 277532 580094
rect 279712 580094 280002 580122
rect 282932 580094 283222 580122
rect 285798 580094 285904 580122
rect 279712 577794 279740 580094
rect 279700 577788 279752 577794
rect 279700 577730 279752 577736
rect 282932 577726 282960 580094
rect 282920 577720 282972 577726
rect 282920 577662 282972 577668
rect 280804 577652 280856 577658
rect 280804 577594 280856 577600
rect 277412 567166 277532 567194
rect 277412 566574 277440 567166
rect 277400 566568 277452 566574
rect 277400 566510 277452 566516
rect 279516 566568 279568 566574
rect 279516 566510 279568 566516
rect 275192 565276 275244 565282
rect 275192 565218 275244 565224
rect 274640 554940 274692 554946
rect 274640 554882 274692 554888
rect 274652 554062 274680 554882
rect 274640 554056 274692 554062
rect 274640 553998 274692 554004
rect 275204 552976 275232 565218
rect 278044 555756 278096 555762
rect 278044 555698 278096 555704
rect 276572 555348 276624 555354
rect 276572 555290 276624 555296
rect 275928 555212 275980 555218
rect 275928 555154 275980 555160
rect 275940 552976 275968 555154
rect 276584 552976 276612 555290
rect 277308 555280 277360 555286
rect 277308 555222 277360 555228
rect 277320 552976 277348 555222
rect 278056 552976 278084 555698
rect 278780 553512 278832 553518
rect 278780 553454 278832 553460
rect 278792 552976 278820 553454
rect 279528 552976 279556 566510
rect 280816 563786 280844 577594
rect 280896 577584 280948 577590
rect 280896 577526 280948 577532
rect 280804 563780 280856 563786
rect 280804 563722 280856 563728
rect 280160 555076 280212 555082
rect 280160 555018 280212 555024
rect 280172 552976 280200 555018
rect 280908 552976 280936 577526
rect 282184 576904 282236 576910
rect 282184 576846 282236 576852
rect 282196 562358 282224 576846
rect 285876 567866 285904 580094
rect 288728 580094 289018 580122
rect 291212 580094 291594 580122
rect 293972 580094 294814 580122
rect 297008 580094 297390 580122
rect 300320 580094 300610 580122
rect 288072 579420 288124 579426
rect 288072 579362 288124 579368
rect 286324 579352 286376 579358
rect 286324 579294 286376 579300
rect 285864 567860 285916 567866
rect 285864 567802 285916 567808
rect 282184 562352 282236 562358
rect 282184 562294 282236 562300
rect 283748 558340 283800 558346
rect 283748 558282 283800 558288
rect 283104 557864 283156 557870
rect 283104 557806 283156 557812
rect 282368 556912 282420 556918
rect 282368 556854 282420 556860
rect 281632 554872 281684 554878
rect 281632 554814 281684 554820
rect 281644 552976 281672 554814
rect 282380 552976 282408 556854
rect 283116 552976 283144 557806
rect 283760 552976 283788 558282
rect 284944 557796 284996 557802
rect 284944 557738 284996 557744
rect 284956 555490 284984 557738
rect 285220 556640 285272 556646
rect 285220 556582 285272 556588
rect 284944 555484 284996 555490
rect 284944 555426 284996 555432
rect 284484 553648 284536 553654
rect 284484 553590 284536 553596
rect 284496 552976 284524 553590
rect 285232 552976 285260 556582
rect 286336 555558 286364 579294
rect 287336 557932 287388 557938
rect 287336 557874 287388 557880
rect 286324 555552 286376 555558
rect 286324 555494 286376 555500
rect 286690 555248 286746 555257
rect 286690 555183 286746 555192
rect 285954 554840 286010 554849
rect 285954 554775 286010 554784
rect 285968 552976 285996 554775
rect 286704 552976 286732 555183
rect 287348 552976 287376 557874
rect 288084 552976 288112 579362
rect 288728 576910 288756 580094
rect 289544 579556 289596 579562
rect 289544 579498 289596 579504
rect 288808 579488 288860 579494
rect 288808 579430 288860 579436
rect 288716 576904 288768 576910
rect 288716 576846 288768 576852
rect 288820 552976 288848 579430
rect 289084 577720 289136 577726
rect 289084 577662 289136 577668
rect 289096 566506 289124 577662
rect 289084 566500 289136 566506
rect 289084 566442 289136 566448
rect 289556 552976 289584 579498
rect 290188 578876 290240 578882
rect 290188 578818 290240 578824
rect 290200 552976 290228 578818
rect 291212 565146 291240 580094
rect 292396 578740 292448 578746
rect 292396 578682 292448 578688
rect 291200 565140 291252 565146
rect 291200 565082 291252 565088
rect 291660 556708 291712 556714
rect 291660 556650 291712 556656
rect 290924 555144 290976 555150
rect 290924 555086 290976 555092
rect 290936 552976 290964 555086
rect 291672 552976 291700 556650
rect 292408 552976 292436 578682
rect 293972 570654 294000 580094
rect 295248 579624 295300 579630
rect 295248 579566 295300 579572
rect 293960 570648 294012 570654
rect 293960 570590 294012 570596
rect 293130 553752 293186 553761
rect 293130 553687 293186 553696
rect 293144 552976 293172 553687
rect 293774 553616 293830 553625
rect 293774 553551 293830 553560
rect 293788 552976 293816 553551
rect 294510 553480 294566 553489
rect 294510 553415 294566 553424
rect 294524 552976 294552 553415
rect 295260 552976 295288 579566
rect 297008 577658 297036 580094
rect 297364 578808 297416 578814
rect 297364 578750 297416 578756
rect 296996 577652 297048 577658
rect 296996 577594 297048 577600
rect 295984 554804 296036 554810
rect 295984 554746 296036 554752
rect 296812 554804 296864 554810
rect 296812 554746 296864 554752
rect 295996 552976 296024 554746
rect 296824 553058 296852 554746
rect 296748 553030 296852 553058
rect 296748 552976 296776 553030
rect 297376 552976 297404 578750
rect 300320 577726 300348 580094
rect 300308 577720 300360 577726
rect 300308 577662 300360 577668
rect 300688 560998 300716 581567
rect 300872 576230 300900 639367
rect 300950 636712 301006 636721
rect 300950 636647 301006 636656
rect 300964 576366 300992 636647
rect 302238 633448 302294 633457
rect 302238 633383 302294 633392
rect 301042 630728 301098 630737
rect 301042 630663 301098 630672
rect 301056 579018 301084 630663
rect 301134 624472 301190 624481
rect 301134 624407 301190 624416
rect 301044 579012 301096 579018
rect 301044 578954 301096 578960
rect 300952 576360 301004 576366
rect 300952 576302 301004 576308
rect 300860 576224 300912 576230
rect 300860 576166 300912 576172
rect 301148 573374 301176 624407
rect 301226 612912 301282 612921
rect 301226 612847 301282 612856
rect 301136 573368 301188 573374
rect 301136 573310 301188 573316
rect 301240 572082 301268 612847
rect 301318 606248 301374 606257
rect 301318 606183 301374 606192
rect 301332 574870 301360 606183
rect 301410 600672 301466 600681
rect 301410 600607 301466 600616
rect 301424 579154 301452 600607
rect 301502 593872 301558 593881
rect 301502 593807 301558 593816
rect 301412 579148 301464 579154
rect 301412 579090 301464 579096
rect 301320 574864 301372 574870
rect 301320 574806 301372 574812
rect 301516 573442 301544 593807
rect 301594 588024 301650 588033
rect 301594 587959 301650 587968
rect 301608 578950 301636 587959
rect 301596 578944 301648 578950
rect 301596 578886 301648 578892
rect 301504 573436 301556 573442
rect 301504 573378 301556 573384
rect 301228 572076 301280 572082
rect 301228 572018 301280 572024
rect 300676 560992 300728 560998
rect 300676 560934 300728 560940
rect 302252 559570 302280 633383
rect 302330 627192 302386 627201
rect 302330 627127 302386 627136
rect 302344 574938 302372 627127
rect 302422 621072 302478 621081
rect 302422 621007 302478 621016
rect 302332 574932 302384 574938
rect 302332 574874 302384 574880
rect 302436 563718 302464 621007
rect 302606 618352 302662 618361
rect 302606 618287 302662 618296
rect 302514 614952 302570 614961
rect 302514 614887 302570 614896
rect 302424 563712 302476 563718
rect 302424 563654 302476 563660
rect 302240 559564 302292 559570
rect 302240 559506 302292 559512
rect 302528 558210 302556 614887
rect 302620 579086 302648 618287
rect 303158 609512 303214 609521
rect 303158 609447 303214 609456
rect 303172 609278 303200 609447
rect 302792 609272 302844 609278
rect 302792 609214 302844 609220
rect 303160 609272 303212 609278
rect 303160 609214 303212 609220
rect 302698 603392 302754 603401
rect 302698 603327 302754 603336
rect 302608 579080 302660 579086
rect 302608 579022 302660 579028
rect 302712 570722 302740 603327
rect 302804 580922 302832 609214
rect 302974 596728 303030 596737
rect 302974 596663 303030 596672
rect 302882 590744 302938 590753
rect 302882 590679 302938 590688
rect 302792 580916 302844 580922
rect 302792 580858 302844 580864
rect 302700 570716 302752 570722
rect 302700 570658 302752 570664
rect 302516 558204 302568 558210
rect 302516 558146 302568 558152
rect 300308 555756 300360 555762
rect 300308 555698 300360 555704
rect 298652 555552 298704 555558
rect 298652 555494 298704 555500
rect 298098 555384 298154 555393
rect 298098 555319 298154 555328
rect 298112 552976 298140 555319
rect 298664 555218 298692 555494
rect 299572 555484 299624 555490
rect 299572 555426 299624 555432
rect 298836 555280 298888 555286
rect 298836 555222 298888 555228
rect 298652 555212 298704 555218
rect 298652 555154 298704 555160
rect 298848 552976 298876 555222
rect 299388 553512 299440 553518
rect 299388 553454 299440 553460
rect 299400 553382 299428 553454
rect 299388 553376 299440 553382
rect 299388 553318 299440 553324
rect 299584 552976 299612 555426
rect 300214 554976 300270 554985
rect 300214 554911 300270 554920
rect 300124 554804 300176 554810
rect 300124 554746 300176 554752
rect 300136 531078 300164 554746
rect 300228 534070 300256 554911
rect 300216 534064 300268 534070
rect 300216 534006 300268 534012
rect 300320 534002 300348 555698
rect 302056 555552 302108 555558
rect 302056 555494 302108 555500
rect 300400 555348 300452 555354
rect 300400 555290 300452 555296
rect 300308 533996 300360 534002
rect 300308 533938 300360 533944
rect 300412 532778 300440 555290
rect 301872 555212 301924 555218
rect 301872 555154 301924 555160
rect 300582 555112 300638 555121
rect 300582 555047 300638 555056
rect 300492 555008 300544 555014
rect 300492 554950 300544 554956
rect 300504 533934 300532 554950
rect 300596 534585 300624 555047
rect 301504 554940 301556 554946
rect 301504 554882 301556 554888
rect 300676 553784 300728 553790
rect 300676 553726 300728 553732
rect 300688 543726 300716 553726
rect 300676 543720 300728 543726
rect 300676 543662 300728 543668
rect 300582 534576 300638 534585
rect 300582 534511 300638 534520
rect 300492 533928 300544 533934
rect 300492 533870 300544 533876
rect 300400 532772 300452 532778
rect 300400 532714 300452 532720
rect 300124 531072 300176 531078
rect 300124 531014 300176 531020
rect 301516 530806 301544 554882
rect 301596 554872 301648 554878
rect 301596 554814 301648 554820
rect 301608 530942 301636 554814
rect 301780 553852 301832 553858
rect 301780 553794 301832 553800
rect 301688 553444 301740 553450
rect 301688 553386 301740 553392
rect 301700 532302 301728 553386
rect 301688 532296 301740 532302
rect 301688 532238 301740 532244
rect 301792 532166 301820 553794
rect 301884 533866 301912 555154
rect 301962 553888 302018 553897
rect 301962 553823 302018 553832
rect 301872 533860 301924 533866
rect 301872 533802 301924 533808
rect 301976 532681 302004 553823
rect 302068 532914 302096 555494
rect 302238 545456 302294 545465
rect 302238 545391 302294 545400
rect 302252 545154 302280 545391
rect 302240 545148 302292 545154
rect 302240 545090 302292 545096
rect 302056 532908 302108 532914
rect 302056 532850 302108 532856
rect 301962 532672 302018 532681
rect 301962 532607 302018 532616
rect 301780 532160 301832 532166
rect 301780 532102 301832 532108
rect 301596 530936 301648 530942
rect 301596 530878 301648 530884
rect 301504 530800 301556 530806
rect 301504 530742 301556 530748
rect 302422 530496 302478 530505
rect 302422 530431 302478 530440
rect 302436 529990 302464 530431
rect 302424 529984 302476 529990
rect 302424 529926 302476 529932
rect 57702 523016 57758 523025
rect 57702 522951 57758 522960
rect 57886 523016 57942 523025
rect 57886 522951 57942 522960
rect 57716 521762 57744 522951
rect 53748 521756 53800 521762
rect 53748 521698 53800 521704
rect 57704 521756 57756 521762
rect 57704 521698 57756 521704
rect 49424 492176 49476 492182
rect 49424 492118 49476 492124
rect 49056 490680 49108 490686
rect 49056 490622 49108 490628
rect 41052 490612 41104 490618
rect 41052 490554 41104 490560
rect 40960 482452 41012 482458
rect 40960 482394 41012 482400
rect 40868 467492 40920 467498
rect 40868 467434 40920 467440
rect 40880 378078 40908 467434
rect 40868 378072 40920 378078
rect 40868 378014 40920 378020
rect 18604 358760 18656 358766
rect 18604 358702 18656 358708
rect 40972 268258 41000 482394
rect 41064 271658 41092 490554
rect 47952 488504 48004 488510
rect 47952 488446 48004 488452
rect 46388 488300 46440 488306
rect 46388 488242 46440 488248
rect 46296 488164 46348 488170
rect 46296 488106 46348 488112
rect 44088 485648 44140 485654
rect 41326 485616 41382 485625
rect 44088 485590 44140 485596
rect 41326 485551 41382 485560
rect 41144 467424 41196 467430
rect 41144 467366 41196 467372
rect 41052 271652 41104 271658
rect 41052 271594 41104 271600
rect 40960 268252 41012 268258
rect 40960 268194 41012 268200
rect 41156 166326 41184 467366
rect 41236 467356 41288 467362
rect 41236 467298 41288 467304
rect 41144 166320 41196 166326
rect 41144 166262 41196 166268
rect 41248 56574 41276 467298
rect 41340 70378 41368 485551
rect 43994 485072 44050 485081
rect 43994 485007 44050 485016
rect 43628 482724 43680 482730
rect 43628 482666 43680 482672
rect 43260 482316 43312 482322
rect 43260 482258 43312 482264
rect 42616 471300 42668 471306
rect 42616 471242 42668 471248
rect 42524 467560 42576 467566
rect 42524 467502 42576 467508
rect 42536 377058 42564 467502
rect 42524 377052 42576 377058
rect 42524 376994 42576 377000
rect 42628 273630 42656 471242
rect 42708 467288 42760 467294
rect 42708 467230 42760 467236
rect 42616 273624 42668 273630
rect 42616 273566 42668 273572
rect 42720 166394 42748 467230
rect 43272 391950 43300 482258
rect 43352 474700 43404 474706
rect 43352 474642 43404 474648
rect 43260 391944 43312 391950
rect 43260 391886 43312 391892
rect 43364 273562 43392 474642
rect 43536 474292 43588 474298
rect 43536 474234 43588 474240
rect 43444 473952 43496 473958
rect 43444 473894 43496 473900
rect 43352 273556 43404 273562
rect 43352 273498 43404 273504
rect 43456 271726 43484 473894
rect 43444 271720 43496 271726
rect 43444 271662 43496 271668
rect 43548 268326 43576 474234
rect 43640 268870 43668 482666
rect 43812 482656 43864 482662
rect 43812 482598 43864 482604
rect 43720 482520 43772 482526
rect 43720 482462 43772 482468
rect 43628 268864 43680 268870
rect 43628 268806 43680 268812
rect 43732 268530 43760 482462
rect 43720 268524 43772 268530
rect 43720 268466 43772 268472
rect 43824 268394 43852 482598
rect 43904 482588 43956 482594
rect 43904 482530 43956 482536
rect 43916 268462 43944 482530
rect 44008 268666 44036 485007
rect 44100 268938 44128 485590
rect 44640 485240 44692 485246
rect 44640 485182 44692 485188
rect 44652 379166 44680 485182
rect 44824 485172 44876 485178
rect 44824 485114 44876 485120
rect 44732 471164 44784 471170
rect 44732 471106 44784 471112
rect 44640 379160 44692 379166
rect 44640 379102 44692 379108
rect 44744 378214 44772 471106
rect 44836 379098 44864 485114
rect 46204 485104 46256 485110
rect 46204 485046 46256 485052
rect 45192 474428 45244 474434
rect 45192 474370 45244 474376
rect 45100 474360 45152 474366
rect 45100 474302 45152 474308
rect 45008 474224 45060 474230
rect 45008 474166 45060 474172
rect 44916 467152 44968 467158
rect 44916 467094 44968 467100
rect 44824 379092 44876 379098
rect 44824 379034 44876 379040
rect 44732 378208 44784 378214
rect 44732 378150 44784 378156
rect 44928 270502 44956 467094
rect 45020 273426 45048 474166
rect 45008 273420 45060 273426
rect 45008 273362 45060 273368
rect 45112 273358 45140 474302
rect 45204 273494 45232 474370
rect 45376 474156 45428 474162
rect 45376 474098 45428 474104
rect 45284 474088 45336 474094
rect 45284 474030 45336 474036
rect 45296 273698 45324 474030
rect 45284 273692 45336 273698
rect 45284 273634 45336 273640
rect 45192 273488 45244 273494
rect 45192 273430 45244 273436
rect 45100 273352 45152 273358
rect 45100 273294 45152 273300
rect 45388 271862 45416 474098
rect 46112 468376 46164 468382
rect 46112 468318 46164 468324
rect 46020 464296 46072 464302
rect 46020 464238 46072 464244
rect 46032 418130 46060 464238
rect 46020 418124 46072 418130
rect 46020 418066 46072 418072
rect 45468 388476 45520 388482
rect 45468 388418 45520 388424
rect 45480 281518 45508 388418
rect 46124 379409 46152 468318
rect 46110 379400 46166 379409
rect 46110 379335 46166 379344
rect 45468 281512 45520 281518
rect 45468 281454 45520 281460
rect 45376 271856 45428 271862
rect 45376 271798 45428 271804
rect 46124 271454 46152 379335
rect 46216 379030 46244 485046
rect 46204 379024 46256 379030
rect 46204 378966 46256 378972
rect 46308 300830 46336 488106
rect 46296 300824 46348 300830
rect 46296 300766 46348 300772
rect 46400 272134 46428 488242
rect 46662 488064 46718 488073
rect 46662 487999 46718 488008
rect 46848 488028 46900 488034
rect 46478 487928 46534 487937
rect 46478 487863 46534 487872
rect 46492 272950 46520 487863
rect 46570 485208 46626 485217
rect 46570 485143 46626 485152
rect 46480 272944 46532 272950
rect 46480 272886 46532 272892
rect 46388 272128 46440 272134
rect 46388 272070 46440 272076
rect 46112 271448 46164 271454
rect 46112 271390 46164 271396
rect 44916 270496 44968 270502
rect 44916 270438 44968 270444
rect 44088 268932 44140 268938
rect 44088 268874 44140 268880
rect 43996 268660 44048 268666
rect 43996 268602 44048 268608
rect 43904 268456 43956 268462
rect 43904 268398 43956 268404
rect 43812 268388 43864 268394
rect 43812 268330 43864 268336
rect 43536 268320 43588 268326
rect 43536 268262 43588 268268
rect 46400 267734 46428 272070
rect 46584 268598 46612 485143
rect 46676 271590 46704 487999
rect 46848 487970 46900 487976
rect 46756 485036 46808 485042
rect 46756 484978 46808 484984
rect 46664 271584 46716 271590
rect 46664 271526 46716 271532
rect 46664 271448 46716 271454
rect 46664 271390 46716 271396
rect 46676 271046 46704 271390
rect 46664 271040 46716 271046
rect 46664 270982 46716 270988
rect 46572 268592 46624 268598
rect 46572 268534 46624 268540
rect 46400 267706 46520 267734
rect 42708 166388 42760 166394
rect 42708 166330 42760 166336
rect 46492 145382 46520 267706
rect 46676 146266 46704 270982
rect 46768 268734 46796 484978
rect 46860 269006 46888 487970
rect 47768 485444 47820 485450
rect 47768 485386 47820 485392
rect 47676 471096 47728 471102
rect 47676 471038 47728 471044
rect 47584 464364 47636 464370
rect 47584 464306 47636 464312
rect 47596 418062 47624 464306
rect 47584 418056 47636 418062
rect 47584 417998 47636 418004
rect 47492 414044 47544 414050
rect 47492 413986 47544 413992
rect 47400 412684 47452 412690
rect 47400 412626 47452 412632
rect 47412 380866 47440 412626
rect 47400 380860 47452 380866
rect 47400 380802 47452 380808
rect 47504 380798 47532 413986
rect 47584 411324 47636 411330
rect 47584 411266 47636 411272
rect 47492 380792 47544 380798
rect 47492 380734 47544 380740
rect 47490 379128 47546 379137
rect 47490 379063 47546 379072
rect 47504 271833 47532 379063
rect 47596 376990 47624 411266
rect 47688 379273 47716 471038
rect 47780 389162 47808 485386
rect 47860 485376 47912 485382
rect 47860 485318 47912 485324
rect 47768 389156 47820 389162
rect 47768 389098 47820 389104
rect 47674 379264 47730 379273
rect 47674 379199 47730 379208
rect 47584 376984 47636 376990
rect 47584 376926 47636 376932
rect 47490 271824 47546 271833
rect 47490 271759 47546 271768
rect 47688 271726 47716 379199
rect 47872 378622 47900 485318
rect 47860 378616 47912 378622
rect 47860 378558 47912 378564
rect 47768 378208 47820 378214
rect 47768 378150 47820 378156
rect 47780 287054 47808 378150
rect 47780 287026 47900 287054
rect 47676 271720 47728 271726
rect 47872 271697 47900 287026
rect 47964 272542 47992 488446
rect 48044 488368 48096 488374
rect 48044 488310 48096 488316
rect 47952 272536 48004 272542
rect 47952 272478 48004 272484
rect 48056 272406 48084 488310
rect 48964 488096 49016 488102
rect 48964 488038 49016 488044
rect 48872 487824 48924 487830
rect 48872 487766 48924 487772
rect 48134 485344 48190 485353
rect 48134 485279 48190 485288
rect 48044 272400 48096 272406
rect 48044 272342 48096 272348
rect 47952 271720 48004 271726
rect 47676 271662 47728 271668
rect 47858 271688 47914 271697
rect 47952 271662 48004 271668
rect 47858 271623 47914 271632
rect 46848 269000 46900 269006
rect 46848 268942 46900 268948
rect 46756 268728 46808 268734
rect 46756 268670 46808 268676
rect 47584 268524 47636 268530
rect 47584 268466 47636 268472
rect 47596 164218 47624 268466
rect 47768 268456 47820 268462
rect 47768 268398 47820 268404
rect 47676 268388 47728 268394
rect 47676 268330 47728 268336
rect 47584 164212 47636 164218
rect 47584 164154 47636 164160
rect 47688 148306 47716 268330
rect 47780 148850 47808 268398
rect 47768 148844 47820 148850
rect 47768 148786 47820 148792
rect 47872 148714 47900 271623
rect 47964 270978 47992 271662
rect 47952 270972 48004 270978
rect 47952 270914 48004 270920
rect 47964 148782 47992 270914
rect 47952 148776 48004 148782
rect 47952 148718 48004 148724
rect 47860 148708 47912 148714
rect 47860 148650 47912 148656
rect 47676 148300 47728 148306
rect 47676 148242 47728 148248
rect 46664 146260 46716 146266
rect 46664 146202 46716 146208
rect 48056 145450 48084 272342
rect 48148 269074 48176 485279
rect 48228 484968 48280 484974
rect 48228 484910 48280 484916
rect 48136 269068 48188 269074
rect 48136 269010 48188 269016
rect 48240 268802 48268 484910
rect 48780 482384 48832 482390
rect 48780 482326 48832 482332
rect 48792 380322 48820 482326
rect 48780 380316 48832 380322
rect 48780 380258 48832 380264
rect 48884 380186 48912 487766
rect 48872 380180 48924 380186
rect 48872 380122 48924 380128
rect 48976 272338 49004 488038
rect 49068 272746 49096 490622
rect 49146 488200 49202 488209
rect 49146 488135 49202 488144
rect 49056 272740 49108 272746
rect 49056 272682 49108 272688
rect 48964 272332 49016 272338
rect 48964 272274 49016 272280
rect 49054 271824 49110 271833
rect 49054 271759 49110 271768
rect 49068 271289 49096 271759
rect 49054 271280 49110 271289
rect 49054 271215 49110 271224
rect 48228 268796 48280 268802
rect 48228 268738 48280 268744
rect 48136 268660 48188 268666
rect 48136 268602 48188 268608
rect 48044 145444 48096 145450
rect 48044 145386 48096 145392
rect 46480 145376 46532 145382
rect 46480 145318 46532 145324
rect 48148 144702 48176 268602
rect 48228 268592 48280 268598
rect 48228 268534 48280 268540
rect 48136 144696 48188 144702
rect 48136 144638 48188 144644
rect 48240 144634 48268 268534
rect 49068 148646 49096 271215
rect 49160 250510 49188 488135
rect 49332 471776 49384 471782
rect 49332 471718 49384 471724
rect 49240 468512 49292 468518
rect 49240 468454 49292 468460
rect 49148 250504 49200 250510
rect 49148 250446 49200 250452
rect 49252 164665 49280 468454
rect 49344 166938 49372 471718
rect 49332 166932 49384 166938
rect 49332 166874 49384 166880
rect 49436 164694 49464 492118
rect 50988 492108 51040 492114
rect 50988 492050 51040 492056
rect 50896 491020 50948 491026
rect 50896 490962 50948 490968
rect 50908 490521 50936 490962
rect 50894 490512 50950 490521
rect 50894 490447 50950 490456
rect 50068 489932 50120 489938
rect 50068 489874 50120 489880
rect 49976 468444 50028 468450
rect 49976 468386 50028 468392
rect 49516 465860 49568 465866
rect 49516 465802 49568 465808
rect 49424 164688 49476 164694
rect 49238 164656 49294 164665
rect 49424 164630 49476 164636
rect 49238 164591 49294 164600
rect 49056 148640 49108 148646
rect 49056 148582 49108 148588
rect 48228 144628 48280 144634
rect 48228 144570 48280 144576
rect 41328 70372 41380 70378
rect 41328 70314 41380 70320
rect 49528 57662 49556 465802
rect 49608 465656 49660 465662
rect 49608 465598 49660 465604
rect 49620 57730 49648 465598
rect 49988 464710 50016 468386
rect 49976 464704 50028 464710
rect 49976 464646 50028 464652
rect 50080 58682 50108 489874
rect 50528 488232 50580 488238
rect 50528 488174 50580 488180
rect 50436 487756 50488 487762
rect 50436 487698 50488 487704
rect 50160 485308 50212 485314
rect 50160 485250 50212 485256
rect 50172 378690 50200 485250
rect 50344 482792 50396 482798
rect 50344 482734 50396 482740
rect 50252 474564 50304 474570
rect 50252 474506 50304 474512
rect 50160 378684 50212 378690
rect 50160 378626 50212 378632
rect 50264 271114 50292 474506
rect 50356 273057 50384 482734
rect 50342 273048 50398 273057
rect 50342 272983 50398 272992
rect 50252 271108 50304 271114
rect 50252 271050 50304 271056
rect 50356 163606 50384 272983
rect 50448 272678 50476 487698
rect 50540 273018 50568 488174
rect 51000 480254 51028 492050
rect 51908 492040 51960 492046
rect 51908 491982 51960 491988
rect 51816 487688 51868 487694
rect 51816 487630 51868 487636
rect 50908 480226 51028 480254
rect 50712 466404 50764 466410
rect 50712 466346 50764 466352
rect 50620 465724 50672 465730
rect 50620 465666 50672 465672
rect 50528 273012 50580 273018
rect 50528 272954 50580 272960
rect 50526 272912 50582 272921
rect 50526 272847 50582 272856
rect 50436 272672 50488 272678
rect 50436 272614 50488 272620
rect 50344 163600 50396 163606
rect 50344 163542 50396 163548
rect 50540 144838 50568 272847
rect 50632 165481 50660 465666
rect 50724 465225 50752 466346
rect 50804 465792 50856 465798
rect 50804 465734 50856 465740
rect 50710 465216 50766 465225
rect 50710 465151 50766 465160
rect 50712 464704 50764 464710
rect 50712 464646 50764 464652
rect 50724 166802 50752 464646
rect 50712 166796 50764 166802
rect 50712 166738 50764 166744
rect 50816 166258 50844 465734
rect 50804 166252 50856 166258
rect 50804 166194 50856 166200
rect 50618 165472 50674 165481
rect 50618 165407 50674 165416
rect 50908 164830 50936 480226
rect 51724 474632 51776 474638
rect 51724 474574 51776 474580
rect 51632 474496 51684 474502
rect 51632 474438 51684 474444
rect 50988 471980 51040 471986
rect 50988 471922 51040 471928
rect 51000 465798 51028 471922
rect 51540 465996 51592 466002
rect 51540 465938 51592 465944
rect 50988 465792 51040 465798
rect 50988 465734 51040 465740
rect 50988 272944 51040 272950
rect 50988 272886 51040 272892
rect 50896 164824 50948 164830
rect 50896 164766 50948 164772
rect 51000 163742 51028 272886
rect 50988 163736 51040 163742
rect 50988 163678 51040 163684
rect 50528 144832 50580 144838
rect 50528 144774 50580 144780
rect 50068 58676 50120 58682
rect 50068 58618 50120 58624
rect 49608 57724 49660 57730
rect 49608 57666 49660 57672
rect 49516 57656 49568 57662
rect 49516 57598 49568 57604
rect 51552 57390 51580 465938
rect 51644 410650 51672 474438
rect 51632 410644 51684 410650
rect 51632 410586 51684 410592
rect 51632 409896 51684 409902
rect 51632 409838 51684 409844
rect 51644 380730 51672 409838
rect 51632 380724 51684 380730
rect 51632 380666 51684 380672
rect 51630 272776 51686 272785
rect 51630 272711 51686 272720
rect 51644 144770 51672 272711
rect 51736 271250 51764 474574
rect 51828 272610 51856 487630
rect 51816 272604 51868 272610
rect 51816 272546 51868 272552
rect 51724 271244 51776 271250
rect 51724 271186 51776 271192
rect 51920 271182 51948 491982
rect 52276 490952 52328 490958
rect 52276 490894 52328 490900
rect 52092 471232 52144 471238
rect 52092 471174 52144 471180
rect 52000 468784 52052 468790
rect 52000 468726 52052 468732
rect 51908 271176 51960 271182
rect 51908 271118 51960 271124
rect 51724 270020 51776 270026
rect 51724 269962 51776 269968
rect 51736 269006 51764 269962
rect 51724 269000 51776 269006
rect 51724 268942 51776 268948
rect 51736 144906 51764 268942
rect 52012 164966 52040 468726
rect 52104 167006 52132 471174
rect 52184 464432 52236 464438
rect 52184 464374 52236 464380
rect 52196 380390 52224 464374
rect 52184 380384 52236 380390
rect 52184 380326 52236 380332
rect 52182 379536 52238 379545
rect 52182 379471 52238 379480
rect 52092 167000 52144 167006
rect 52092 166942 52144 166948
rect 52000 164960 52052 164966
rect 52000 164902 52052 164908
rect 52092 148776 52144 148782
rect 52092 148718 52144 148724
rect 52000 148708 52052 148714
rect 52000 148650 52052 148656
rect 51908 146260 51960 146266
rect 51908 146202 51960 146208
rect 51920 145518 51948 146202
rect 51908 145512 51960 145518
rect 51908 145454 51960 145460
rect 51724 144900 51776 144906
rect 51724 144842 51776 144848
rect 51632 144764 51684 144770
rect 51632 144706 51684 144712
rect 51540 57384 51592 57390
rect 51540 57326 51592 57332
rect 41236 56568 41288 56574
rect 41236 56510 41288 56516
rect 51920 55962 51948 145454
rect 52012 56030 52040 148650
rect 52000 56024 52052 56030
rect 52000 55966 52052 55972
rect 51908 55956 51960 55962
rect 51908 55898 51960 55904
rect 52104 54670 52132 148718
rect 52196 58818 52224 379471
rect 52288 166870 52316 490894
rect 53564 490884 53616 490890
rect 53564 490826 53616 490832
rect 53472 471912 53524 471918
rect 53472 471854 53524 471860
rect 53196 471504 53248 471510
rect 53196 471446 53248 471452
rect 52828 471436 52880 471442
rect 52828 471378 52880 471384
rect 52368 408536 52420 408542
rect 52368 408478 52420 408484
rect 52380 380662 52408 408478
rect 52460 389224 52512 389230
rect 52460 389166 52512 389172
rect 52472 388482 52500 389166
rect 52460 388476 52512 388482
rect 52460 388418 52512 388424
rect 52368 380656 52420 380662
rect 52368 380598 52420 380604
rect 52368 273284 52420 273290
rect 52368 273226 52420 273232
rect 52276 166864 52328 166870
rect 52276 166806 52328 166812
rect 52276 164212 52328 164218
rect 52276 164154 52328 164160
rect 52288 163674 52316 164154
rect 52276 163668 52328 163674
rect 52276 163610 52328 163616
rect 52184 58812 52236 58818
rect 52184 58754 52236 58760
rect 52288 56506 52316 163610
rect 52380 145625 52408 273226
rect 52460 271584 52512 271590
rect 52458 271552 52460 271561
rect 52512 271552 52514 271561
rect 52458 271487 52514 271496
rect 52734 271552 52790 271561
rect 52734 271487 52790 271496
rect 52748 163538 52776 271487
rect 52840 271454 52868 471378
rect 53012 464704 53064 464710
rect 53012 464646 53064 464652
rect 52920 410644 52972 410650
rect 52920 410586 52972 410592
rect 52828 271448 52880 271454
rect 52828 271390 52880 271396
rect 52932 271318 52960 410586
rect 53024 271522 53052 464646
rect 53012 271516 53064 271522
rect 53012 271458 53064 271464
rect 53208 271386 53236 471446
rect 53380 468648 53432 468654
rect 53380 468590 53432 468596
rect 53288 468580 53340 468586
rect 53288 468522 53340 468528
rect 53196 271380 53248 271386
rect 53196 271322 53248 271328
rect 52920 271312 52972 271318
rect 52920 271254 52972 271260
rect 53010 271144 53066 271153
rect 53010 271079 53066 271088
rect 53024 164014 53052 271079
rect 53104 269952 53156 269958
rect 53104 269894 53156 269900
rect 53116 269074 53144 269894
rect 53104 269068 53156 269074
rect 53104 269010 53156 269016
rect 53012 164008 53064 164014
rect 53012 163950 53064 163956
rect 52736 163532 52788 163538
rect 52736 163474 52788 163480
rect 52366 145616 52422 145625
rect 52366 145551 52422 145560
rect 52276 56500 52328 56506
rect 52276 56442 52328 56448
rect 53024 56438 53052 163950
rect 53116 161474 53144 269010
rect 53300 165345 53328 468522
rect 53286 165336 53342 165345
rect 53286 165271 53342 165280
rect 53392 165238 53420 468590
rect 53380 165232 53432 165238
rect 53380 165174 53432 165180
rect 53484 164082 53512 471854
rect 53576 165034 53604 490826
rect 53656 490476 53708 490482
rect 53656 490418 53708 490424
rect 53564 165028 53616 165034
rect 53564 164970 53616 164976
rect 53472 164076 53524 164082
rect 53472 164018 53524 164024
rect 53564 163600 53616 163606
rect 53564 163542 53616 163548
rect 53116 161446 53328 161474
rect 53196 148368 53248 148374
rect 53196 148310 53248 148316
rect 53208 58954 53236 148310
rect 53300 146062 53328 161446
rect 53380 148640 53432 148646
rect 53380 148582 53432 148588
rect 53288 146056 53340 146062
rect 53288 145998 53340 146004
rect 53196 58948 53248 58954
rect 53196 58890 53248 58896
rect 53012 56432 53064 56438
rect 53012 56374 53064 56380
rect 53300 56166 53328 145998
rect 53288 56160 53340 56166
rect 53288 56102 53340 56108
rect 53392 54738 53420 148582
rect 53576 55146 53604 163542
rect 53668 57798 53696 490418
rect 53760 389230 53788 521698
rect 302804 515545 302832 580858
rect 302896 572014 302924 590679
rect 302988 576298 303016 596663
rect 303066 584352 303122 584361
rect 303066 584287 303122 584296
rect 302976 576292 303028 576298
rect 302976 576234 303028 576240
rect 302884 572008 302936 572014
rect 302884 571950 302936 571956
rect 303080 569226 303108 584287
rect 303068 569220 303120 569226
rect 303068 569162 303120 569168
rect 304276 555286 304304 644846
rect 305644 644564 305696 644570
rect 305644 644506 305696 644512
rect 304356 556572 304408 556578
rect 304356 556514 304408 556520
rect 304264 555280 304316 555286
rect 304264 555222 304316 555228
rect 302882 554840 302938 554849
rect 302882 554775 302938 554784
rect 302896 531282 302924 554775
rect 303068 554328 303120 554334
rect 303068 554270 303120 554276
rect 302976 554124 303028 554130
rect 302976 554066 303028 554072
rect 302988 532506 303016 554066
rect 303080 539578 303108 554270
rect 304264 545148 304316 545154
rect 304264 545090 304316 545096
rect 303068 539572 303120 539578
rect 303068 539514 303120 539520
rect 302976 532500 303028 532506
rect 302976 532442 303028 532448
rect 302884 531276 302936 531282
rect 302884 531218 302936 531224
rect 302790 515536 302846 515545
rect 302790 515471 302846 515480
rect 302882 500576 302938 500585
rect 302882 500511 302938 500520
rect 302896 499594 302924 500511
rect 302884 499588 302936 499594
rect 302884 499530 302936 499536
rect 304276 494766 304304 545090
rect 304368 531894 304396 556514
rect 305656 555393 305684 644506
rect 305736 625184 305788 625190
rect 305736 625126 305788 625132
rect 305748 565214 305776 625126
rect 305828 596216 305880 596222
rect 305828 596158 305880 596164
rect 305840 580990 305868 596158
rect 305828 580984 305880 580990
rect 305828 580926 305880 580932
rect 305736 565208 305788 565214
rect 305736 565150 305788 565156
rect 305642 555384 305698 555393
rect 305642 555319 305698 555328
rect 305644 553988 305696 553994
rect 305644 553930 305696 553936
rect 305656 531962 305684 553930
rect 307036 532846 307064 700334
rect 364352 692102 364380 702406
rect 429856 700398 429884 703520
rect 429844 700392 429896 700398
rect 429844 700334 429896 700340
rect 434720 700392 434772 700398
rect 434720 700334 434772 700340
rect 364340 692096 364392 692102
rect 364340 692038 364392 692044
rect 427820 692096 427872 692102
rect 427820 692038 427872 692044
rect 427832 654134 427860 692038
rect 427832 654106 428320 654134
rect 405832 652044 405884 652050
rect 405832 651986 405884 651992
rect 324228 649324 324280 649330
rect 324228 649266 324280 649272
rect 311164 648168 311216 648174
rect 311164 648110 311216 648116
rect 309876 638988 309928 638994
rect 309876 638930 309928 638936
rect 307116 633480 307168 633486
rect 307116 633422 307168 633428
rect 307128 566574 307156 633422
rect 309784 629332 309836 629338
rect 309784 629274 309836 629280
rect 308404 600364 308456 600370
rect 308404 600306 308456 600312
rect 307116 566568 307168 566574
rect 307116 566510 307168 566516
rect 308416 556918 308444 600306
rect 308404 556912 308456 556918
rect 308404 556854 308456 556860
rect 307024 532840 307076 532846
rect 307024 532782 307076 532788
rect 305644 531956 305696 531962
rect 305644 531898 305696 531904
rect 304356 531888 304408 531894
rect 304356 531830 304408 531836
rect 304264 494760 304316 494766
rect 304264 494702 304316 494708
rect 59464 493054 60214 493082
rect 196298 493054 196664 493082
rect 59360 491496 59412 491502
rect 59360 491438 59412 491444
rect 59084 490816 59136 490822
rect 59084 490758 59136 490764
rect 55128 490748 55180 490754
rect 55128 490690 55180 490696
rect 54852 487620 54904 487626
rect 54852 487562 54904 487568
rect 54484 485580 54536 485586
rect 54484 485522 54536 485528
rect 54392 466200 54444 466206
rect 54392 466142 54444 466148
rect 54300 466064 54352 466070
rect 54300 466006 54352 466012
rect 53748 389224 53800 389230
rect 53748 389166 53800 389172
rect 53746 388512 53802 388521
rect 53746 388447 53802 388456
rect 53760 57866 53788 388447
rect 54312 378010 54340 466006
rect 54300 378004 54352 378010
rect 54300 377946 54352 377952
rect 54404 377942 54432 466142
rect 54496 379506 54524 485522
rect 54758 485480 54814 485489
rect 54758 485415 54814 485424
rect 54668 471572 54720 471578
rect 54668 471514 54720 471520
rect 54576 464568 54628 464574
rect 54576 464510 54628 464516
rect 54484 379500 54536 379506
rect 54484 379442 54536 379448
rect 54482 378040 54538 378049
rect 54482 377975 54538 377984
rect 54392 377936 54444 377942
rect 54392 377878 54444 377884
rect 54496 282198 54524 377975
rect 54484 282192 54536 282198
rect 54484 282134 54536 282140
rect 53840 273012 53892 273018
rect 53840 272954 53892 272960
rect 53852 272202 53880 272954
rect 54588 272921 54616 464510
rect 54574 272912 54630 272921
rect 54574 272847 54630 272856
rect 54300 272332 54352 272338
rect 54300 272274 54352 272280
rect 53840 272196 53892 272202
rect 53840 272138 53892 272144
rect 54116 272196 54168 272202
rect 54116 272138 54168 272144
rect 53840 251864 53892 251870
rect 53840 251806 53892 251812
rect 53852 251025 53880 251806
rect 53838 251016 53894 251025
rect 53838 250951 53894 250960
rect 54128 145994 54156 272138
rect 54208 271992 54260 271998
rect 54208 271934 54260 271940
rect 54220 146198 54248 271934
rect 54208 146192 54260 146198
rect 54208 146134 54260 146140
rect 54116 145988 54168 145994
rect 54116 145930 54168 145936
rect 54312 145926 54340 272274
rect 54680 271658 54708 471514
rect 54772 271998 54800 485415
rect 54864 272882 54892 487562
rect 55036 469056 55088 469062
rect 55036 468998 55088 469004
rect 54944 468852 54996 468858
rect 54944 468794 54996 468800
rect 54852 272876 54904 272882
rect 54852 272818 54904 272824
rect 54760 271992 54812 271998
rect 54760 271934 54812 271940
rect 54668 271652 54720 271658
rect 54668 271594 54720 271600
rect 54574 270600 54630 270609
rect 54574 270535 54630 270544
rect 54390 251016 54446 251025
rect 54390 250951 54446 250960
rect 54404 165646 54432 250951
rect 54392 165640 54444 165646
rect 54392 165582 54444 165588
rect 54300 145920 54352 145926
rect 54300 145862 54352 145868
rect 53748 57860 53800 57866
rect 53748 57802 53800 57808
rect 53656 57792 53708 57798
rect 53656 57734 53708 57740
rect 53564 55140 53616 55146
rect 53564 55082 53616 55088
rect 54404 55078 54432 165582
rect 54588 164218 54616 270535
rect 54852 250504 54904 250510
rect 54852 250446 54904 250452
rect 54576 164212 54628 164218
rect 54576 164154 54628 164160
rect 54760 145988 54812 145994
rect 54760 145930 54812 145936
rect 54484 145920 54536 145926
rect 54484 145862 54536 145868
rect 54496 59634 54524 145862
rect 54574 145616 54630 145625
rect 54574 145551 54630 145560
rect 54484 59628 54536 59634
rect 54484 59570 54536 59576
rect 54588 59566 54616 145551
rect 54668 145444 54720 145450
rect 54668 145386 54720 145392
rect 54680 59838 54708 145386
rect 54668 59832 54720 59838
rect 54668 59774 54720 59780
rect 54576 59560 54628 59566
rect 54576 59502 54628 59508
rect 54772 59362 54800 145930
rect 54864 145897 54892 250446
rect 54956 165374 54984 468794
rect 54944 165368 54996 165374
rect 54944 165310 54996 165316
rect 55048 165102 55076 468998
rect 55140 165510 55168 490690
rect 58532 490544 58584 490550
rect 58532 490486 58584 490492
rect 56324 490408 56376 490414
rect 56324 490350 56376 490356
rect 56336 490113 56364 490350
rect 56322 490104 56378 490113
rect 56322 490039 56378 490048
rect 56416 487892 56468 487898
rect 56416 487834 56468 487840
rect 56324 471844 56376 471850
rect 56324 471786 56376 471792
rect 56230 471336 56286 471345
rect 56230 471271 56286 471280
rect 56048 469192 56100 469198
rect 56048 469134 56100 469140
rect 55956 468988 56008 468994
rect 55956 468930 56008 468936
rect 55864 468920 55916 468926
rect 55864 468862 55916 468868
rect 55588 465928 55640 465934
rect 55588 465870 55640 465876
rect 55494 381032 55550 381041
rect 55494 380967 55550 380976
rect 55128 165504 55180 165510
rect 55128 165446 55180 165452
rect 55036 165096 55088 165102
rect 55036 165038 55088 165044
rect 55036 163736 55088 163742
rect 55036 163678 55088 163684
rect 54944 148436 54996 148442
rect 54944 148378 54996 148384
rect 54850 145888 54906 145897
rect 54850 145823 54906 145832
rect 54852 145376 54904 145382
rect 54852 145318 54904 145324
rect 54760 59356 54812 59362
rect 54760 59298 54812 59304
rect 54864 57186 54892 145318
rect 54852 57180 54904 57186
rect 54852 57122 54904 57128
rect 54956 55214 54984 148378
rect 55048 59226 55076 163678
rect 55036 59220 55088 59226
rect 55036 59162 55088 59168
rect 55508 58750 55536 380967
rect 55600 58886 55628 465870
rect 55772 464636 55824 464642
rect 55772 464578 55824 464584
rect 55784 380934 55812 464578
rect 55772 380928 55824 380934
rect 55772 380870 55824 380876
rect 55772 357400 55824 357406
rect 55772 357342 55824 357348
rect 55784 272474 55812 357342
rect 55772 272468 55824 272474
rect 55772 272410 55824 272416
rect 55772 268728 55824 268734
rect 55772 268670 55824 268676
rect 55680 164144 55732 164150
rect 55680 164086 55732 164092
rect 55692 96626 55720 164086
rect 55784 146266 55812 268670
rect 55876 165578 55904 468862
rect 55864 165572 55916 165578
rect 55864 165514 55916 165520
rect 55968 165442 55996 468930
rect 55956 165436 56008 165442
rect 55956 165378 56008 165384
rect 56060 164626 56088 469134
rect 56140 469124 56192 469130
rect 56140 469066 56192 469072
rect 56152 165306 56180 469066
rect 56244 166734 56272 471271
rect 56232 166728 56284 166734
rect 56232 166670 56284 166676
rect 56140 165300 56192 165306
rect 56140 165242 56192 165248
rect 56336 165209 56364 471786
rect 56428 378826 56456 487834
rect 57152 485784 57204 485790
rect 57152 485726 57204 485732
rect 56876 471640 56928 471646
rect 56876 471582 56928 471588
rect 56692 471368 56744 471374
rect 56692 471310 56744 471316
rect 56508 392012 56560 392018
rect 56508 391954 56560 391960
rect 56520 380458 56548 391954
rect 56508 380452 56560 380458
rect 56508 380394 56560 380400
rect 56416 378820 56468 378826
rect 56416 378762 56468 378768
rect 56704 311137 56732 471310
rect 56784 388544 56836 388550
rect 56784 388486 56836 388492
rect 56690 311128 56746 311137
rect 56690 311063 56746 311072
rect 56508 270156 56560 270162
rect 56508 270098 56560 270104
rect 56520 268734 56548 270098
rect 56508 268728 56560 268734
rect 56508 268670 56560 268676
rect 56690 204232 56746 204241
rect 56690 204167 56746 204176
rect 56704 203017 56732 204167
rect 56690 203008 56746 203017
rect 56690 202943 56746 202952
rect 56322 165200 56378 165209
rect 56322 165135 56378 165144
rect 56048 164620 56100 164626
rect 56048 164562 56100 164568
rect 56048 148572 56100 148578
rect 56048 148514 56100 148520
rect 55772 146260 55824 146266
rect 55772 146202 55824 146208
rect 55956 144900 56008 144906
rect 55956 144842 56008 144848
rect 55864 144832 55916 144838
rect 55864 144774 55916 144780
rect 55680 96620 55732 96626
rect 55680 96562 55732 96568
rect 55876 59702 55904 144774
rect 55968 59770 55996 144842
rect 55956 59764 56008 59770
rect 55956 59706 56008 59712
rect 55864 59696 55916 59702
rect 55864 59638 55916 59644
rect 56060 59498 56088 148514
rect 56140 147688 56192 147694
rect 56140 147630 56192 147636
rect 56048 59492 56100 59498
rect 56048 59434 56100 59440
rect 56152 59090 56180 147630
rect 56232 146260 56284 146266
rect 56232 146202 56284 146208
rect 56244 145314 56272 146202
rect 56324 146192 56376 146198
rect 56324 146134 56376 146140
rect 56336 145790 56364 146134
rect 56416 145852 56468 145858
rect 56416 145794 56468 145800
rect 56324 145784 56376 145790
rect 56324 145726 56376 145732
rect 56232 145308 56284 145314
rect 56232 145250 56284 145256
rect 56140 59084 56192 59090
rect 56140 59026 56192 59032
rect 55588 58880 55640 58886
rect 55588 58822 55640 58828
rect 55496 58744 55548 58750
rect 55496 58686 55548 58692
rect 54944 55208 54996 55214
rect 54944 55150 54996 55156
rect 54392 55072 54444 55078
rect 54392 55014 54444 55020
rect 56244 54806 56272 145250
rect 56336 54874 56364 145726
rect 56428 144906 56456 145794
rect 56506 145752 56562 145761
rect 56506 145687 56562 145696
rect 56416 144900 56468 144906
rect 56416 144842 56468 144848
rect 56520 144838 56548 145687
rect 56508 144832 56560 144838
rect 56508 144774 56560 144780
rect 56704 96529 56732 202943
rect 56796 175137 56824 388486
rect 56888 271590 56916 471582
rect 57060 464500 57112 464506
rect 57060 464442 57112 464448
rect 57072 392018 57100 464442
rect 57060 392012 57112 392018
rect 57060 391954 57112 391960
rect 57164 390674 57192 485726
rect 57888 485512 57940 485518
rect 57888 485454 57940 485460
rect 57704 482996 57756 483002
rect 57704 482938 57756 482944
rect 57612 472660 57664 472666
rect 57612 472602 57664 472608
rect 57520 469872 57572 469878
rect 57520 469814 57572 469820
rect 57336 468716 57388 468722
rect 57336 468658 57388 468664
rect 57244 418056 57296 418062
rect 57244 417998 57296 418004
rect 57256 417625 57284 417998
rect 57242 417616 57298 417625
rect 57242 417551 57298 417560
rect 57072 390646 57192 390674
rect 57072 388482 57100 390646
rect 57152 390584 57204 390590
rect 57152 390526 57204 390532
rect 57060 388476 57112 388482
rect 57060 388418 57112 388424
rect 57164 388006 57192 390526
rect 57244 389156 57296 389162
rect 57244 389098 57296 389104
rect 57256 389065 57284 389098
rect 57242 389056 57298 389065
rect 57242 388991 57298 389000
rect 57152 388000 57204 388006
rect 57152 387942 57204 387948
rect 57060 380928 57112 380934
rect 57060 380870 57112 380876
rect 56966 301608 57022 301617
rect 56966 301543 57022 301552
rect 56980 300830 57008 301543
rect 57072 300830 57100 380870
rect 57150 310448 57206 310457
rect 57150 310383 57206 310392
rect 56968 300824 57020 300830
rect 56968 300766 57020 300772
rect 57060 300824 57112 300830
rect 57060 300766 57112 300772
rect 56876 271584 56928 271590
rect 56876 271526 56928 271532
rect 56876 269816 56928 269822
rect 56876 269758 56928 269764
rect 56888 268870 56916 269758
rect 56876 268864 56928 268870
rect 56876 268806 56928 268812
rect 56782 175128 56838 175137
rect 56782 175063 56838 175072
rect 56888 165170 56916 268806
rect 56980 195265 57008 300766
rect 57164 204241 57192 310383
rect 57348 306785 57376 468658
rect 57428 467220 57480 467226
rect 57428 467162 57480 467168
rect 57440 389450 57468 467162
rect 57532 389586 57560 469814
rect 57624 389722 57652 472602
rect 57716 402974 57744 482938
rect 57796 418124 57848 418130
rect 57796 418066 57848 418072
rect 57808 417897 57836 418066
rect 57794 417888 57850 417897
rect 57794 417823 57850 417832
rect 57794 414216 57850 414225
rect 57794 414151 57850 414160
rect 57808 414050 57836 414151
rect 57796 414044 57848 414050
rect 57796 413986 57848 413992
rect 57794 413264 57850 413273
rect 57794 413199 57850 413208
rect 57808 412690 57836 413199
rect 57796 412684 57848 412690
rect 57796 412626 57848 412632
rect 57794 411496 57850 411505
rect 57794 411431 57850 411440
rect 57808 411330 57836 411431
rect 57796 411324 57848 411330
rect 57796 411266 57848 411272
rect 57794 410408 57850 410417
rect 57794 410343 57850 410352
rect 57808 409902 57836 410343
rect 57796 409896 57848 409902
rect 57796 409838 57848 409844
rect 57794 408640 57850 408649
rect 57794 408575 57850 408584
rect 57808 408542 57836 408575
rect 57796 408536 57848 408542
rect 57796 408478 57848 408484
rect 57716 402946 57836 402974
rect 57704 391944 57756 391950
rect 57704 391886 57756 391892
rect 57716 391649 57744 391886
rect 57702 391640 57758 391649
rect 57702 391575 57758 391584
rect 57624 389694 57744 389722
rect 57532 389558 57652 389586
rect 57440 389422 57560 389450
rect 57426 389328 57482 389337
rect 57426 389263 57482 389272
rect 57440 389230 57468 389263
rect 57428 389224 57480 389230
rect 57428 389166 57480 389172
rect 57532 388498 57560 389422
rect 57440 388470 57560 388498
rect 57334 306776 57390 306785
rect 57334 306711 57390 306720
rect 57244 281512 57296 281518
rect 57244 281454 57296 281460
rect 57150 204232 57206 204241
rect 57150 204167 57206 204176
rect 57058 203960 57114 203969
rect 57058 203895 57114 203904
rect 56966 195256 57022 195265
rect 56966 195191 57022 195200
rect 56876 165164 56928 165170
rect 56876 165106 56928 165112
rect 56968 144696 57020 144702
rect 56968 144638 57020 144644
rect 56690 96520 56746 96529
rect 56690 96455 56746 96464
rect 56980 55010 57008 144638
rect 57072 97481 57100 203895
rect 57150 198792 57206 198801
rect 57150 198727 57206 198736
rect 57058 97472 57114 97481
rect 57058 97407 57114 97416
rect 57060 96620 57112 96626
rect 57060 96562 57112 96568
rect 57072 57594 57100 96562
rect 57164 93401 57192 198727
rect 57256 175409 57284 281454
rect 57348 199889 57376 306711
rect 57440 303929 57468 388470
rect 57624 388362 57652 389558
rect 57532 388334 57652 388362
rect 57532 305017 57560 388334
rect 57716 388226 57744 389694
rect 57624 388198 57744 388226
rect 57624 307873 57652 388198
rect 57808 388090 57836 402946
rect 57716 388062 57836 388090
rect 57716 310457 57744 388062
rect 57796 388000 57848 388006
rect 57796 387942 57848 387948
rect 57808 382090 57836 387942
rect 57796 382084 57848 382090
rect 57796 382026 57848 382032
rect 57900 380254 57928 485454
rect 58440 482860 58492 482866
rect 58440 482802 58492 482808
rect 58346 390688 58402 390697
rect 58346 390623 58402 390632
rect 58360 380934 58388 390623
rect 58452 390590 58480 482802
rect 58440 390584 58492 390590
rect 58440 390526 58492 390532
rect 58544 388550 58572 490486
rect 58624 485716 58676 485722
rect 58624 485658 58676 485664
rect 58532 388544 58584 388550
rect 58532 388486 58584 388492
rect 58440 388476 58492 388482
rect 58440 388418 58492 388424
rect 58348 380928 58400 380934
rect 58348 380870 58400 380876
rect 57888 380248 57940 380254
rect 57888 380190 57940 380196
rect 58452 378894 58480 388418
rect 58636 378962 58664 485658
rect 58808 484900 58860 484906
rect 58808 484842 58860 484848
rect 58716 483676 58768 483682
rect 58716 483618 58768 483624
rect 58624 378956 58676 378962
rect 58624 378898 58676 378904
rect 58440 378888 58492 378894
rect 58440 378830 58492 378836
rect 58624 356040 58676 356046
rect 58624 355982 58676 355988
rect 57886 311128 57942 311137
rect 57886 311063 57942 311072
rect 57702 310448 57758 310457
rect 57702 310383 57758 310392
rect 57610 307864 57666 307873
rect 57610 307799 57666 307808
rect 57518 305008 57574 305017
rect 57518 304943 57574 304952
rect 57426 303920 57482 303929
rect 57426 303855 57482 303864
rect 57334 199880 57390 199889
rect 57334 199815 57390 199824
rect 57348 198801 57376 199815
rect 57334 198792 57390 198801
rect 57334 198727 57390 198736
rect 57440 196353 57468 303855
rect 57532 282418 57560 304943
rect 57624 287054 57652 307799
rect 57624 287026 57744 287054
rect 57532 282390 57652 282418
rect 57518 282296 57574 282305
rect 57518 282231 57574 282240
rect 57532 281518 57560 282231
rect 57520 281512 57572 281518
rect 57520 281454 57572 281460
rect 57624 281330 57652 282390
rect 57532 281302 57652 281330
rect 57532 197441 57560 281302
rect 57716 277394 57744 287026
rect 57624 277366 57744 277394
rect 57624 200841 57652 277366
rect 57900 203969 57928 311063
rect 58532 300824 58584 300830
rect 58532 300766 58584 300772
rect 57980 282192 58032 282198
rect 57980 282134 58032 282140
rect 57992 273290 58020 282134
rect 57980 273284 58032 273290
rect 57980 273226 58032 273232
rect 58544 271930 58572 300766
rect 58636 277394 58664 355982
rect 58728 282033 58756 483618
rect 58820 284209 58848 484842
rect 58900 471708 58952 471714
rect 58900 471650 58952 471656
rect 58806 284200 58862 284209
rect 58806 284135 58862 284144
rect 58714 282024 58770 282033
rect 58714 281959 58770 281968
rect 58636 277366 58756 277394
rect 58532 271924 58584 271930
rect 58532 271866 58584 271872
rect 58544 270314 58572 271866
rect 58728 270609 58756 277366
rect 58808 273284 58860 273290
rect 58808 273226 58860 273232
rect 58820 272814 58848 273226
rect 58808 272808 58860 272814
rect 58808 272750 58860 272756
rect 58714 270600 58770 270609
rect 58714 270535 58770 270544
rect 58728 270434 58756 270535
rect 58716 270428 58768 270434
rect 58716 270370 58768 270376
rect 58544 270286 58848 270314
rect 58624 270224 58676 270230
rect 58624 270166 58676 270172
rect 57980 269884 58032 269890
rect 57980 269826 58032 269832
rect 57992 268258 58020 269826
rect 58636 268802 58664 270166
rect 58624 268796 58676 268802
rect 58624 268738 58676 268744
rect 57980 268252 58032 268258
rect 57980 268194 58032 268200
rect 57886 203960 57942 203969
rect 57886 203895 57942 203904
rect 57610 200832 57666 200841
rect 57610 200767 57666 200776
rect 57518 197432 57574 197441
rect 57518 197367 57574 197376
rect 57426 196344 57482 196353
rect 57426 196279 57482 196288
rect 57242 175400 57298 175409
rect 57242 175335 57298 175344
rect 57336 165164 57388 165170
rect 57336 165106 57388 165112
rect 57348 164898 57376 165106
rect 57336 164892 57388 164898
rect 57336 164834 57388 164840
rect 57150 93392 57206 93401
rect 57150 93327 57206 93336
rect 57348 59022 57376 164834
rect 57440 90545 57468 196279
rect 57520 164212 57572 164218
rect 57520 164154 57572 164160
rect 57532 163305 57560 164154
rect 57518 163296 57574 163305
rect 57518 163231 57574 163240
rect 57520 145716 57572 145722
rect 57520 145658 57572 145664
rect 57532 144702 57560 145658
rect 57520 144696 57572 144702
rect 57520 144638 57572 144644
rect 57624 93809 57652 200767
rect 57702 197432 57758 197441
rect 57702 197367 57758 197376
rect 57610 93800 57666 93809
rect 57610 93735 57666 93744
rect 57716 91089 57744 197367
rect 57794 195256 57850 195265
rect 57794 195191 57850 195200
rect 57702 91080 57758 91089
rect 57702 91015 57758 91024
rect 57426 90536 57482 90545
rect 57426 90471 57482 90480
rect 57808 88233 57836 195191
rect 57886 175400 57942 175409
rect 57886 175335 57942 175344
rect 57794 88224 57850 88233
rect 57794 88159 57850 88168
rect 57520 70372 57572 70378
rect 57520 70314 57572 70320
rect 57532 70145 57560 70314
rect 57518 70136 57574 70145
rect 57518 70071 57574 70080
rect 57900 68921 57928 175335
rect 57992 149054 58020 268194
rect 58532 252000 58584 252006
rect 58532 251942 58584 251948
rect 58544 251161 58572 251942
rect 58530 251152 58586 251161
rect 58530 251087 58586 251096
rect 57980 149048 58032 149054
rect 57980 148990 58032 148996
rect 57992 147694 58020 148990
rect 58544 148510 58572 251087
rect 58532 148504 58584 148510
rect 58532 148446 58584 148452
rect 58532 148300 58584 148306
rect 58532 148242 58584 148248
rect 57980 147688 58032 147694
rect 57980 147630 58032 147636
rect 58544 146112 58572 148242
rect 58636 146266 58664 268738
rect 58716 252068 58768 252074
rect 58716 252010 58768 252016
rect 58624 146260 58676 146266
rect 58624 146202 58676 146208
rect 58728 146198 58756 252010
rect 58820 148986 58848 270286
rect 58912 177585 58940 471650
rect 58992 464772 59044 464778
rect 58992 464714 59044 464720
rect 58898 177576 58954 177585
rect 58898 177511 58954 177520
rect 59004 166462 59032 464714
rect 59096 166598 59124 490758
rect 59372 487966 59400 491438
rect 59464 489190 59492 493054
rect 60292 493023 60582 493051
rect 60292 491502 60320 493023
rect 60280 491496 60332 491502
rect 60280 491438 60332 491444
rect 59452 489184 59504 489190
rect 59452 489126 59504 489132
rect 59728 488436 59780 488442
rect 59728 488378 59780 488384
rect 59360 487960 59412 487966
rect 59360 487902 59412 487908
rect 59636 482928 59688 482934
rect 59636 482870 59688 482876
rect 59268 467084 59320 467090
rect 59268 467026 59320 467032
rect 59176 466132 59228 466138
rect 59176 466074 59228 466080
rect 59084 166592 59136 166598
rect 59084 166534 59136 166540
rect 58992 166456 59044 166462
rect 58992 166398 59044 166404
rect 59084 163804 59136 163810
rect 59084 163746 59136 163752
rect 59096 163538 59124 163746
rect 59084 163532 59136 163538
rect 59084 163474 59136 163480
rect 58808 148980 58860 148986
rect 58808 148922 58860 148928
rect 58820 148578 58848 148922
rect 58808 148572 58860 148578
rect 58808 148514 58860 148520
rect 58992 148572 59044 148578
rect 58992 148514 59044 148520
rect 59004 148306 59032 148514
rect 58992 148300 59044 148306
rect 58992 148242 59044 148248
rect 58900 146260 58952 146266
rect 58900 146202 58952 146208
rect 58992 146260 59044 146266
rect 58992 146202 59044 146208
rect 58716 146192 58768 146198
rect 58716 146134 58768 146140
rect 58544 146084 58664 146112
rect 58530 146024 58586 146033
rect 58530 145959 58586 145968
rect 58544 145738 58572 145959
rect 58636 145874 58664 146084
rect 58636 145846 58848 145874
rect 58544 145710 58756 145738
rect 58624 145580 58676 145586
rect 58624 145522 58676 145528
rect 58636 144770 58664 145522
rect 58624 144764 58676 144770
rect 58624 144706 58676 144712
rect 57886 68912 57942 68921
rect 57886 68847 57942 68856
rect 57336 59016 57388 59022
rect 57336 58958 57388 58964
rect 57900 57934 57928 68847
rect 57244 57928 57296 57934
rect 57244 57870 57296 57876
rect 57888 57928 57940 57934
rect 57888 57870 57940 57876
rect 57060 57588 57112 57594
rect 57060 57530 57112 57536
rect 56968 55004 57020 55010
rect 56968 54946 57020 54952
rect 56324 54868 56376 54874
rect 56324 54810 56376 54816
rect 56232 54800 56284 54806
rect 56232 54742 56284 54748
rect 53380 54732 53432 54738
rect 53380 54674 53432 54680
rect 52092 54664 52144 54670
rect 52092 54606 52144 54612
rect 2780 20392 2832 20398
rect 2780 20334 2832 20340
rect 4804 20392 4856 20398
rect 4804 20334 4856 20340
rect 2792 19417 2820 20334
rect 2778 19408 2834 19417
rect 2778 19343 2834 19352
rect 57256 3466 57284 57870
rect 58636 56370 58664 144706
rect 58728 144634 58756 145710
rect 58716 144628 58768 144634
rect 58716 144570 58768 144576
rect 58624 56364 58676 56370
rect 58624 56306 58676 56312
rect 58728 56234 58756 144570
rect 58820 59430 58848 145846
rect 58808 59424 58860 59430
rect 58808 59366 58860 59372
rect 58716 56228 58768 56234
rect 58716 56170 58768 56176
rect 58912 56098 58940 146202
rect 58900 56092 58952 56098
rect 58900 56034 58952 56040
rect 59004 54942 59032 146202
rect 59096 59294 59124 163474
rect 59084 59288 59136 59294
rect 59084 59230 59136 59236
rect 59188 57322 59216 466074
rect 59176 57316 59228 57322
rect 59176 57258 59228 57264
rect 59280 57254 59308 467026
rect 59360 382084 59412 382090
rect 59360 382026 59412 382032
rect 59372 357377 59400 382026
rect 59358 357368 59414 357377
rect 59358 357303 59414 357312
rect 59648 356046 59676 482870
rect 59636 356040 59688 356046
rect 59636 355982 59688 355988
rect 59634 272640 59690 272649
rect 59634 272575 59690 272584
rect 59648 272474 59676 272575
rect 59740 272474 59768 488378
rect 59910 471472 59966 471481
rect 59910 471407 59966 471416
rect 59820 465656 59872 465662
rect 59820 465598 59872 465604
rect 59636 272468 59688 272474
rect 59636 272410 59688 272416
rect 59728 272468 59780 272474
rect 59728 272410 59780 272416
rect 59360 270088 59412 270094
rect 59360 270030 59412 270036
rect 59372 268938 59400 270030
rect 59360 268932 59412 268938
rect 59360 268874 59412 268880
rect 59372 146266 59400 268874
rect 59450 164248 59506 164257
rect 59450 164183 59506 164192
rect 59464 163538 59492 164183
rect 59648 164150 59676 272410
rect 59832 166666 59860 465598
rect 59820 166660 59872 166666
rect 59820 166602 59872 166608
rect 59924 166530 59952 471407
rect 60004 468308 60056 468314
rect 60004 468250 60056 468256
rect 59912 166524 59964 166530
rect 59912 166466 59964 166472
rect 59820 165164 59872 165170
rect 59820 165106 59872 165112
rect 59832 164966 59860 165106
rect 59820 164960 59872 164966
rect 59820 164902 59872 164908
rect 59912 164960 59964 164966
rect 59912 164902 59964 164908
rect 59924 164830 59952 164902
rect 59912 164824 59964 164830
rect 59912 164766 59964 164772
rect 59636 164144 59688 164150
rect 59636 164086 59688 164092
rect 59452 163532 59504 163538
rect 59452 163474 59504 163480
rect 59360 146260 59412 146266
rect 59360 146202 59412 146208
rect 59464 140865 59492 163474
rect 59912 148844 59964 148850
rect 59912 148786 59964 148792
rect 59820 148504 59872 148510
rect 59820 148446 59872 148452
rect 59636 146192 59688 146198
rect 59636 146134 59688 146140
rect 59648 145654 59676 146134
rect 59636 145648 59688 145654
rect 59636 145590 59688 145596
rect 59648 142154 59676 145590
rect 59648 142126 59768 142154
rect 59450 140856 59506 140865
rect 59450 140791 59506 140800
rect 59268 57248 59320 57254
rect 59268 57190 59320 57196
rect 59740 56302 59768 142126
rect 59832 59158 59860 148446
rect 59820 59152 59872 59158
rect 59820 59094 59872 59100
rect 59924 57526 59952 148786
rect 59912 57520 59964 57526
rect 59912 57462 59964 57468
rect 60016 57458 60044 468250
rect 61028 467566 61056 493037
rect 61488 474026 61516 493037
rect 61948 475386 61976 493037
rect 61936 475380 61988 475386
rect 61936 475322 61988 475328
rect 61476 474020 61528 474026
rect 61476 473962 61528 473968
rect 61016 467560 61068 467566
rect 61016 467502 61068 467508
rect 62316 467498 62344 493037
rect 62776 476814 62804 493037
rect 62856 491156 62908 491162
rect 62856 491098 62908 491104
rect 62764 476808 62816 476814
rect 62764 476750 62816 476756
rect 62304 467492 62356 467498
rect 62304 467434 62356 467440
rect 62868 465662 62896 491098
rect 63236 466206 63264 493037
rect 63224 466200 63276 466206
rect 63224 466142 63276 466148
rect 63696 466070 63724 493037
rect 64156 491298 64184 493037
rect 64144 491292 64196 491298
rect 64144 491234 64196 491240
rect 64524 468382 64552 493037
rect 64984 471102 65012 493037
rect 65444 471170 65472 493037
rect 65904 471753 65932 493037
rect 66364 490657 66392 493037
rect 66350 490648 66406 490657
rect 66350 490583 66406 490592
rect 65890 471744 65946 471753
rect 65890 471679 65946 471688
rect 65432 471164 65484 471170
rect 65432 471106 65484 471112
rect 64972 471096 65024 471102
rect 64972 471038 65024 471044
rect 64512 468376 64564 468382
rect 64512 468318 64564 468324
rect 63684 466064 63736 466070
rect 63684 466006 63736 466012
rect 66732 466002 66760 493037
rect 67192 467090 67220 493037
rect 67180 467084 67232 467090
rect 67180 467026 67232 467032
rect 67652 466138 67680 493037
rect 67732 490000 67784 490006
rect 67732 489942 67784 489948
rect 67744 468314 67772 489942
rect 67732 468308 67784 468314
rect 67732 468250 67784 468256
rect 68112 467129 68140 493037
rect 68204 493023 68494 493051
rect 68664 493023 68954 493051
rect 68204 490006 68232 493023
rect 68284 491224 68336 491230
rect 68284 491166 68336 491172
rect 68192 490000 68244 490006
rect 68192 489942 68244 489948
rect 68296 467430 68324 491166
rect 68664 490385 68692 493023
rect 68928 491020 68980 491026
rect 68928 490962 68980 490968
rect 68940 490657 68968 490962
rect 68926 490648 68982 490657
rect 68926 490583 68982 490592
rect 68650 490376 68706 490385
rect 68376 490340 68428 490346
rect 68650 490311 68706 490320
rect 68376 490282 68428 490288
rect 68388 468450 68416 490282
rect 68376 468444 68428 468450
rect 68376 468386 68428 468392
rect 68284 467424 68336 467430
rect 68284 467366 68336 467372
rect 68098 467120 68154 467129
rect 68098 467055 68154 467064
rect 67640 466132 67692 466138
rect 67640 466074 67692 466080
rect 66720 465996 66772 466002
rect 66720 465938 66772 465944
rect 62856 465656 62908 465662
rect 69400 465633 69428 493037
rect 69860 469849 69888 493037
rect 69846 469840 69902 469849
rect 69846 469775 69902 469784
rect 70320 468761 70348 493037
rect 70688 468897 70716 493037
rect 70674 468888 70730 468897
rect 70674 468823 70730 468832
rect 70306 468752 70362 468761
rect 70306 468687 70362 468696
rect 71148 465866 71176 493037
rect 71608 491201 71636 493037
rect 71594 491192 71650 491201
rect 71594 491127 71650 491136
rect 71778 491192 71834 491201
rect 71778 491127 71834 491136
rect 71792 490414 71820 491127
rect 72068 490929 72096 493037
rect 72160 493023 72542 493051
rect 72054 490920 72110 490929
rect 72054 490855 72110 490864
rect 71780 490408 71832 490414
rect 71780 490350 71832 490356
rect 72160 489914 72188 493023
rect 72424 491088 72476 491094
rect 72238 491056 72294 491065
rect 72424 491030 72476 491036
rect 72238 490991 72294 491000
rect 72252 489938 72280 490991
rect 71792 489886 72188 489914
rect 72240 489932 72292 489938
rect 71136 465860 71188 465866
rect 71136 465802 71188 465808
rect 71792 465730 71820 489886
rect 72240 489874 72292 489880
rect 72436 473958 72464 491030
rect 72516 491020 72568 491026
rect 72516 490962 72568 490968
rect 72528 474706 72556 490962
rect 72516 474700 72568 474706
rect 72516 474642 72568 474648
rect 72424 473952 72476 473958
rect 72424 473894 72476 473900
rect 72896 467362 72924 493037
rect 73356 490249 73384 493037
rect 73816 490793 73844 493037
rect 73802 490784 73858 490793
rect 73802 490719 73858 490728
rect 74276 490482 74304 493037
rect 74644 490521 74672 493037
rect 74630 490512 74686 490521
rect 74264 490476 74316 490482
rect 74630 490447 74686 490456
rect 74264 490418 74316 490424
rect 73342 490240 73398 490249
rect 73342 490175 73398 490184
rect 72884 467356 72936 467362
rect 72884 467298 72936 467304
rect 75104 466449 75132 493037
rect 75090 466440 75146 466449
rect 75090 466375 75146 466384
rect 75564 465934 75592 493037
rect 76024 466313 76052 493037
rect 76010 466304 76066 466313
rect 76010 466239 76066 466248
rect 76484 466041 76512 493037
rect 76852 466177 76880 493037
rect 77312 491065 77340 493037
rect 77772 491201 77800 493037
rect 77758 491192 77814 491201
rect 77758 491127 77814 491136
rect 77298 491056 77354 491065
rect 77298 490991 77354 491000
rect 76838 466168 76894 466177
rect 76838 466103 76894 466112
rect 76470 466032 76526 466041
rect 76470 465967 76526 465976
rect 75552 465928 75604 465934
rect 78232 465905 78260 493037
rect 78692 490657 78720 493037
rect 78678 490648 78734 490657
rect 78678 490583 78734 490592
rect 75552 465870 75604 465876
rect 78218 465896 78274 465905
rect 78218 465831 78274 465840
rect 79060 465769 79088 493037
rect 79520 466410 79548 493037
rect 79980 468625 80008 493037
rect 79966 468616 80022 468625
rect 79966 468551 80022 468560
rect 80440 468489 80468 493037
rect 80808 485625 80836 493037
rect 81268 490550 81296 493037
rect 81256 490544 81308 490550
rect 81256 490486 81308 490492
rect 80794 485616 80850 485625
rect 80794 485551 80850 485560
rect 81728 469198 81756 493037
rect 82188 492182 82216 493037
rect 82176 492176 82228 492182
rect 82176 492118 82228 492124
rect 82648 471209 82676 493037
rect 83016 471986 83044 493037
rect 83004 471980 83056 471986
rect 83004 471922 83056 471928
rect 83476 471782 83504 493037
rect 83464 471776 83516 471782
rect 83464 471718 83516 471724
rect 83936 471238 83964 493037
rect 84396 492114 84424 493037
rect 84384 492108 84436 492114
rect 84384 492050 84436 492056
rect 84856 490958 84884 493037
rect 84844 490952 84896 490958
rect 84844 490894 84896 490900
rect 85224 490346 85252 493037
rect 85212 490340 85264 490346
rect 85212 490282 85264 490288
rect 85684 471918 85712 493037
rect 86144 490890 86172 493037
rect 86224 491292 86276 491298
rect 86224 491234 86276 491240
rect 86132 490884 86184 490890
rect 86132 490826 86184 490832
rect 85672 471912 85724 471918
rect 85672 471854 85724 471860
rect 83924 471232 83976 471238
rect 82634 471200 82690 471209
rect 83924 471174 83976 471180
rect 82634 471135 82690 471144
rect 81716 469192 81768 469198
rect 81716 469134 81768 469140
rect 80426 468480 80482 468489
rect 80426 468415 80482 468424
rect 79508 466404 79560 466410
rect 79508 466346 79560 466352
rect 79046 465760 79102 465769
rect 71780 465724 71832 465730
rect 86236 465730 86264 491234
rect 86604 468790 86632 493037
rect 87064 469062 87092 493037
rect 87052 469056 87104 469062
rect 87052 468998 87104 469004
rect 86592 468784 86644 468790
rect 86592 468726 86644 468732
rect 87432 468654 87460 493037
rect 87892 469130 87920 493037
rect 87880 469124 87932 469130
rect 87880 469066 87932 469072
rect 88352 468858 88380 493037
rect 88812 468994 88840 493037
rect 89180 490754 89208 493037
rect 89168 490748 89220 490754
rect 89168 490690 89220 490696
rect 88800 468988 88852 468994
rect 88800 468930 88852 468936
rect 89640 468926 89668 493037
rect 90100 471850 90128 493037
rect 90088 471844 90140 471850
rect 90088 471786 90140 471792
rect 90560 471345 90588 493037
rect 91020 471617 91048 493037
rect 91388 491162 91416 493037
rect 91376 491156 91428 491162
rect 91376 491098 91428 491104
rect 91848 490822 91876 493037
rect 91836 490816 91888 490822
rect 91836 490758 91888 490764
rect 91006 471608 91062 471617
rect 91006 471543 91062 471552
rect 90546 471336 90602 471345
rect 90546 471271 90602 471280
rect 89628 468920 89680 468926
rect 89628 468862 89680 468868
rect 88340 468852 88392 468858
rect 88340 468794 88392 468800
rect 87420 468648 87472 468654
rect 87420 468590 87472 468596
rect 79046 465695 79102 465704
rect 86224 465724 86276 465730
rect 71780 465666 71832 465672
rect 86224 465666 86276 465672
rect 62856 465598 62908 465604
rect 69386 465624 69442 465633
rect 69386 465559 69442 465568
rect 92308 464409 92336 493037
rect 92768 471481 92796 493037
rect 92754 471472 92810 471481
rect 92754 471407 92810 471416
rect 93228 464778 93256 493037
rect 93596 465798 93624 493037
rect 94056 468586 94084 493037
rect 94044 468580 94096 468586
rect 94044 468522 94096 468528
rect 94516 468518 94544 493037
rect 94504 468512 94556 468518
rect 94504 468454 94556 468460
rect 94976 467294 95004 493037
rect 95344 491230 95372 493037
rect 95332 491224 95384 491230
rect 95332 491166 95384 491172
rect 95804 471714 95832 493037
rect 96264 483682 96292 493037
rect 96738 493023 96844 493051
rect 96816 487626 96844 493023
rect 97184 490686 97212 493037
rect 97172 490680 97224 490686
rect 97172 490622 97224 490628
rect 97552 487762 97580 493037
rect 98012 488510 98040 493037
rect 98000 488504 98052 488510
rect 98000 488446 98052 488452
rect 97540 487756 97592 487762
rect 97540 487698 97592 487704
rect 98472 487694 98500 493037
rect 98460 487688 98512 487694
rect 98460 487630 98512 487636
rect 96804 487620 96856 487626
rect 96804 487562 96856 487568
rect 96252 483676 96304 483682
rect 96252 483618 96304 483624
rect 98932 474570 98960 493037
rect 99392 492046 99420 493037
rect 99380 492040 99432 492046
rect 99380 491982 99432 491988
rect 99760 474638 99788 493037
rect 100220 490618 100248 493037
rect 100208 490612 100260 490618
rect 100208 490554 100260 490560
rect 99748 474632 99800 474638
rect 99748 474574 99800 474580
rect 98920 474564 98972 474570
rect 98920 474506 98972 474512
rect 100680 474502 100708 493037
rect 100668 474496 100720 474502
rect 100668 474438 100720 474444
rect 95792 471708 95844 471714
rect 95792 471650 95844 471656
rect 101140 471510 101168 493037
rect 101128 471504 101180 471510
rect 101128 471446 101180 471452
rect 101508 471442 101536 493037
rect 101496 471436 101548 471442
rect 101496 471378 101548 471384
rect 94964 467288 95016 467294
rect 94964 467230 95016 467236
rect 93584 465792 93636 465798
rect 93584 465734 93636 465740
rect 93216 464772 93268 464778
rect 93216 464714 93268 464720
rect 101968 464710 101996 493037
rect 102428 471578 102456 493037
rect 102888 471646 102916 493037
rect 103348 491094 103376 493037
rect 103336 491088 103388 491094
rect 103336 491030 103388 491036
rect 103716 474298 103744 493037
rect 103704 474292 103756 474298
rect 103704 474234 103756 474240
rect 102876 471640 102928 471646
rect 102876 471582 102928 471588
rect 102416 471572 102468 471578
rect 102416 471514 102468 471520
rect 104176 471306 104204 493037
rect 104636 491026 104664 493037
rect 104624 491020 104676 491026
rect 104624 490962 104676 490968
rect 105096 474434 105124 493037
rect 105084 474428 105136 474434
rect 105084 474370 105136 474376
rect 105556 474230 105584 493037
rect 105924 474366 105952 493037
rect 105912 474360 105964 474366
rect 105912 474302 105964 474308
rect 105544 474224 105596 474230
rect 105544 474166 105596 474172
rect 106384 474162 106412 493037
rect 106372 474156 106424 474162
rect 106372 474098 106424 474104
rect 106844 474094 106872 493037
rect 106832 474088 106884 474094
rect 106832 474030 106884 474036
rect 104164 471300 104216 471306
rect 104164 471242 104216 471248
rect 107304 467158 107332 493037
rect 107292 467152 107344 467158
rect 107292 467094 107344 467100
rect 107764 465769 107792 493037
rect 108132 468586 108160 493037
rect 108120 468580 108172 468586
rect 108120 468522 108172 468528
rect 108592 468518 108620 493037
rect 109052 492046 109080 493037
rect 109040 492040 109092 492046
rect 109040 491982 109092 491988
rect 109512 471306 109540 493037
rect 109500 471300 109552 471306
rect 109500 471242 109552 471248
rect 109880 468654 109908 493037
rect 110340 490618 110368 493037
rect 110328 490612 110380 490618
rect 110328 490554 110380 490560
rect 110800 484906 110828 493037
rect 111260 488306 111288 493037
rect 111720 488374 111748 493037
rect 111708 488368 111760 488374
rect 111708 488310 111760 488316
rect 111248 488300 111300 488306
rect 111248 488242 111300 488248
rect 112088 488170 112116 493037
rect 112076 488164 112128 488170
rect 112076 488106 112128 488112
rect 110788 484900 110840 484906
rect 110788 484842 110840 484848
rect 109868 468648 109920 468654
rect 109868 468590 109920 468596
rect 108580 468512 108632 468518
rect 108580 468454 108632 468460
rect 112548 467226 112576 493037
rect 113008 469878 113036 493037
rect 112996 469872 113048 469878
rect 112996 469814 113048 469820
rect 113468 468722 113496 493037
rect 113928 472666 113956 493037
rect 114296 483002 114324 493037
rect 114284 482996 114336 483002
rect 114284 482938 114336 482944
rect 113916 472660 113968 472666
rect 113916 472602 113968 472608
rect 114756 471374 114784 493037
rect 115216 488102 115244 493037
rect 115204 488096 115256 488102
rect 115204 488038 115256 488044
rect 115676 488034 115704 493037
rect 116044 488238 116072 493037
rect 116032 488232 116084 488238
rect 116032 488174 116084 488180
rect 115664 488028 115716 488034
rect 115664 487970 115716 487976
rect 116504 485353 116532 493037
rect 116490 485344 116546 485353
rect 116490 485279 116546 485288
rect 116964 485042 116992 493037
rect 117424 485489 117452 493037
rect 117410 485480 117466 485489
rect 117410 485415 117466 485424
rect 116952 485036 117004 485042
rect 116952 484978 117004 484984
rect 117884 484974 117912 493037
rect 118252 485081 118280 493037
rect 118712 485217 118740 493037
rect 119172 485654 119200 493037
rect 119632 488442 119660 493037
rect 119620 488436 119672 488442
rect 119620 488378 119672 488384
rect 120092 488073 120120 493037
rect 120460 488209 120488 493037
rect 120446 488200 120502 488209
rect 120446 488135 120502 488144
rect 120078 488064 120134 488073
rect 120078 487999 120134 488008
rect 120920 487937 120948 493037
rect 121380 488345 121408 493037
rect 121366 488336 121422 488345
rect 121366 488271 121422 488280
rect 120906 487928 120962 487937
rect 120906 487863 120962 487872
rect 119160 485648 119212 485654
rect 119160 485590 119212 485596
rect 118698 485208 118754 485217
rect 118698 485143 118754 485152
rect 118238 485072 118294 485081
rect 118238 485007 118294 485016
rect 117872 484968 117924 484974
rect 117872 484910 117924 484916
rect 114744 471368 114796 471374
rect 114744 471310 114796 471316
rect 113456 468716 113508 468722
rect 113456 468658 113508 468664
rect 112536 467220 112588 467226
rect 112536 467162 112588 467168
rect 107750 465760 107806 465769
rect 107750 465695 107806 465704
rect 101956 464704 102008 464710
rect 101956 464646 102008 464652
rect 121840 464574 121868 493037
rect 122208 474065 122236 493037
rect 122194 474056 122250 474065
rect 122194 473991 122250 474000
rect 122668 464642 122696 493037
rect 123128 482458 123156 493037
rect 123588 482730 123616 493037
rect 123576 482724 123628 482730
rect 123576 482666 123628 482672
rect 123116 482452 123168 482458
rect 123116 482394 123168 482400
rect 124048 482225 124076 493037
rect 124416 482662 124444 493037
rect 124404 482656 124456 482662
rect 124404 482598 124456 482604
rect 124876 482594 124904 493037
rect 124864 482588 124916 482594
rect 124864 482530 124916 482536
rect 125336 482361 125364 493037
rect 125796 482526 125824 493037
rect 126256 482798 126284 493037
rect 126624 487801 126652 493037
rect 126610 487792 126666 487801
rect 126610 487727 126666 487736
rect 126244 482792 126296 482798
rect 126244 482734 126296 482740
rect 125784 482520 125836 482526
rect 125784 482462 125836 482468
rect 125322 482352 125378 482361
rect 125322 482287 125378 482296
rect 124034 482216 124090 482225
rect 124034 482151 124090 482160
rect 127084 471374 127112 493037
rect 127544 474094 127572 493037
rect 128004 482934 128032 493037
rect 127992 482928 128044 482934
rect 127992 482870 128044 482876
rect 128464 482497 128492 493037
rect 128832 482866 128860 493037
rect 129292 485450 129320 493037
rect 129752 485586 129780 493037
rect 129740 485580 129792 485586
rect 129740 485522 129792 485528
rect 129280 485444 129332 485450
rect 129280 485386 129332 485392
rect 130212 485246 130240 493037
rect 130200 485240 130252 485246
rect 130200 485182 130252 485188
rect 130580 485178 130608 493037
rect 131040 485382 131068 493037
rect 131028 485376 131080 485382
rect 131028 485318 131080 485324
rect 131500 485314 131528 493037
rect 131960 487898 131988 493037
rect 131948 487892 132000 487898
rect 131948 487834 132000 487840
rect 132420 485790 132448 493037
rect 132408 485784 132460 485790
rect 132408 485726 132460 485732
rect 132788 485722 132816 493037
rect 133144 487960 133196 487966
rect 133144 487902 133196 487908
rect 132776 485716 132828 485722
rect 132776 485658 132828 485664
rect 131488 485308 131540 485314
rect 131488 485250 131540 485256
rect 130568 485172 130620 485178
rect 130568 485114 130620 485120
rect 128820 482860 128872 482866
rect 128820 482802 128872 482808
rect 128450 482488 128506 482497
rect 128450 482423 128506 482432
rect 127532 474088 127584 474094
rect 127532 474030 127584 474036
rect 127072 471368 127124 471374
rect 127072 471310 127124 471316
rect 133156 467838 133184 487902
rect 133248 485110 133276 493037
rect 133236 485104 133288 485110
rect 133236 485046 133288 485052
rect 133708 482390 133736 493037
rect 133696 482384 133748 482390
rect 133696 482326 133748 482332
rect 133144 467832 133196 467838
rect 133144 467774 133196 467780
rect 122656 464636 122708 464642
rect 122656 464578 122708 464584
rect 121828 464568 121880 464574
rect 121828 464510 121880 464516
rect 134168 464438 134196 493037
rect 134628 487830 134656 493037
rect 134616 487824 134668 487830
rect 134616 487766 134668 487772
rect 134996 464506 135024 493037
rect 135456 487898 135484 493037
rect 135444 487892 135496 487898
rect 135444 487834 135496 487840
rect 135916 485518 135944 493037
rect 136376 488034 136404 493037
rect 136744 488102 136772 493037
rect 136732 488096 136784 488102
rect 136732 488038 136784 488044
rect 136364 488028 136416 488034
rect 136364 487970 136416 487976
rect 135904 485512 135956 485518
rect 135904 485454 135956 485460
rect 134984 464500 135036 464506
rect 134984 464442 135036 464448
rect 137204 464438 137232 493037
rect 137664 488170 137692 493037
rect 137652 488164 137704 488170
rect 137652 488106 137704 488112
rect 138124 487966 138152 493037
rect 138584 488238 138612 493037
rect 138952 490686 138980 493037
rect 139412 490754 139440 493037
rect 139400 490748 139452 490754
rect 139400 490690 139452 490696
rect 138940 490680 138992 490686
rect 138940 490622 138992 490628
rect 138572 488232 138624 488238
rect 138572 488174 138624 488180
rect 138112 487960 138164 487966
rect 138112 487902 138164 487908
rect 139872 474162 139900 493037
rect 139860 474156 139912 474162
rect 139860 474098 139912 474104
rect 140332 471646 140360 493037
rect 140792 492114 140820 493037
rect 140780 492108 140832 492114
rect 140780 492050 140832 492056
rect 140320 471640 140372 471646
rect 140320 471582 140372 471588
rect 141160 471578 141188 493037
rect 141148 471572 141200 471578
rect 141148 471514 141200 471520
rect 141620 471510 141648 493037
rect 141608 471504 141660 471510
rect 141608 471446 141660 471452
rect 142080 471442 142108 493037
rect 142068 471436 142120 471442
rect 142068 471378 142120 471384
rect 142540 465798 142568 493037
rect 142528 465792 142580 465798
rect 142528 465734 142580 465740
rect 142908 464506 142936 493037
rect 143368 465866 143396 493037
rect 143828 482322 143856 493037
rect 144288 486470 144316 493037
rect 144748 487830 144776 493037
rect 145116 490521 145144 493037
rect 145102 490512 145158 490521
rect 145102 490447 145158 490456
rect 144736 487824 144788 487830
rect 144736 487766 144788 487772
rect 144276 486464 144328 486470
rect 144276 486406 144328 486412
rect 143816 482316 143868 482322
rect 143816 482258 143868 482264
rect 145576 479505 145604 493037
rect 145562 479496 145618 479505
rect 145562 479431 145618 479440
rect 146036 474337 146064 493037
rect 146496 490657 146524 493037
rect 146482 490648 146538 490657
rect 146482 490583 146538 490592
rect 146956 482225 146984 493037
rect 146942 482216 146998 482225
rect 146942 482151 146998 482160
rect 146022 474328 146078 474337
rect 146022 474263 146078 474272
rect 147324 468489 147352 493037
rect 147784 490793 147812 493037
rect 147770 490784 147826 490793
rect 147770 490719 147826 490728
rect 148244 475454 148272 493037
rect 148704 476785 148732 493037
rect 149164 489161 149192 493037
rect 149532 491094 149560 493037
rect 149520 491088 149572 491094
rect 149520 491030 149572 491036
rect 149992 490958 150020 493037
rect 149980 490952 150032 490958
rect 149980 490894 150032 490900
rect 149150 489152 149206 489161
rect 149150 489087 149206 489096
rect 150452 481001 150480 493037
rect 150912 491230 150940 493037
rect 150900 491224 150952 491230
rect 150900 491166 150952 491172
rect 151280 483721 151308 493037
rect 151266 483712 151322 483721
rect 151266 483647 151322 483656
rect 150438 480992 150494 481001
rect 150438 480927 150494 480936
rect 148690 476776 148746 476785
rect 148690 476711 148746 476720
rect 148232 475448 148284 475454
rect 148232 475390 148284 475396
rect 151740 474201 151768 493037
rect 152200 491162 152228 493037
rect 152188 491156 152240 491162
rect 152188 491098 152240 491104
rect 152660 485081 152688 493037
rect 153120 490414 153148 493037
rect 153488 491298 153516 493037
rect 153476 491292 153528 491298
rect 153476 491234 153528 491240
rect 153108 490408 153160 490414
rect 153108 490350 153160 490356
rect 152646 485072 152702 485081
rect 152646 485007 152702 485016
rect 153948 475425 153976 493037
rect 154408 490482 154436 493037
rect 154396 490476 154448 490482
rect 154396 490418 154448 490424
rect 153934 475416 153990 475425
rect 153934 475351 153990 475360
rect 151726 474192 151782 474201
rect 151726 474127 151782 474136
rect 154868 468625 154896 493037
rect 155328 490822 155356 493037
rect 155316 490816 155368 490822
rect 155316 490758 155368 490764
rect 155696 482497 155724 493037
rect 155682 482488 155738 482497
rect 155682 482423 155738 482432
rect 156156 482361 156184 493037
rect 156616 490890 156644 493037
rect 156604 490884 156656 490890
rect 156604 490826 156656 490832
rect 156142 482352 156198 482361
rect 156142 482287 156198 482296
rect 157076 476921 157104 493037
rect 157444 490550 157472 493037
rect 157904 491026 157932 493037
rect 157892 491020 157944 491026
rect 157892 490962 157944 490968
rect 157432 490544 157484 490550
rect 157432 490486 157484 490492
rect 158364 478145 158392 493037
rect 158824 483857 158852 493037
rect 158810 483848 158866 483857
rect 158810 483783 158866 483792
rect 159284 478242 159312 493037
rect 159652 485110 159680 493037
rect 160112 488306 160140 493037
rect 160100 488300 160152 488306
rect 160100 488242 160152 488248
rect 159640 485104 159692 485110
rect 159640 485046 159692 485052
rect 159272 478236 159324 478242
rect 159272 478178 159324 478184
rect 158350 478136 158406 478145
rect 158350 478071 158406 478080
rect 157062 476912 157118 476921
rect 157062 476847 157118 476856
rect 160572 471345 160600 493037
rect 160744 489184 160796 489190
rect 160744 489126 160796 489132
rect 160558 471336 160614 471345
rect 160558 471271 160614 471280
rect 154854 468616 154910 468625
rect 154854 468551 154910 468560
rect 147310 468480 147366 468489
rect 147310 468415 147366 468424
rect 160756 467770 160784 489126
rect 161032 472666 161060 493037
rect 161020 472660 161072 472666
rect 161020 472602 161072 472608
rect 161492 469878 161520 493037
rect 161480 469872 161532 469878
rect 161480 469814 161532 469820
rect 161860 468897 161888 493037
rect 162320 480962 162348 493037
rect 162308 480956 162360 480962
rect 162308 480898 162360 480904
rect 162780 471481 162808 493037
rect 163240 476882 163268 493037
rect 163228 476876 163280 476882
rect 163228 476818 163280 476824
rect 162766 471472 162822 471481
rect 162766 471407 162822 471416
rect 163608 471209 163636 493037
rect 164068 489190 164096 493037
rect 164056 489184 164108 489190
rect 164056 489126 164108 489132
rect 164528 486538 164556 493037
rect 164516 486532 164568 486538
rect 164516 486474 164568 486480
rect 163594 471200 163650 471209
rect 163594 471135 163650 471144
rect 161846 468888 161902 468897
rect 161846 468823 161902 468832
rect 160744 467764 160796 467770
rect 160744 467706 160796 467712
rect 164988 465934 165016 493037
rect 165448 467158 165476 493037
rect 165816 474473 165844 493037
rect 166276 479602 166304 493037
rect 166264 479596 166316 479602
rect 166264 479538 166316 479544
rect 165802 474464 165858 474473
rect 165802 474399 165858 474408
rect 165436 467152 165488 467158
rect 165436 467094 165488 467100
rect 166736 466070 166764 493037
rect 166724 466064 166776 466070
rect 167196 466041 167224 493037
rect 167656 489258 167684 493037
rect 167644 489252 167696 489258
rect 167644 489194 167696 489200
rect 168024 466206 168052 493037
rect 168484 468858 168512 493037
rect 168472 468852 168524 468858
rect 168472 468794 168524 468800
rect 168012 466200 168064 466206
rect 168012 466142 168064 466148
rect 166724 466006 166776 466012
rect 167182 466032 167238 466041
rect 167182 465967 167238 465976
rect 164976 465928 165028 465934
rect 168944 465905 168972 493037
rect 169404 468790 169432 493037
rect 169392 468784 169444 468790
rect 169864 468761 169892 493037
rect 169392 468726 169444 468732
rect 169850 468752 169906 468761
rect 170232 468722 170260 493037
rect 170692 475522 170720 493037
rect 170680 475516 170732 475522
rect 170680 475458 170732 475464
rect 169850 468687 169906 468696
rect 170220 468716 170272 468722
rect 170220 468658 170272 468664
rect 171152 467129 171180 493037
rect 171612 467226 171640 493037
rect 171980 482322 172008 493037
rect 171968 482316 172020 482322
rect 171968 482258 172020 482264
rect 172440 471753 172468 493037
rect 172900 472569 172928 493037
rect 172886 472560 172942 472569
rect 172886 472495 172942 472504
rect 173360 471889 173388 493037
rect 173346 471880 173402 471889
rect 173346 471815 173402 471824
rect 172426 471744 172482 471753
rect 172426 471679 172482 471688
rect 173820 470014 173848 493037
rect 173808 470008 173860 470014
rect 173808 469950 173860 469956
rect 171600 467220 171652 467226
rect 171600 467162 171652 467168
rect 171138 467120 171194 467129
rect 171138 467055 171194 467064
rect 174188 466274 174216 493037
rect 174176 466268 174228 466274
rect 174176 466210 174228 466216
rect 174648 466002 174676 493037
rect 175108 471782 175136 493037
rect 175096 471776 175148 471782
rect 175096 471718 175148 471724
rect 175568 470082 175596 493037
rect 176028 472802 176056 493037
rect 176396 479670 176424 493037
rect 176384 479664 176436 479670
rect 176384 479606 176436 479612
rect 176016 472796 176068 472802
rect 176016 472738 176068 472744
rect 176856 472734 176884 493037
rect 177316 486606 177344 493037
rect 177304 486600 177356 486606
rect 177304 486542 177356 486548
rect 177776 481030 177804 493037
rect 177764 481024 177816 481030
rect 177764 480966 177816 480972
rect 176844 472728 176896 472734
rect 176844 472670 176896 472676
rect 175556 470076 175608 470082
rect 175556 470018 175608 470024
rect 178144 469946 178172 493037
rect 178604 476950 178632 493037
rect 178592 476944 178644 476950
rect 178592 476886 178644 476892
rect 179064 471714 179092 493037
rect 179052 471708 179104 471714
rect 179052 471650 179104 471656
rect 178132 469940 178184 469946
rect 178132 469882 178184 469888
rect 178040 467832 178092 467838
rect 178040 467774 178092 467780
rect 178052 466614 178080 467774
rect 179420 467764 179472 467770
rect 179420 467706 179472 467712
rect 178040 466608 178092 466614
rect 178038 466576 178040 466585
rect 179432 466585 179460 467706
rect 178092 466576 178094 466585
rect 178038 466511 178094 466520
rect 179418 466576 179474 466585
rect 179418 466511 179420 466520
rect 179472 466511 179474 466520
rect 179420 466482 179472 466488
rect 179432 466451 179460 466482
rect 179524 466138 179552 493037
rect 179984 490929 180012 493037
rect 179970 490920 180026 490929
rect 179970 490855 180026 490864
rect 180064 490612 180116 490618
rect 180064 490554 180116 490560
rect 180076 466177 180104 490554
rect 180352 466342 180380 493037
rect 180340 466336 180392 466342
rect 180340 466278 180392 466284
rect 180062 466168 180118 466177
rect 179512 466132 179564 466138
rect 180062 466103 180118 466112
rect 179512 466074 179564 466080
rect 174636 465996 174688 466002
rect 174636 465938 174688 465944
rect 164976 465870 165028 465876
rect 168930 465896 168986 465905
rect 143356 465860 143408 465866
rect 168930 465831 168986 465840
rect 143356 465802 143408 465808
rect 180812 464574 180840 493037
rect 181272 469033 181300 493037
rect 181732 469130 181760 493037
rect 181720 469124 181772 469130
rect 181720 469066 181772 469072
rect 181258 469024 181314 469033
rect 181258 468959 181314 468968
rect 182192 467362 182220 493037
rect 182560 471617 182588 493037
rect 183020 471850 183048 493037
rect 183008 471844 183060 471850
rect 183008 471786 183060 471792
rect 182546 471608 182602 471617
rect 182546 471543 182602 471552
rect 182180 467356 182232 467362
rect 182180 467298 182232 467304
rect 180800 464568 180852 464574
rect 180800 464510 180852 464516
rect 142896 464500 142948 464506
rect 142896 464442 142948 464448
rect 134156 464432 134208 464438
rect 92294 464400 92350 464409
rect 134156 464374 134208 464380
rect 137192 464432 137244 464438
rect 183480 464409 183508 493037
rect 183940 468382 183968 493037
rect 184308 483682 184336 493037
rect 184768 491065 184796 493037
rect 184754 491056 184810 491065
rect 184754 490991 184810 491000
rect 184296 483676 184348 483682
rect 184296 483618 184348 483624
rect 183928 468376 183980 468382
rect 183928 468318 183980 468324
rect 185228 467430 185256 493037
rect 185688 491201 185716 493037
rect 185674 491192 185730 491201
rect 185674 491127 185730 491136
rect 186148 474230 186176 493037
rect 186136 474224 186188 474230
rect 186136 474166 186188 474172
rect 186516 469198 186544 493037
rect 186976 490385 187004 493037
rect 186962 490376 187018 490385
rect 186962 490311 187018 490320
rect 187436 472870 187464 493037
rect 187424 472864 187476 472870
rect 187424 472806 187476 472812
rect 186504 469192 186556 469198
rect 186504 469134 186556 469140
rect 185216 467424 185268 467430
rect 185216 467366 185268 467372
rect 187896 465662 187924 493037
rect 188356 467294 188384 493037
rect 188724 471170 188752 493037
rect 188712 471164 188764 471170
rect 188712 471106 188764 471112
rect 188344 467288 188396 467294
rect 188344 467230 188396 467236
rect 187884 465656 187936 465662
rect 187884 465598 187936 465604
rect 189184 465594 189212 493037
rect 189644 468926 189672 493037
rect 189632 468920 189684 468926
rect 189632 468862 189684 468868
rect 190104 467498 190132 493037
rect 190472 468994 190500 493037
rect 190932 471918 190960 493037
rect 190920 471912 190972 471918
rect 190920 471854 190972 471860
rect 191392 471238 191420 493037
rect 191380 471232 191432 471238
rect 191380 471174 191432 471180
rect 190460 468988 190512 468994
rect 190460 468930 190512 468936
rect 190092 467492 190144 467498
rect 190092 467434 190144 467440
rect 190918 466576 190974 466585
rect 190918 466511 190974 466520
rect 190932 466478 190960 466511
rect 190920 466472 190972 466478
rect 190920 466414 190972 466420
rect 189172 465588 189224 465594
rect 189172 465530 189224 465536
rect 191852 464710 191880 493037
rect 192312 464778 192340 493037
rect 192680 469062 192708 493037
rect 193140 471986 193168 493037
rect 193128 471980 193180 471986
rect 193128 471922 193180 471928
rect 192668 469056 192720 469062
rect 192668 468998 192720 469004
rect 193600 468450 193628 493037
rect 193956 490748 194008 490754
rect 193956 490690 194008 490696
rect 193864 490680 193916 490686
rect 193864 490622 193916 490628
rect 193876 470626 193904 490622
rect 193968 474298 193996 490690
rect 193956 474292 194008 474298
rect 193956 474234 194008 474240
rect 193864 470620 193916 470626
rect 193864 470562 193916 470568
rect 193588 468444 193640 468450
rect 193588 468386 193640 468392
rect 194060 466410 194088 493037
rect 194048 466404 194100 466410
rect 194048 466346 194100 466352
rect 192300 464772 192352 464778
rect 192300 464714 192352 464720
rect 191840 464704 191892 464710
rect 191840 464646 191892 464652
rect 194520 464642 194548 493037
rect 194888 490754 194916 493037
rect 194876 490748 194928 490754
rect 194876 490690 194928 490696
rect 195348 490686 195376 493037
rect 195336 490680 195388 490686
rect 195336 490622 195388 490628
rect 195808 465526 195836 493037
rect 195796 465520 195848 465526
rect 195796 465462 195848 465468
rect 194508 464636 194560 464642
rect 194508 464578 194560 464584
rect 137192 464374 137244 464380
rect 183466 464400 183522 464409
rect 92294 464335 92350 464344
rect 183466 464335 183522 464344
rect 195060 380996 195112 381002
rect 195060 380938 195112 380944
rect 60740 380928 60792 380934
rect 60740 380870 60792 380876
rect 194600 380928 194652 380934
rect 194600 380870 194652 380876
rect 60752 357406 60780 380870
rect 155960 380588 156012 380594
rect 155960 380530 156012 380536
rect 143632 380520 143684 380526
rect 143632 380462 143684 380468
rect 118332 380452 118384 380458
rect 118332 380394 118384 380400
rect 121000 380452 121052 380458
rect 121000 380394 121052 380400
rect 113548 380384 113600 380390
rect 110970 380352 111026 380361
rect 110970 380287 110972 380296
rect 111024 380287 111026 380296
rect 113546 380352 113548 380361
rect 118344 380361 118372 380394
rect 121012 380361 121040 380394
rect 143644 380361 143672 380462
rect 155972 380361 156000 380530
rect 163504 380384 163556 380390
rect 113600 380352 113602 380361
rect 113546 380287 113602 380296
rect 115938 380352 115994 380361
rect 115938 380287 115994 380296
rect 118330 380352 118386 380361
rect 118330 380287 118386 380296
rect 120998 380352 121054 380361
rect 120998 380287 121054 380296
rect 123482 380352 123538 380361
rect 123482 380287 123538 380296
rect 128358 380352 128414 380361
rect 128358 380287 128414 380296
rect 135902 380352 135958 380361
rect 135902 380287 135958 380296
rect 143630 380352 143686 380361
rect 143630 380287 143686 380296
rect 148598 380352 148654 380361
rect 148598 380287 148600 380296
rect 110972 380258 111024 380264
rect 99378 380216 99434 380225
rect 115952 380186 115980 380287
rect 123496 380254 123524 380287
rect 123484 380248 123536 380254
rect 123484 380190 123536 380196
rect 128372 380186 128400 380287
rect 135916 380254 135944 380287
rect 148652 380287 148654 380296
rect 155958 380352 156014 380361
rect 155958 380287 156014 380296
rect 158534 380352 158590 380361
rect 158534 380287 158590 380296
rect 160926 380352 160982 380361
rect 160926 380287 160982 380296
rect 163502 380352 163504 380361
rect 163556 380352 163558 380361
rect 163502 380287 163558 380296
rect 166078 380352 166134 380361
rect 166078 380287 166134 380296
rect 148600 380258 148652 380264
rect 135904 380248 135956 380254
rect 135904 380190 135956 380196
rect 99378 380151 99434 380160
rect 115940 380180 115992 380186
rect 88340 379500 88392 379506
rect 88340 379442 88392 379448
rect 92388 379500 92440 379506
rect 92388 379442 92440 379448
rect 86592 379432 86644 379438
rect 77206 379400 77262 379409
rect 77206 379335 77262 379344
rect 80426 379400 80482 379409
rect 80426 379335 80482 379344
rect 85486 379400 85542 379409
rect 85486 379335 85488 379344
rect 76838 379264 76894 379273
rect 76838 379199 76894 379208
rect 76852 378865 76880 379199
rect 76838 378856 76894 378865
rect 76838 378791 76894 378800
rect 77220 378758 77248 379335
rect 77208 378752 77260 378758
rect 80440 378729 80468 379335
rect 85540 379335 85542 379344
rect 86590 379400 86592 379409
rect 88352 379409 88380 379442
rect 92400 379409 92428 379442
rect 86644 379400 86646 379409
rect 86590 379335 86646 379344
rect 88338 379400 88394 379409
rect 88338 379335 88394 379344
rect 88798 379400 88854 379409
rect 88798 379335 88854 379344
rect 90730 379400 90786 379409
rect 90730 379335 90786 379344
rect 91374 379400 91430 379409
rect 91374 379335 91430 379344
rect 92386 379400 92442 379409
rect 92386 379335 92442 379344
rect 93582 379400 93638 379409
rect 93582 379335 93638 379344
rect 96066 379400 96122 379409
rect 96066 379335 96122 379344
rect 98458 379400 98514 379409
rect 98458 379335 98514 379344
rect 85488 379306 85540 379312
rect 88812 379302 88840 379335
rect 88800 379296 88852 379302
rect 88800 379238 88852 379244
rect 90744 379166 90772 379335
rect 90822 379264 90878 379273
rect 91388 379234 91416 379335
rect 93490 379264 93546 379273
rect 90822 379199 90878 379208
rect 91376 379228 91428 379234
rect 90836 379166 90864 379199
rect 93490 379199 93546 379208
rect 91376 379170 91428 379176
rect 90732 379160 90784 379166
rect 90732 379102 90784 379108
rect 90824 379160 90876 379166
rect 90824 379102 90876 379108
rect 93504 379098 93532 379199
rect 93596 379098 93624 379335
rect 93492 379092 93544 379098
rect 93492 379034 93544 379040
rect 93584 379092 93636 379098
rect 93584 379034 93636 379040
rect 77208 378694 77260 378700
rect 80426 378720 80482 378729
rect 80426 378655 80482 378664
rect 77114 378584 77170 378593
rect 77114 378519 77170 378528
rect 77128 376106 77156 378519
rect 80440 378214 80468 378655
rect 96080 378622 96108 379335
rect 98472 378690 98500 379335
rect 99392 378758 99420 380151
rect 115940 380122 115992 380128
rect 128360 380180 128412 380186
rect 128360 380122 128412 380128
rect 158548 380118 158576 380287
rect 158536 380112 158588 380118
rect 158536 380054 158588 380060
rect 160940 380050 160968 380287
rect 160928 380044 160980 380050
rect 160928 379986 160980 379992
rect 166092 379982 166120 380287
rect 166080 379976 166132 379982
rect 166080 379918 166132 379924
rect 101034 379400 101090 379409
rect 101034 379335 101090 379344
rect 103518 379400 103574 379409
rect 103518 379335 103574 379344
rect 105358 379400 105414 379409
rect 105358 379335 105414 379344
rect 108210 379400 108266 379409
rect 108210 379335 108266 379344
rect 108854 379400 108910 379409
rect 108854 379335 108910 379344
rect 109774 379400 109830 379409
rect 109774 379335 109830 379344
rect 111246 379400 111302 379409
rect 111246 379335 111302 379344
rect 112350 379400 112406 379409
rect 112350 379335 112406 379344
rect 113454 379400 113510 379409
rect 113454 379335 113510 379344
rect 114466 379400 114522 379409
rect 114466 379335 114522 379344
rect 115846 379400 115902 379409
rect 115846 379335 115902 379344
rect 117134 379400 117190 379409
rect 117134 379335 117190 379344
rect 141054 379400 141110 379409
rect 141054 379335 141110 379344
rect 146022 379400 146078 379409
rect 146022 379335 146078 379344
rect 150990 379400 151046 379409
rect 150990 379335 151046 379344
rect 153566 379400 153622 379409
rect 153566 379335 153622 379344
rect 99470 379264 99526 379273
rect 99470 379199 99526 379208
rect 99380 378752 99432 378758
rect 99380 378694 99432 378700
rect 98460 378684 98512 378690
rect 98460 378626 98512 378632
rect 96068 378616 96120 378622
rect 96068 378558 96120 378564
rect 97078 378584 97134 378593
rect 97078 378519 97134 378528
rect 98550 378584 98606 378593
rect 98550 378519 98606 378528
rect 80428 378208 80480 378214
rect 80428 378150 80480 378156
rect 97092 376514 97120 378519
rect 97080 376508 97132 376514
rect 97080 376450 97132 376456
rect 77116 376100 77168 376106
rect 77116 376042 77168 376048
rect 98564 376038 98592 378519
rect 99484 376650 99512 379199
rect 101048 378826 101076 379335
rect 102966 379264 103022 379273
rect 102966 379199 103022 379208
rect 101036 378820 101088 378826
rect 101036 378762 101088 378768
rect 101862 378584 101918 378593
rect 101862 378519 101918 378528
rect 100758 378312 100814 378321
rect 100758 378247 100814 378256
rect 99472 376644 99524 376650
rect 99472 376586 99524 376592
rect 98552 376032 98604 376038
rect 98552 375974 98604 375980
rect 100772 375358 100800 378247
rect 101876 376582 101904 378519
rect 101864 376576 101916 376582
rect 101864 376518 101916 376524
rect 100760 375352 100812 375358
rect 100760 375294 100812 375300
rect 102980 374746 103008 379199
rect 103532 378894 103560 379335
rect 104254 379264 104310 379273
rect 104254 379199 104310 379208
rect 103520 378888 103572 378894
rect 103520 378830 103572 378836
rect 104268 377262 104296 379199
rect 105372 378962 105400 379335
rect 108224 379030 108252 379335
rect 108212 379024 108264 379030
rect 108212 378966 108264 378972
rect 105360 378956 105412 378962
rect 105360 378898 105412 378904
rect 107566 378584 107622 378593
rect 107566 378519 107622 378528
rect 104256 377256 104308 377262
rect 104256 377198 104308 377204
rect 107580 376446 107608 378519
rect 108868 377777 108896 379335
rect 109788 378214 109816 379335
rect 111260 378350 111288 379335
rect 112364 378962 112392 379335
rect 112352 378956 112404 378962
rect 112352 378898 112404 378904
rect 113468 378554 113496 379335
rect 113456 378548 113508 378554
rect 113456 378490 113508 378496
rect 114480 378418 114508 379335
rect 115860 379030 115888 379335
rect 115848 379024 115900 379030
rect 115848 378966 115900 378972
rect 117148 378894 117176 379335
rect 117136 378888 117188 378894
rect 117136 378830 117188 378836
rect 125966 378448 126022 378457
rect 114468 378412 114520 378418
rect 125966 378383 126022 378392
rect 131026 378448 131082 378457
rect 131026 378383 131082 378392
rect 133510 378448 133566 378457
rect 133510 378383 133566 378392
rect 138478 378448 138534 378457
rect 138478 378383 138534 378392
rect 114468 378354 114520 378360
rect 111248 378344 111300 378350
rect 111248 378286 111300 378292
rect 109776 378208 109828 378214
rect 109776 378150 109828 378156
rect 108854 377768 108910 377777
rect 108854 377703 108910 377712
rect 107568 376440 107620 376446
rect 107568 376382 107620 376388
rect 125980 376378 126008 378383
rect 125968 376372 126020 376378
rect 125968 376314 126020 376320
rect 131040 376310 131068 378383
rect 131028 376304 131080 376310
rect 131028 376246 131080 376252
rect 133524 376242 133552 378383
rect 133512 376236 133564 376242
rect 133512 376178 133564 376184
rect 138492 376174 138520 378383
rect 141068 377194 141096 379335
rect 146036 377330 146064 379335
rect 151004 377806 151032 379335
rect 150992 377800 151044 377806
rect 150992 377742 151044 377748
rect 146024 377324 146076 377330
rect 146024 377266 146076 377272
rect 141056 377188 141108 377194
rect 141056 377130 141108 377136
rect 153580 377126 153608 379335
rect 182362 378448 182418 378457
rect 182362 378383 182418 378392
rect 182270 378312 182326 378321
rect 182270 378247 182326 378256
rect 182284 377942 182312 378247
rect 182376 378010 182404 378383
rect 182822 378312 182878 378321
rect 182822 378247 182878 378256
rect 182364 378004 182416 378010
rect 182364 377946 182416 377952
rect 182272 377936 182324 377942
rect 182272 377878 182324 377884
rect 153568 377120 153620 377126
rect 153568 377062 153620 377068
rect 138480 376168 138532 376174
rect 138480 376110 138532 376116
rect 102968 374740 103020 374746
rect 102968 374682 103020 374688
rect 179696 358896 179748 358902
rect 178590 358864 178646 358873
rect 178590 358799 178592 358808
rect 178644 358799 178646 358808
rect 179694 358864 179696 358873
rect 179748 358864 179750 358873
rect 179694 358799 179750 358808
rect 178592 358770 178644 358776
rect 182836 358086 182864 378247
rect 182916 378004 182968 378010
rect 182916 377946 182968 377952
rect 182928 367810 182956 377946
rect 194612 376242 194640 380870
rect 194600 376236 194652 376242
rect 194600 376178 194652 376184
rect 195072 376174 195100 380938
rect 195980 379160 196032 379166
rect 195980 379102 196032 379108
rect 195992 378826 196020 379102
rect 195980 378820 196032 378826
rect 195980 378762 196032 378768
rect 196636 377874 196664 493054
rect 196624 377868 196676 377874
rect 196624 377810 196676 377816
rect 196728 377534 196756 493037
rect 196808 490748 196860 490754
rect 196808 490690 196860 490696
rect 196716 377528 196768 377534
rect 196716 377470 196768 377476
rect 196820 377398 196848 490690
rect 196992 488232 197044 488238
rect 196992 488174 197044 488180
rect 196900 471640 196952 471646
rect 196900 471582 196952 471588
rect 196912 380322 196940 471582
rect 197004 465050 197032 488174
rect 196992 465044 197044 465050
rect 196992 464986 197044 464992
rect 196900 380316 196952 380322
rect 196900 380258 196952 380264
rect 197096 377602 197124 493037
rect 197452 492040 197504 492046
rect 197452 491982 197504 491988
rect 197360 490408 197412 490414
rect 197360 490350 197412 490356
rect 197372 490249 197400 490350
rect 197358 490240 197414 490249
rect 197358 490175 197414 490184
rect 197464 470594 197492 491982
rect 197372 470566 197492 470594
rect 197268 468308 197320 468314
rect 197268 468250 197320 468256
rect 197280 378826 197308 468250
rect 197268 378820 197320 378826
rect 197268 378762 197320 378768
rect 197084 377596 197136 377602
rect 197084 377538 197136 377544
rect 196808 377392 196860 377398
rect 196808 377334 196860 377340
rect 195060 376168 195112 376174
rect 195060 376110 195112 376116
rect 182916 367804 182968 367810
rect 182916 367746 182968 367752
rect 190920 359508 190972 359514
rect 190920 359450 190972 359456
rect 190932 358873 190960 359450
rect 190918 358864 190974 358873
rect 190918 358799 190974 358808
rect 182824 358080 182876 358086
rect 182824 358022 182876 358028
rect 60740 357400 60792 357406
rect 60740 357342 60792 357348
rect 95974 273864 96030 273873
rect 95974 273799 96030 273808
rect 77114 273184 77170 273193
rect 77114 273119 77170 273128
rect 88338 273184 88394 273193
rect 88338 273119 88394 273128
rect 90730 273184 90786 273193
rect 90730 273119 90786 273128
rect 93674 273184 93730 273193
rect 93674 273119 93730 273128
rect 60922 272504 60978 272513
rect 60832 272468 60884 272474
rect 60922 272439 60978 272448
rect 60832 272410 60884 272416
rect 60844 272066 60872 272410
rect 60832 272060 60884 272066
rect 60832 272002 60884 272008
rect 60740 270360 60792 270366
rect 60740 270302 60792 270308
rect 60752 268666 60780 270302
rect 60740 268660 60792 268666
rect 60740 268602 60792 268608
rect 60740 268252 60792 268258
rect 60740 268194 60792 268200
rect 60752 252521 60780 268194
rect 60738 252512 60794 252521
rect 60738 252447 60794 252456
rect 60844 252074 60872 272002
rect 60936 268258 60964 272439
rect 77128 272406 77156 273119
rect 88352 272882 88380 273119
rect 88340 272876 88392 272882
rect 88340 272818 88392 272824
rect 90744 272746 90772 273119
rect 90732 272740 90784 272746
rect 90732 272682 90784 272688
rect 93688 272678 93716 273119
rect 95698 272776 95754 272785
rect 95698 272711 95754 272720
rect 95882 272776 95938 272785
rect 95882 272711 95938 272720
rect 93676 272672 93728 272678
rect 93676 272614 93728 272620
rect 77116 272400 77168 272406
rect 95712 272377 95740 272711
rect 95896 272542 95924 272711
rect 95884 272536 95936 272542
rect 95884 272478 95936 272484
rect 77116 272342 77168 272348
rect 83002 272368 83058 272377
rect 83002 272303 83004 272312
rect 83056 272303 83058 272312
rect 95698 272368 95754 272377
rect 95698 272303 95754 272312
rect 83004 272274 83056 272280
rect 95988 272270 96016 273799
rect 131026 273728 131082 273737
rect 131026 273663 131082 273672
rect 145930 273728 145986 273737
rect 145930 273663 145932 273672
rect 131040 273630 131068 273663
rect 145984 273663 145986 273672
rect 145932 273634 145984 273640
rect 131028 273624 131080 273630
rect 131028 273566 131080 273572
rect 133418 273592 133474 273601
rect 133418 273527 133420 273536
rect 133472 273527 133474 273536
rect 135902 273592 135958 273601
rect 135902 273527 135958 273536
rect 138478 273592 138534 273601
rect 138478 273527 138534 273536
rect 140870 273592 140926 273601
rect 140870 273527 140926 273536
rect 133420 273498 133472 273504
rect 135916 273494 135944 273527
rect 135904 273488 135956 273494
rect 135904 273430 135956 273436
rect 138492 273426 138520 273527
rect 138480 273420 138532 273426
rect 138480 273362 138532 273368
rect 140884 273358 140912 273527
rect 140872 273352 140924 273358
rect 140872 273294 140924 273300
rect 98090 273184 98146 273193
rect 98090 273119 98146 273128
rect 98104 272950 98132 273119
rect 98092 272944 98144 272950
rect 98092 272886 98144 272892
rect 98458 272912 98514 272921
rect 98458 272847 98514 272856
rect 99378 272912 99434 272921
rect 99378 272847 99434 272856
rect 98472 272610 98500 272847
rect 99392 272814 99420 272847
rect 99380 272808 99432 272814
rect 99380 272750 99432 272756
rect 98460 272604 98512 272610
rect 98460 272546 98512 272552
rect 67548 272264 67600 272270
rect 95976 272264 96028 272270
rect 67548 272206 67600 272212
rect 85394 272232 85450 272241
rect 67560 271561 67588 272206
rect 95976 272206 96028 272212
rect 113546 272232 113602 272241
rect 85394 272167 85396 272176
rect 85448 272167 85450 272176
rect 113546 272167 113602 272176
rect 85396 272138 85448 272144
rect 75920 272128 75972 272134
rect 75920 272070 75972 272076
rect 75932 271833 75960 272070
rect 94228 272060 94280 272066
rect 94228 272002 94280 272008
rect 88340 271992 88392 271998
rect 88340 271934 88392 271940
rect 88352 271833 88380 271934
rect 94240 271833 94268 272002
rect 102140 271924 102192 271930
rect 102140 271866 102192 271872
rect 102152 271833 102180 271866
rect 75918 271824 75974 271833
rect 75918 271759 75974 271768
rect 84198 271824 84254 271833
rect 84198 271759 84254 271768
rect 88338 271824 88394 271833
rect 88338 271759 88394 271768
rect 94226 271824 94282 271833
rect 94226 271759 94282 271768
rect 102138 271824 102194 271833
rect 102138 271759 102194 271768
rect 107658 271824 107714 271833
rect 107658 271759 107714 271768
rect 67546 271552 67602 271561
rect 67546 271487 67602 271496
rect 77298 271416 77354 271425
rect 77298 271351 77354 271360
rect 77312 271046 77340 271351
rect 77300 271040 77352 271046
rect 77300 270982 77352 270988
rect 78678 271008 78734 271017
rect 78678 270943 78680 270952
rect 78732 270943 78734 270952
rect 78680 270914 78732 270920
rect 79048 270292 79100 270298
rect 79048 270234 79100 270240
rect 62120 269748 62172 269754
rect 62120 269690 62172 269696
rect 62132 268598 62160 269690
rect 62120 268592 62172 268598
rect 62120 268534 62172 268540
rect 79060 268530 79088 270234
rect 84212 270026 84240 271759
rect 107672 271726 107700 271759
rect 107660 271720 107712 271726
rect 103518 271688 103574 271697
rect 107660 271662 107712 271668
rect 110418 271688 110474 271697
rect 103518 271623 103574 271632
rect 110418 271623 110474 271632
rect 100758 271552 100814 271561
rect 100758 271487 100814 271496
rect 91190 271416 91246 271425
rect 91190 271351 91246 271360
rect 85578 270736 85634 270745
rect 85578 270671 85634 270680
rect 89718 270736 89774 270745
rect 89718 270671 89774 270680
rect 84200 270020 84252 270026
rect 84200 269962 84252 269968
rect 85592 269958 85620 270671
rect 86958 270600 87014 270609
rect 86958 270535 87014 270544
rect 86972 270162 87000 270535
rect 89732 270230 89760 270671
rect 91098 270600 91154 270609
rect 91098 270535 91154 270544
rect 91112 270366 91140 270535
rect 91100 270360 91152 270366
rect 91100 270302 91152 270308
rect 89720 270224 89772 270230
rect 89720 270166 89772 270172
rect 86960 270156 87012 270162
rect 86960 270098 87012 270104
rect 85580 269952 85632 269958
rect 85580 269894 85632 269900
rect 88248 269952 88300 269958
rect 88248 269894 88300 269900
rect 81440 269680 81492 269686
rect 81440 269622 81492 269628
rect 79048 268524 79100 268530
rect 79048 268466 79100 268472
rect 81452 268462 81480 269622
rect 83464 269612 83516 269618
rect 83464 269554 83516 269560
rect 81440 268456 81492 268462
rect 81440 268398 81492 268404
rect 60924 268252 60976 268258
rect 60924 268194 60976 268200
rect 60832 252068 60884 252074
rect 60832 252010 60884 252016
rect 83476 252006 83504 269554
rect 88260 268394 88288 269894
rect 91204 269754 91232 271351
rect 100772 271114 100800 271487
rect 103532 271182 103560 271623
rect 104898 271416 104954 271425
rect 104898 271351 104954 271360
rect 104912 271250 104940 271351
rect 110432 271318 110460 271623
rect 113560 271386 113588 272167
rect 143540 271856 143592 271862
rect 125598 271824 125654 271833
rect 125598 271759 125600 271768
rect 125652 271759 125654 271768
rect 143538 271824 143540 271833
rect 154488 271856 154540 271862
rect 143592 271824 143594 271833
rect 143538 271759 143594 271768
rect 154486 271824 154488 271833
rect 154540 271824 154542 271833
rect 154486 271759 154542 271768
rect 157246 271824 157302 271833
rect 157246 271759 157248 271768
rect 125600 271730 125652 271736
rect 157300 271759 157302 271768
rect 158626 271824 158682 271833
rect 158626 271759 158682 271768
rect 157248 271730 157300 271736
rect 158640 271726 158668 271759
rect 197372 271726 197400 470566
rect 197452 468648 197504 468654
rect 197452 468590 197504 468596
rect 158628 271720 158680 271726
rect 120078 271688 120134 271697
rect 120078 271623 120080 271632
rect 120132 271623 120134 271632
rect 123114 271688 123170 271697
rect 197360 271720 197412 271726
rect 158628 271662 158680 271668
rect 161386 271688 161442 271697
rect 123114 271623 123170 271632
rect 161386 271623 161442 271632
rect 164146 271688 164202 271697
rect 197360 271662 197412 271668
rect 164146 271623 164202 271632
rect 120080 271594 120132 271600
rect 123128 271590 123156 271623
rect 123116 271584 123168 271590
rect 115938 271552 115994 271561
rect 115938 271487 115994 271496
rect 117318 271552 117374 271561
rect 123116 271526 123168 271532
rect 161400 271522 161428 271623
rect 164160 271590 164188 271623
rect 197464 271590 197492 468590
rect 197556 377670 197584 493037
rect 197728 488164 197780 488170
rect 197728 488106 197780 488112
rect 197636 488096 197688 488102
rect 197636 488038 197688 488044
rect 197648 380186 197676 488038
rect 197740 380934 197768 488106
rect 197820 464500 197872 464506
rect 197820 464442 197872 464448
rect 197728 380928 197780 380934
rect 197728 380870 197780 380876
rect 197832 380390 197860 464442
rect 197820 380384 197872 380390
rect 197820 380326 197872 380332
rect 197636 380180 197688 380186
rect 197636 380122 197688 380128
rect 198016 377738 198044 493037
rect 198096 488028 198148 488034
rect 198096 487970 198148 487976
rect 198108 410582 198136 487970
rect 198188 487892 198240 487898
rect 198188 487834 198240 487840
rect 198200 416090 198228 487834
rect 198188 416084 198240 416090
rect 198188 416026 198240 416032
rect 198096 410576 198148 410582
rect 198096 410518 198148 410524
rect 198096 397452 198148 397458
rect 198096 397394 198148 397400
rect 198108 377806 198136 397394
rect 198476 377806 198504 493037
rect 198740 465724 198792 465730
rect 198740 465666 198792 465672
rect 198752 465118 198780 465666
rect 198740 465112 198792 465118
rect 198740 465054 198792 465060
rect 198752 460193 198780 465054
rect 198738 460184 198794 460193
rect 198738 460119 198794 460128
rect 198646 396672 198702 396681
rect 198646 396607 198702 396616
rect 198554 381032 198610 381041
rect 198554 380967 198610 380976
rect 198096 377800 198148 377806
rect 198096 377742 198148 377748
rect 198464 377800 198516 377806
rect 198464 377742 198516 377748
rect 198004 377732 198056 377738
rect 198004 377674 198056 377680
rect 197544 377664 197596 377670
rect 197544 377606 197596 377612
rect 197544 360188 197596 360194
rect 197544 360130 197596 360136
rect 197556 358902 197584 360130
rect 197728 359576 197780 359582
rect 197728 359518 197780 359524
rect 197544 358896 197596 358902
rect 197544 358838 197596 358844
rect 164148 271584 164200 271590
rect 164148 271526 164200 271532
rect 197452 271584 197504 271590
rect 197452 271526 197504 271532
rect 117318 271487 117320 271496
rect 115952 271454 115980 271487
rect 117372 271487 117374 271496
rect 161388 271516 161440 271522
rect 117320 271458 117372 271464
rect 161388 271458 161440 271464
rect 115940 271448 115992 271454
rect 197360 271448 197412 271454
rect 115940 271390 115992 271396
rect 183466 271416 183522 271425
rect 113548 271380 113600 271386
rect 197360 271390 197412 271396
rect 183466 271351 183522 271360
rect 113548 271322 113600 271328
rect 183480 271318 183508 271351
rect 197372 271318 197400 271390
rect 110420 271312 110472 271318
rect 106278 271280 106334 271289
rect 104900 271244 104952 271250
rect 110420 271254 110472 271260
rect 183468 271312 183520 271318
rect 183468 271254 183520 271260
rect 197360 271312 197412 271318
rect 197360 271254 197412 271260
rect 106278 271215 106334 271224
rect 104900 271186 104952 271192
rect 103520 271176 103572 271182
rect 103520 271118 103572 271124
rect 100760 271108 100812 271114
rect 100760 271050 100812 271056
rect 104898 271008 104954 271017
rect 104898 270943 104954 270952
rect 96618 270872 96674 270881
rect 96618 270807 96674 270816
rect 92478 270736 92534 270745
rect 92478 270671 92534 270680
rect 92492 270094 92520 270671
rect 92480 270088 92532 270094
rect 92480 270030 92532 270036
rect 91192 269748 91244 269754
rect 91192 269690 91244 269696
rect 88248 268388 88300 268394
rect 88248 268330 88300 268336
rect 83464 252000 83516 252006
rect 83464 251942 83516 251948
rect 96632 251938 96660 270807
rect 103702 270600 103758 270609
rect 102784 270564 102836 270570
rect 103702 270535 103758 270544
rect 102784 270506 102836 270512
rect 68376 251932 68428 251938
rect 68376 251874 68428 251880
rect 96620 251932 96672 251938
rect 96620 251874 96672 251880
rect 68388 250510 68416 251874
rect 102796 251870 102824 270506
rect 103716 269890 103744 270535
rect 103704 269884 103756 269890
rect 103704 269826 103756 269832
rect 104912 269822 104940 270943
rect 106292 269958 106320 271215
rect 183468 271176 183520 271182
rect 128358 271144 128414 271153
rect 128358 271079 128414 271088
rect 183466 271144 183468 271153
rect 183520 271144 183522 271153
rect 183466 271079 183522 271088
rect 115938 270872 115994 270881
rect 115938 270807 115994 270816
rect 106370 270600 106426 270609
rect 106370 270535 106426 270544
rect 107658 270600 107714 270609
rect 107658 270535 107714 270544
rect 110418 270600 110474 270609
rect 110418 270535 110474 270544
rect 113178 270600 113234 270609
rect 113178 270535 113180 270544
rect 106280 269952 106332 269958
rect 106280 269894 106332 269900
rect 104900 269816 104952 269822
rect 104900 269758 104952 269764
rect 106384 269618 106412 270535
rect 107672 269686 107700 270535
rect 110432 270298 110460 270535
rect 113232 270535 113234 270544
rect 114466 270600 114522 270609
rect 114466 270535 114522 270544
rect 115846 270600 115902 270609
rect 115846 270535 115902 270544
rect 113180 270506 113232 270512
rect 110420 270292 110472 270298
rect 110420 270234 110472 270240
rect 114480 269822 114508 270535
rect 115860 269890 115888 270535
rect 115952 270434 115980 270807
rect 115940 270428 115992 270434
rect 115940 270370 115992 270376
rect 115848 269884 115900 269890
rect 115848 269826 115900 269832
rect 114468 269816 114520 269822
rect 114468 269758 114520 269764
rect 107660 269680 107712 269686
rect 107660 269622 107712 269628
rect 106372 269612 106424 269618
rect 106372 269554 106424 269560
rect 128372 268326 128400 271079
rect 147678 270872 147734 270881
rect 147678 270807 147734 270816
rect 147692 270502 147720 270807
rect 147680 270496 147732 270502
rect 147680 270438 147732 270444
rect 196716 269884 196768 269890
rect 196716 269826 196768 269832
rect 196624 269816 196676 269822
rect 196624 269758 196676 269764
rect 128360 268320 128412 268326
rect 128360 268262 128412 268268
rect 180156 253360 180208 253366
rect 180154 253328 180156 253337
rect 180208 253328 180210 253337
rect 180154 253263 180210 253272
rect 179328 253224 179380 253230
rect 179326 253192 179328 253201
rect 179380 253192 179382 253201
rect 179326 253127 179382 253136
rect 191746 252648 191802 252657
rect 191746 252583 191748 252592
rect 191800 252583 191802 252592
rect 191748 252554 191800 252560
rect 102784 251864 102836 251870
rect 102784 251806 102836 251812
rect 68376 250504 68428 250510
rect 68376 250446 68428 250452
rect 101036 167000 101088 167006
rect 101036 166942 101088 166948
rect 98460 166932 98512 166938
rect 98460 166874 98512 166880
rect 98472 166705 98500 166874
rect 101048 166705 101076 166942
rect 105820 166864 105872 166870
rect 105820 166806 105872 166812
rect 138478 166832 138534 166841
rect 105832 166705 105860 166806
rect 108212 166796 108264 166802
rect 138478 166767 138534 166776
rect 143538 166832 143594 166841
rect 143538 166767 143594 166776
rect 145930 166832 145986 166841
rect 145930 166767 145986 166776
rect 108212 166738 108264 166744
rect 108224 166705 108252 166738
rect 138492 166734 138520 166767
rect 138480 166728 138532 166734
rect 98458 166696 98514 166705
rect 98458 166631 98514 166640
rect 101034 166696 101090 166705
rect 101034 166631 101090 166640
rect 105818 166696 105874 166705
rect 105818 166631 105874 166640
rect 108210 166696 108266 166705
rect 138480 166670 138532 166676
rect 143552 166666 143580 166767
rect 108210 166631 108266 166640
rect 143540 166660 143592 166666
rect 143540 166602 143592 166608
rect 145944 166598 145972 166767
rect 163318 166696 163374 166705
rect 163318 166631 163374 166640
rect 165894 166696 165950 166705
rect 165894 166631 165950 166640
rect 145932 166592 145984 166598
rect 113270 166560 113326 166569
rect 145932 166534 145984 166540
rect 150898 166560 150954 166569
rect 113270 166495 113326 166504
rect 150898 166495 150900 166504
rect 96066 166288 96122 166297
rect 96066 166223 96068 166232
rect 96120 166223 96122 166232
rect 96068 166194 96120 166200
rect 113284 165646 113312 166495
rect 150952 166495 150954 166504
rect 153290 166560 153346 166569
rect 153290 166495 153346 166504
rect 150900 166466 150952 166472
rect 153304 166462 153332 166495
rect 153292 166456 153344 166462
rect 153292 166398 153344 166404
rect 163332 166394 163360 166631
rect 163320 166388 163372 166394
rect 163320 166330 163372 166336
rect 165908 166326 165936 166631
rect 165896 166320 165948 166326
rect 165896 166262 165948 166268
rect 113272 165640 113324 165646
rect 81438 165608 81494 165617
rect 81438 165543 81494 165552
rect 84290 165608 84346 165617
rect 84290 165543 84346 165552
rect 89902 165608 89958 165617
rect 89902 165543 89958 165552
rect 91098 165608 91154 165617
rect 91098 165543 91154 165552
rect 95238 165608 95294 165617
rect 95238 165543 95294 165552
rect 99378 165608 99434 165617
rect 99378 165543 99434 165552
rect 103518 165608 103574 165617
rect 103518 165543 103574 165552
rect 109682 165608 109738 165617
rect 109682 165543 109738 165552
rect 110878 165608 110934 165617
rect 110878 165543 110934 165552
rect 111154 165608 111210 165617
rect 111154 165543 111210 165552
rect 111890 165608 111946 165617
rect 113272 165582 113324 165588
rect 113546 165608 113602 165617
rect 111890 165543 111946 165552
rect 113546 165543 113602 165552
rect 115938 165608 115994 165617
rect 115938 165543 115994 165552
rect 116398 165608 116454 165617
rect 116398 165543 116454 165552
rect 117870 165608 117926 165617
rect 117870 165543 117926 165552
rect 118330 165608 118386 165617
rect 118330 165543 118386 165552
rect 120906 165608 120962 165617
rect 120906 165543 120962 165552
rect 123482 165608 123538 165617
rect 123482 165543 123538 165552
rect 125874 165608 125930 165617
rect 125874 165543 125930 165552
rect 128358 165608 128414 165617
rect 128358 165543 128414 165552
rect 129738 165608 129794 165617
rect 129738 165543 129794 165552
rect 132498 165608 132554 165617
rect 132498 165543 132500 165552
rect 76010 164384 76066 164393
rect 76010 164319 76066 164328
rect 75918 164248 75974 164257
rect 75918 164183 75974 164192
rect 60096 146328 60148 146334
rect 60096 146270 60148 146276
rect 60108 146062 60136 146270
rect 60924 146124 60976 146130
rect 60924 146066 60976 146072
rect 60096 146056 60148 146062
rect 60096 145998 60148 146004
rect 60936 145314 60964 146066
rect 75932 145382 75960 164183
rect 76024 145450 76052 164319
rect 77298 164248 77354 164257
rect 77298 164183 77354 164192
rect 78678 164248 78734 164257
rect 78678 164183 78734 164192
rect 80058 164248 80114 164257
rect 80058 164183 80114 164192
rect 77312 145518 77340 164183
rect 78692 148782 78720 164183
rect 78680 148776 78732 148782
rect 78680 148718 78732 148724
rect 80072 148714 80100 164183
rect 80060 148708 80112 148714
rect 80060 148650 80112 148656
rect 81452 148646 81480 165543
rect 83464 164484 83516 164490
rect 83464 164426 83516 164432
rect 82818 164248 82874 164257
rect 82818 164183 82874 164192
rect 81440 148640 81492 148646
rect 81440 148582 81492 148588
rect 82832 145926 82860 164183
rect 83476 148850 83504 164426
rect 84198 164248 84254 164257
rect 84198 164183 84254 164192
rect 83464 148844 83516 148850
rect 83464 148786 83516 148792
rect 82820 145920 82872 145926
rect 82820 145862 82872 145868
rect 84212 145858 84240 164183
rect 84304 145994 84332 165543
rect 89916 164830 89944 165543
rect 89904 164824 89956 164830
rect 88338 164792 88394 164801
rect 89904 164766 89956 164772
rect 88338 164727 88340 164736
rect 88392 164727 88394 164736
rect 88340 164698 88392 164704
rect 88984 164348 89036 164354
rect 88984 164290 89036 164296
rect 85578 164248 85634 164257
rect 85578 164183 85634 164192
rect 86958 164248 87014 164257
rect 86958 164183 87014 164192
rect 88430 164248 88486 164257
rect 88430 164183 88486 164192
rect 85592 146198 85620 164183
rect 85580 146192 85632 146198
rect 85580 146134 85632 146140
rect 86972 146130 87000 164183
rect 86960 146124 87012 146130
rect 86960 146066 87012 146072
rect 84292 145988 84344 145994
rect 84292 145930 84344 145936
rect 84200 145852 84252 145858
rect 84200 145794 84252 145800
rect 88444 145790 88472 164183
rect 88996 148578 89024 164290
rect 89810 164248 89866 164257
rect 89810 164183 89866 164192
rect 88984 148572 89036 148578
rect 88984 148514 89036 148520
rect 89824 146062 89852 164183
rect 89812 146056 89864 146062
rect 91112 146033 91140 165543
rect 91190 164248 91246 164257
rect 91190 164183 91246 164192
rect 92478 164248 92534 164257
rect 92478 164183 92534 164192
rect 93858 164248 93914 164257
rect 93858 164183 93914 164192
rect 89812 145998 89864 146004
rect 91098 146024 91154 146033
rect 91098 145959 91154 145968
rect 88432 145784 88484 145790
rect 88432 145726 88484 145732
rect 91204 145722 91232 164183
rect 92492 146266 92520 164183
rect 92480 146260 92532 146266
rect 92480 146202 92532 146208
rect 91192 145716 91244 145722
rect 91192 145658 91244 145664
rect 93872 145654 93900 164183
rect 95252 163810 95280 165543
rect 97264 164416 97316 164422
rect 97264 164358 97316 164364
rect 96618 164248 96674 164257
rect 96618 164183 96674 164192
rect 95240 163804 95292 163810
rect 95240 163746 95292 163752
rect 96632 145897 96660 164183
rect 96618 145888 96674 145897
rect 96618 145823 96674 145832
rect 97276 145761 97304 164358
rect 97998 164248 98054 164257
rect 97998 164183 98054 164192
rect 98012 163742 98040 164183
rect 98000 163736 98052 163742
rect 98000 163678 98052 163684
rect 97262 145752 97318 145761
rect 97262 145687 97318 145696
rect 93860 145648 93912 145654
rect 99392 145625 99420 165543
rect 103532 164966 103560 165543
rect 103520 164960 103572 164966
rect 103520 164902 103572 164908
rect 104898 164928 104954 164937
rect 104898 164863 104900 164872
rect 104952 164863 104954 164872
rect 107566 164928 107622 164937
rect 107622 164886 107700 164914
rect 107566 164863 107622 164872
rect 104900 164834 104952 164840
rect 106278 164792 106334 164801
rect 106278 164727 106334 164736
rect 100758 164520 100814 164529
rect 100758 164455 100814 164464
rect 100772 164422 100800 164455
rect 100760 164416 100812 164422
rect 100760 164358 100812 164364
rect 106292 164354 106320 164727
rect 106280 164348 106332 164354
rect 106280 164290 106332 164296
rect 100758 164248 100814 164257
rect 100758 164183 100814 164192
rect 102138 164248 102194 164257
rect 102138 164183 102194 164192
rect 103610 164248 103666 164257
rect 103610 164183 103666 164192
rect 93860 145590 93912 145596
rect 99378 145616 99434 145625
rect 100772 145586 100800 164183
rect 102152 148986 102180 164183
rect 103624 149054 103652 164183
rect 103612 149048 103664 149054
rect 103612 148990 103664 148996
rect 102140 148980 102192 148986
rect 102140 148922 102192 148928
rect 107672 148510 107700 164886
rect 107750 164520 107806 164529
rect 107750 164455 107752 164464
rect 107804 164455 107806 164464
rect 107752 164426 107804 164432
rect 109696 164014 109724 165543
rect 110892 164082 110920 165543
rect 110880 164076 110932 164082
rect 110880 164018 110932 164024
rect 109684 164008 109736 164014
rect 109684 163950 109736 163956
rect 111168 163674 111196 165543
rect 111156 163668 111208 163674
rect 111156 163610 111208 163616
rect 111904 163606 111932 165543
rect 113560 165034 113588 165543
rect 115952 165170 115980 165543
rect 115940 165164 115992 165170
rect 115940 165106 115992 165112
rect 113548 165028 113600 165034
rect 113548 164970 113600 164976
rect 116032 164960 116084 164966
rect 114466 164928 114522 164937
rect 114522 164898 114600 164914
rect 116032 164902 116084 164908
rect 114522 164892 114612 164898
rect 114522 164886 114560 164892
rect 114466 164863 114522 164872
rect 114560 164834 114612 164840
rect 111892 163600 111944 163606
rect 111892 163542 111944 163548
rect 107660 148504 107712 148510
rect 107660 148446 107712 148452
rect 114572 148374 114600 164834
rect 116044 164529 116072 164902
rect 116030 164520 116086 164529
rect 116030 164455 116086 164464
rect 116044 148442 116072 164455
rect 116412 164218 116440 165543
rect 116400 164212 116452 164218
rect 116400 164154 116452 164160
rect 117884 164150 117912 165543
rect 118344 165102 118372 165543
rect 120920 165238 120948 165543
rect 123496 165306 123524 165543
rect 125888 165374 125916 165543
rect 128372 165442 128400 165543
rect 129752 165510 129780 165543
rect 132552 165543 132554 165552
rect 183190 165608 183246 165617
rect 183190 165543 183246 165552
rect 132500 165514 132552 165520
rect 129740 165504 129792 165510
rect 129740 165446 129792 165452
rect 128360 165436 128412 165442
rect 128360 165378 128412 165384
rect 125876 165368 125928 165374
rect 125876 165310 125928 165316
rect 123484 165300 123536 165306
rect 123484 165242 123536 165248
rect 120908 165232 120960 165238
rect 120908 165174 120960 165180
rect 183204 165170 183232 165543
rect 183192 165164 183244 165170
rect 183192 165106 183244 165112
rect 118332 165096 118384 165102
rect 118332 165038 118384 165044
rect 118882 165064 118938 165073
rect 118882 164999 118938 165008
rect 183466 165064 183522 165073
rect 183466 164999 183468 165008
rect 117872 164144 117924 164150
rect 117872 164086 117924 164092
rect 118896 163538 118924 164999
rect 183520 164999 183522 165008
rect 183468 164970 183520 164976
rect 118884 163532 118936 163538
rect 118884 163474 118936 163480
rect 116032 148436 116084 148442
rect 116032 148378 116084 148384
rect 114560 148368 114612 148374
rect 114560 148310 114612 148316
rect 179052 146260 179104 146266
rect 179052 146202 179104 146208
rect 99378 145551 99434 145560
rect 100760 145580 100812 145586
rect 100760 145522 100812 145528
rect 77300 145512 77352 145518
rect 77300 145454 77352 145460
rect 76012 145444 76064 145450
rect 76012 145386 76064 145392
rect 75920 145376 75972 145382
rect 75920 145318 75972 145324
rect 60924 145308 60976 145314
rect 60924 145250 60976 145256
rect 179064 144945 179092 146202
rect 179696 146192 179748 146198
rect 179696 146134 179748 146140
rect 179708 144945 179736 146134
rect 183480 145654 183508 164970
rect 196636 164898 196664 269758
rect 196728 164966 196756 269826
rect 197372 165170 197400 271254
rect 197556 258074 197584 358838
rect 197740 358834 197768 359518
rect 197728 358828 197780 358834
rect 197728 358770 197780 358776
rect 197740 358170 197768 358770
rect 197464 258046 197584 258074
rect 197648 358142 197768 358170
rect 197464 253366 197492 258046
rect 197452 253360 197504 253366
rect 197452 253302 197504 253308
rect 197360 165164 197412 165170
rect 197360 165106 197412 165112
rect 196716 164960 196768 164966
rect 196716 164902 196768 164908
rect 196624 164892 196676 164898
rect 196624 164834 196676 164840
rect 183468 145648 183520 145654
rect 183468 145590 183520 145596
rect 191748 145580 191800 145586
rect 191748 145522 191800 145528
rect 191760 145489 191788 145522
rect 191746 145480 191802 145489
rect 191746 145415 191802 145424
rect 179050 144936 179106 144945
rect 179050 144871 179106 144880
rect 179694 144936 179750 144945
rect 179694 144871 179750 144880
rect 77116 59832 77168 59838
rect 77114 59800 77116 59809
rect 77168 59800 77170 59809
rect 77114 59735 77170 59744
rect 83094 59800 83150 59809
rect 83094 59735 83150 59744
rect 84198 59800 84254 59809
rect 84198 59735 84200 59744
rect 83108 59634 83136 59735
rect 84252 59735 84254 59744
rect 99470 59800 99526 59809
rect 99470 59735 99526 59744
rect 102782 59800 102838 59809
rect 102782 59735 102838 59744
rect 107566 59800 107622 59809
rect 107566 59735 107622 59744
rect 84200 59706 84252 59712
rect 83096 59628 83148 59634
rect 83096 59570 83148 59576
rect 99484 59566 99512 59735
rect 100760 59696 100812 59702
rect 100758 59664 100760 59673
rect 100812 59664 100814 59673
rect 100758 59599 100814 59608
rect 99472 59560 99524 59566
rect 99472 59502 99524 59508
rect 102796 59498 102824 59735
rect 103886 59664 103942 59673
rect 103886 59599 103942 59608
rect 102784 59492 102836 59498
rect 102784 59434 102836 59440
rect 85394 59392 85450 59401
rect 85394 59327 85396 59336
rect 85448 59327 85450 59336
rect 95882 59392 95938 59401
rect 95882 59327 95938 59336
rect 98090 59392 98146 59401
rect 98090 59327 98146 59336
rect 85396 59298 85448 59304
rect 95896 59294 95924 59327
rect 95884 59288 95936 59294
rect 95884 59230 95936 59236
rect 98104 59226 98132 59327
rect 98092 59220 98144 59226
rect 98092 59162 98144 59168
rect 103900 59090 103928 59599
rect 107580 59430 107608 59735
rect 114374 59664 114430 59673
rect 114374 59599 114430 59608
rect 143538 59664 143594 59673
rect 143538 59599 143594 59608
rect 107568 59424 107620 59430
rect 105266 59392 105322 59401
rect 105266 59327 105322 59336
rect 106370 59392 106426 59401
rect 107568 59366 107620 59372
rect 106370 59327 106426 59336
rect 103888 59084 103940 59090
rect 103888 59026 103940 59032
rect 105280 59022 105308 59327
rect 106384 59158 106412 59327
rect 106372 59152 106424 59158
rect 106372 59094 106424 59100
rect 105268 59016 105320 59022
rect 105268 58958 105320 58964
rect 114388 58954 114416 59599
rect 138386 59120 138442 59129
rect 138386 59055 138442 59064
rect 114376 58948 114428 58954
rect 114376 58890 114428 58896
rect 138400 58886 138428 59055
rect 138388 58880 138440 58886
rect 138388 58822 138440 58828
rect 143552 58818 143580 59599
rect 148506 59256 148562 59265
rect 148506 59191 148562 59200
rect 150898 59256 150954 59265
rect 150898 59191 150954 59200
rect 143540 58812 143592 58818
rect 143540 58754 143592 58760
rect 148520 58682 148548 59191
rect 150912 58750 150940 59191
rect 150900 58744 150952 58750
rect 150900 58686 150952 58692
rect 148508 58676 148560 58682
rect 148508 58618 148560 58624
rect 76010 57896 76066 57905
rect 76010 57831 76066 57840
rect 78218 57896 78274 57905
rect 78218 57831 78274 57840
rect 78678 57896 78734 57905
rect 78678 57831 78734 57840
rect 80426 57896 80482 57905
rect 80426 57831 80482 57840
rect 81438 57896 81494 57905
rect 81438 57831 81494 57840
rect 86498 57896 86554 57905
rect 86498 57831 86554 57840
rect 86958 57896 87014 57905
rect 86958 57831 87014 57840
rect 88338 57896 88394 57905
rect 88338 57831 88394 57840
rect 89994 57896 90050 57905
rect 89994 57831 90050 57840
rect 90730 57896 90786 57905
rect 90730 57831 90786 57840
rect 91190 57896 91246 57905
rect 91190 57831 91246 57840
rect 92202 57896 92258 57905
rect 92202 57831 92258 57840
rect 92478 57896 92534 57905
rect 92478 57831 92534 57840
rect 93674 57896 93730 57905
rect 93674 57831 93730 57840
rect 94410 57896 94466 57905
rect 94410 57831 94466 57840
rect 98458 57896 98514 57905
rect 98458 57831 98514 57840
rect 101770 57896 101826 57905
rect 101770 57831 101826 57840
rect 108578 57896 108634 57905
rect 108578 57831 108634 57840
rect 109498 57896 109554 57905
rect 109498 57831 109554 57840
rect 111154 57896 111210 57905
rect 111154 57831 111210 57840
rect 113546 57896 113602 57905
rect 113546 57831 113602 57840
rect 116490 57896 116546 57905
rect 116490 57831 116546 57840
rect 117962 57896 118018 57905
rect 117962 57831 118018 57840
rect 120722 57896 120778 57905
rect 120722 57831 120778 57840
rect 123482 57896 123538 57905
rect 123482 57831 123538 57840
rect 130842 57896 130898 57905
rect 130842 57831 130898 57840
rect 145562 57896 145618 57905
rect 145562 57831 145564 57840
rect 60004 57452 60056 57458
rect 60004 57394 60056 57400
rect 76024 57186 76052 57831
rect 76012 57180 76064 57186
rect 76012 57122 76064 57128
rect 59728 56296 59780 56302
rect 59728 56238 59780 56244
rect 78232 55962 78260 57831
rect 78220 55956 78272 55962
rect 78220 55898 78272 55904
rect 58992 54936 59044 54942
rect 58992 54878 59044 54884
rect 78692 54670 78720 57831
rect 80440 56030 80468 57831
rect 80428 56024 80480 56030
rect 80428 55966 80480 55972
rect 81452 54738 81480 57831
rect 86512 56166 86540 57831
rect 86500 56160 86552 56166
rect 86500 56102 86552 56108
rect 86972 54806 87000 57831
rect 88352 54874 88380 57831
rect 88432 57384 88484 57390
rect 88432 57326 88484 57332
rect 88444 57089 88472 57326
rect 88430 57080 88486 57089
rect 88430 57015 88486 57024
rect 90008 56098 90036 57831
rect 90744 57254 90772 57831
rect 90732 57248 90784 57254
rect 90732 57190 90784 57196
rect 89996 56092 90048 56098
rect 89996 56034 90048 56040
rect 91204 55010 91232 57831
rect 92216 56234 92244 57831
rect 92204 56228 92256 56234
rect 92204 56170 92256 56176
rect 91192 55004 91244 55010
rect 91192 54946 91244 54952
rect 92492 54942 92520 57831
rect 93688 57322 93716 57831
rect 93676 57316 93728 57322
rect 93676 57258 93728 57264
rect 94424 56302 94452 57831
rect 98472 57458 98500 57831
rect 98642 57488 98698 57497
rect 98460 57452 98512 57458
rect 98642 57423 98698 57432
rect 98460 57394 98512 57400
rect 98656 57225 98684 57423
rect 98642 57216 98698 57225
rect 98642 57151 98698 57160
rect 101784 56370 101812 57831
rect 108592 57526 108620 57831
rect 108580 57520 108632 57526
rect 108580 57462 108632 57468
rect 109512 56438 109540 57831
rect 111168 56506 111196 57831
rect 113560 57662 113588 57831
rect 113548 57656 113600 57662
rect 113548 57598 113600 57604
rect 114558 57624 114614 57633
rect 114558 57559 114614 57568
rect 111798 57488 111854 57497
rect 111798 57423 111854 57432
rect 113178 57488 113234 57497
rect 113178 57423 113234 57432
rect 111156 56500 111208 56506
rect 111156 56442 111208 56448
rect 109500 56432 109552 56438
rect 109500 56374 109552 56380
rect 101772 56364 101824 56370
rect 101772 56306 101824 56312
rect 94412 56296 94464 56302
rect 94412 56238 94464 56244
rect 111812 55146 111840 57423
rect 111800 55140 111852 55146
rect 111800 55082 111852 55088
rect 113192 55078 113220 57423
rect 114572 55214 114600 57559
rect 116504 56137 116532 57831
rect 117976 57594 118004 57831
rect 120736 57730 120764 57831
rect 120724 57724 120776 57730
rect 120724 57666 120776 57672
rect 118698 57624 118754 57633
rect 117964 57588 118016 57594
rect 118698 57559 118754 57568
rect 117964 57530 118016 57536
rect 116490 56128 116546 56137
rect 116490 56063 116546 56072
rect 114560 55208 114612 55214
rect 114560 55150 114612 55156
rect 113180 55072 113232 55078
rect 113180 55014 113232 55020
rect 92480 54936 92532 54942
rect 92480 54878 92532 54884
rect 88340 54868 88392 54874
rect 88340 54810 88392 54816
rect 86960 54800 87012 54806
rect 118712 54777 118740 57559
rect 123496 56574 123524 57831
rect 130856 57798 130884 57831
rect 145616 57831 145618 57840
rect 153290 57896 153346 57905
rect 153290 57831 153346 57840
rect 183466 57896 183522 57905
rect 183466 57831 183468 57840
rect 145564 57802 145616 57808
rect 130844 57792 130896 57798
rect 130844 57734 130896 57740
rect 123484 56568 123536 56574
rect 123484 56510 123536 56516
rect 153304 56273 153332 57831
rect 183520 57831 183522 57840
rect 183468 57802 183520 57808
rect 197372 57798 197400 165106
rect 197464 146198 197492 253302
rect 197648 253230 197676 358142
rect 197728 358080 197780 358086
rect 197728 358022 197780 358028
rect 197740 271454 197768 358022
rect 197728 271448 197780 271454
rect 197728 271390 197780 271396
rect 197636 253224 197688 253230
rect 197636 253166 197688 253172
rect 197648 238754 197676 253166
rect 197556 238726 197676 238754
rect 197556 146266 197584 238726
rect 198004 175976 198056 175982
rect 198004 175918 198056 175924
rect 197544 146260 197596 146266
rect 197544 146202 197596 146208
rect 197452 146192 197504 146198
rect 197452 146134 197504 146140
rect 197452 145648 197504 145654
rect 197452 145590 197504 145596
rect 197464 57866 197492 145590
rect 198016 145586 198044 175918
rect 198004 145580 198056 145586
rect 198004 145522 198056 145528
rect 198568 59022 198596 380967
rect 198660 379098 198688 396607
rect 198648 379092 198700 379098
rect 198648 379034 198700 379040
rect 198752 364334 198780 460119
rect 198844 376718 198872 493037
rect 198924 492108 198976 492114
rect 198924 492050 198976 492056
rect 198936 400466 198964 492050
rect 199108 476808 199160 476814
rect 199108 476750 199160 476756
rect 199016 464432 199068 464438
rect 199016 464374 199068 464380
rect 199028 400586 199056 464374
rect 199120 400586 199148 476750
rect 199200 475380 199252 475386
rect 199200 475322 199252 475328
rect 199016 400580 199068 400586
rect 199016 400522 199068 400528
rect 199108 400580 199160 400586
rect 199108 400522 199160 400528
rect 198936 400438 199148 400466
rect 199016 400376 199068 400382
rect 198922 400344 198978 400353
rect 199016 400318 199068 400324
rect 198922 400279 198978 400288
rect 198936 400246 198964 400279
rect 198924 400240 198976 400246
rect 198924 400182 198976 400188
rect 198922 395312 198978 395321
rect 198922 395247 198978 395256
rect 198936 378146 198964 395247
rect 198924 378140 198976 378146
rect 198924 378082 198976 378088
rect 198832 376712 198884 376718
rect 198832 376654 198884 376660
rect 199028 376310 199056 400318
rect 199120 397458 199148 400438
rect 199108 397452 199160 397458
rect 199108 397394 199160 397400
rect 199212 397361 199240 475322
rect 199198 397352 199254 397361
rect 199198 397287 199254 397296
rect 199304 382974 199332 493037
rect 199384 490680 199436 490686
rect 199384 490622 199436 490628
rect 199292 382968 199344 382974
rect 199292 382910 199344 382916
rect 199396 377466 199424 490622
rect 199476 474020 199528 474026
rect 199476 473962 199528 473968
rect 199488 422294 199516 473962
rect 199488 422266 199608 422294
rect 199580 398313 199608 422266
rect 199566 398304 199622 398313
rect 199566 398239 199622 398248
rect 199474 397352 199530 397361
rect 199474 397287 199530 397296
rect 199384 377460 199436 377466
rect 199384 377402 199436 377408
rect 199016 376304 199068 376310
rect 199016 376246 199068 376252
rect 199384 375284 199436 375290
rect 199384 375226 199436 375232
rect 199396 374678 199424 375226
rect 199384 374672 199436 374678
rect 199384 374614 199436 374620
rect 198752 364306 198872 364334
rect 198844 353161 198872 364306
rect 198830 353152 198886 353161
rect 198830 353087 198886 353096
rect 198738 291680 198794 291689
rect 198738 291615 198794 291624
rect 198648 253904 198700 253910
rect 198648 253846 198700 253852
rect 198660 252618 198688 253846
rect 198648 252612 198700 252618
rect 198648 252554 198700 252560
rect 198660 175982 198688 252554
rect 198752 184929 198780 291615
rect 198844 246265 198872 353087
rect 199198 292768 199254 292777
rect 199198 292703 199254 292712
rect 198922 291000 198978 291009
rect 198922 290935 198978 290944
rect 198830 246256 198886 246265
rect 198830 246191 198886 246200
rect 198738 184920 198794 184929
rect 198738 184855 198794 184864
rect 198738 183560 198794 183569
rect 198738 183495 198794 183504
rect 198648 175976 198700 175982
rect 198648 175918 198700 175924
rect 198752 76401 198780 183495
rect 198844 139233 198872 246191
rect 198936 183569 198964 290935
rect 199106 289776 199162 289785
rect 199106 289711 199162 289720
rect 199120 288833 199148 289711
rect 199106 288824 199162 288833
rect 199106 288759 199162 288768
rect 199014 288416 199070 288425
rect 199014 288351 199070 288360
rect 199028 287609 199056 288351
rect 199014 287600 199070 287609
rect 199014 287535 199070 287544
rect 198922 183560 198978 183569
rect 198922 183495 198978 183504
rect 198922 182064 198978 182073
rect 198922 181999 198978 182008
rect 198830 139224 198886 139233
rect 198830 139159 198886 139168
rect 198738 76392 198794 76401
rect 198738 76327 198794 76336
rect 198936 74905 198964 181999
rect 199028 180713 199056 287535
rect 199120 182073 199148 288759
rect 199212 209774 199240 292703
rect 199396 291689 199424 374614
rect 199488 369170 199516 397287
rect 199580 375290 199608 398239
rect 199764 380322 199792 493037
rect 200120 468580 200172 468586
rect 200120 468522 200172 468528
rect 199844 400580 199896 400586
rect 199844 400522 199896 400528
rect 199856 394641 199884 400522
rect 199842 394632 199898 394641
rect 199842 394567 199898 394576
rect 199752 380316 199804 380322
rect 199752 380258 199804 380264
rect 199660 378140 199712 378146
rect 199660 378082 199712 378088
rect 199568 375284 199620 375290
rect 199568 375226 199620 375232
rect 199568 371204 199620 371210
rect 199568 371146 199620 371152
rect 199476 369164 199528 369170
rect 199476 369106 199528 369112
rect 199382 291680 199438 291689
rect 199382 291615 199438 291624
rect 199488 291009 199516 369106
rect 199580 292777 199608 371146
rect 199672 363662 199700 378082
rect 199752 377052 199804 377058
rect 199752 376994 199804 377000
rect 199764 371210 199792 376994
rect 199752 371204 199804 371210
rect 199752 371146 199804 371152
rect 199856 364334 199884 394567
rect 199764 364306 199884 364334
rect 199660 363656 199712 363662
rect 199660 363598 199712 363604
rect 199566 292768 199622 292777
rect 199566 292703 199622 292712
rect 199474 291000 199530 291009
rect 199474 290935 199530 290944
rect 199672 289785 199700 363598
rect 199764 362234 199792 364306
rect 199752 362228 199804 362234
rect 199752 362170 199804 362176
rect 199658 289776 199714 289785
rect 199658 289711 199714 289720
rect 199764 288425 199792 362170
rect 199750 288416 199806 288425
rect 199750 288351 199806 288360
rect 200132 271862 200160 468522
rect 200224 377942 200252 493037
rect 200684 490618 200712 493037
rect 200764 490952 200816 490958
rect 200762 490920 200764 490929
rect 200816 490920 200818 490929
rect 200762 490855 200818 490864
rect 200672 490612 200724 490618
rect 200672 490554 200724 490560
rect 200580 490476 200632 490482
rect 200580 490418 200632 490424
rect 200592 490385 200620 490418
rect 200578 490376 200634 490385
rect 200578 490311 200634 490320
rect 200304 487960 200356 487966
rect 200304 487902 200356 487908
rect 200316 380254 200344 487902
rect 200856 476944 200908 476950
rect 200856 476886 200908 476892
rect 200396 471572 200448 471578
rect 200396 471514 200448 471520
rect 200304 380248 200356 380254
rect 200304 380190 200356 380196
rect 200212 377936 200264 377942
rect 200212 377878 200264 377884
rect 200408 377126 200436 471514
rect 200764 471164 200816 471170
rect 200764 471106 200816 471112
rect 200488 465860 200540 465866
rect 200488 465802 200540 465808
rect 200500 379982 200528 465802
rect 200580 465044 200632 465050
rect 200580 464986 200632 464992
rect 200592 381002 200620 464986
rect 200580 380996 200632 381002
rect 200580 380938 200632 380944
rect 200488 379976 200540 379982
rect 200488 379918 200540 379924
rect 200396 377120 200448 377126
rect 200396 377062 200448 377068
rect 200776 284306 200804 471106
rect 200764 284300 200816 284306
rect 200764 284242 200816 284248
rect 200764 282464 200816 282470
rect 200764 282406 200816 282412
rect 200120 271856 200172 271862
rect 200120 271798 200172 271804
rect 200776 253910 200804 282406
rect 200868 271726 200896 476886
rect 200948 468376 201000 468382
rect 200948 468318 201000 468324
rect 200960 272542 200988 468318
rect 201052 380254 201080 493037
rect 201406 381032 201462 381041
rect 201406 380967 201462 380976
rect 201040 380248 201092 380254
rect 201040 380190 201092 380196
rect 200948 272536 201000 272542
rect 200948 272478 201000 272484
rect 200856 271720 200908 271726
rect 200856 271662 200908 271668
rect 200764 253904 200816 253910
rect 200764 253846 200816 253852
rect 199212 209746 199332 209774
rect 199304 186425 199332 209746
rect 199290 186416 199346 186425
rect 199290 186351 199346 186360
rect 199198 184920 199254 184929
rect 199198 184855 199254 184864
rect 199106 182064 199162 182073
rect 199106 181999 199162 182008
rect 199014 180704 199070 180713
rect 199014 180639 199070 180648
rect 199028 171134 199056 180639
rect 199028 171106 199148 171134
rect 198922 74896 198978 74905
rect 198922 74831 198978 74840
rect 199120 73681 199148 171106
rect 199212 77761 199240 184855
rect 199304 79393 199332 186351
rect 199290 79384 199346 79393
rect 199290 79319 199346 79328
rect 199198 77752 199254 77761
rect 199198 77687 199254 77696
rect 199106 73672 199162 73681
rect 199106 73607 199162 73616
rect 198556 59016 198608 59022
rect 198556 58958 198608 58964
rect 201420 58886 201448 380967
rect 201512 380186 201540 493037
rect 201972 491230 202000 493037
rect 202064 493023 202446 493051
rect 201960 491224 202012 491230
rect 201960 491166 202012 491172
rect 201592 491088 201644 491094
rect 201590 491056 201592 491065
rect 201644 491056 201646 491065
rect 201590 490991 201646 491000
rect 201684 491020 201736 491026
rect 201684 490962 201736 490968
rect 201696 490686 201724 490962
rect 201684 490680 201736 490686
rect 201684 490622 201736 490628
rect 202064 489914 202092 493023
rect 202892 490657 202920 493037
rect 202878 490648 202934 490657
rect 202878 490583 202934 490592
rect 203260 490346 203288 493037
rect 203352 493023 203734 493051
rect 203248 490340 203300 490346
rect 203248 490282 203300 490288
rect 203352 489914 203380 493023
rect 204076 490476 204128 490482
rect 204076 490418 204128 490424
rect 201604 489886 202092 489914
rect 203076 489886 203380 489914
rect 201604 380390 201632 489886
rect 202328 481024 202380 481030
rect 202328 480966 202380 480972
rect 202234 471336 202290 471345
rect 202234 471271 202290 471280
rect 201868 470620 201920 470626
rect 201868 470562 201920 470568
rect 201684 468512 201736 468518
rect 201684 468454 201736 468460
rect 201592 380384 201644 380390
rect 201592 380326 201644 380332
rect 201500 380180 201552 380186
rect 201500 380122 201552 380128
rect 201592 367804 201644 367810
rect 201592 367746 201644 367752
rect 201500 359508 201552 359514
rect 201500 359450 201552 359456
rect 201512 282878 201540 359450
rect 201500 282872 201552 282878
rect 201500 282814 201552 282820
rect 201512 282470 201540 282814
rect 201500 282464 201552 282470
rect 201500 282406 201552 282412
rect 201604 271182 201632 367746
rect 201696 271794 201724 468454
rect 201776 466540 201828 466546
rect 201776 466482 201828 466488
rect 201788 360194 201816 466482
rect 201880 377194 201908 470562
rect 202144 465588 202196 465594
rect 202144 465530 202196 465536
rect 202156 389162 202184 465530
rect 202144 389156 202196 389162
rect 202144 389098 202196 389104
rect 201868 377188 201920 377194
rect 201868 377130 201920 377136
rect 201776 360188 201828 360194
rect 201776 360130 201828 360136
rect 201684 271788 201736 271794
rect 201684 271730 201736 271736
rect 201592 271176 201644 271182
rect 201592 271118 201644 271124
rect 201604 258074 201632 271118
rect 201512 258046 201632 258074
rect 201512 165034 201540 258046
rect 202248 166870 202276 471271
rect 202340 271658 202368 480966
rect 202418 471472 202474 471481
rect 202418 471407 202474 471416
rect 202328 271652 202380 271658
rect 202328 271594 202380 271600
rect 202236 166864 202288 166870
rect 202236 166806 202288 166812
rect 202432 166734 202460 471407
rect 202880 471368 202932 471374
rect 202880 471310 202932 471316
rect 202512 465656 202564 465662
rect 202512 465598 202564 465604
rect 202524 270473 202552 465598
rect 202788 360868 202840 360874
rect 202788 360810 202840 360816
rect 202800 359514 202828 360810
rect 202788 359508 202840 359514
rect 202788 359450 202840 359456
rect 202510 270464 202566 270473
rect 202510 270399 202566 270408
rect 202892 269822 202920 471310
rect 202972 471300 203024 471306
rect 202972 471242 203024 471248
rect 202984 271522 203012 471242
rect 203076 418062 203104 489886
rect 203708 486600 203760 486606
rect 203708 486542 203760 486548
rect 203524 482316 203576 482322
rect 203524 482258 203576 482264
rect 203064 418056 203116 418062
rect 203064 417998 203116 418004
rect 203064 416084 203116 416090
rect 203064 416026 203116 416032
rect 203076 380458 203104 416026
rect 203064 380452 203116 380458
rect 203064 380394 203116 380400
rect 202972 271516 203024 271522
rect 202972 271458 203024 271464
rect 202880 269816 202932 269822
rect 202880 269758 202932 269764
rect 202420 166728 202472 166734
rect 202420 166670 202472 166676
rect 203536 165481 203564 482258
rect 203616 466200 203668 466206
rect 203616 466142 203668 466148
rect 203628 166462 203656 466142
rect 203720 271590 203748 486542
rect 203800 469124 203852 469130
rect 203800 469066 203852 469072
rect 203812 272678 203840 469066
rect 203892 466268 203944 466274
rect 203892 466210 203944 466216
rect 203904 282810 203932 466210
rect 204088 378962 204116 490418
rect 204180 379574 204208 493037
rect 204654 493023 204760 493051
rect 204444 491496 204496 491502
rect 204444 491438 204496 491444
rect 204260 490952 204312 490958
rect 204258 490920 204260 490929
rect 204312 490920 204314 490929
rect 204258 490855 204314 490864
rect 204260 490544 204312 490550
rect 204258 490512 204260 490521
rect 204312 490512 204314 490521
rect 204258 490447 204314 490456
rect 204352 474088 204404 474094
rect 204352 474030 204404 474036
rect 204168 379568 204220 379574
rect 204168 379510 204220 379516
rect 204076 378956 204128 378962
rect 204076 378898 204128 378904
rect 204180 376106 204208 379510
rect 204258 379128 204314 379137
rect 204258 379063 204314 379072
rect 204272 378457 204300 379063
rect 204258 378448 204314 378457
rect 204258 378383 204314 378392
rect 204168 376100 204220 376106
rect 204168 376042 204220 376048
rect 203892 282804 203944 282810
rect 203892 282746 203944 282752
rect 203800 272672 203852 272678
rect 203800 272614 203852 272620
rect 203708 271584 203760 271590
rect 203708 271526 203760 271532
rect 204364 269890 204392 474030
rect 204456 411534 204484 491438
rect 204628 471504 204680 471510
rect 204628 471446 204680 471452
rect 204536 466608 204588 466614
rect 204536 466550 204588 466556
rect 204444 411528 204496 411534
rect 204444 411470 204496 411476
rect 204444 410576 204496 410582
rect 204444 410518 204496 410524
rect 204456 376378 204484 410518
rect 204444 376372 204496 376378
rect 204444 376314 204496 376320
rect 204548 359582 204576 466550
rect 204640 380594 204668 471446
rect 204628 380588 204680 380594
rect 204628 380530 204680 380536
rect 204732 380225 204760 493023
rect 204824 493023 205022 493051
rect 204824 491502 204852 493023
rect 204812 491496 204864 491502
rect 204812 491438 204864 491444
rect 205468 483750 205496 493037
rect 205640 491088 205692 491094
rect 205638 491056 205640 491065
rect 205692 491056 205694 491065
rect 205638 490991 205694 491000
rect 205640 490884 205692 490890
rect 205640 490826 205692 490832
rect 205652 490385 205680 490826
rect 205638 490376 205694 490385
rect 205638 490311 205694 490320
rect 205456 483744 205508 483750
rect 205456 483686 205508 483692
rect 204904 480956 204956 480962
rect 204904 480898 204956 480904
rect 204718 380216 204774 380225
rect 204718 380151 204774 380160
rect 204732 379953 204760 380151
rect 204718 379944 204774 379953
rect 204718 379879 204774 379888
rect 204718 378992 204774 379001
rect 204718 378927 204774 378936
rect 204732 378185 204760 378927
rect 204810 378584 204866 378593
rect 204810 378519 204866 378528
rect 204824 378282 204852 378519
rect 204812 378276 204864 378282
rect 204812 378218 204864 378224
rect 204718 378176 204774 378185
rect 204718 378111 204774 378120
rect 204536 359576 204588 359582
rect 204536 359518 204588 359524
rect 204352 269884 204404 269890
rect 204352 269826 204404 269832
rect 203616 166456 203668 166462
rect 203616 166398 203668 166404
rect 203522 165472 203578 165481
rect 203522 165407 203578 165416
rect 204916 165102 204944 480898
rect 204996 478236 205048 478242
rect 204996 478178 205048 478184
rect 205008 175234 205036 478178
rect 205732 474292 205784 474298
rect 205732 474234 205784 474240
rect 205088 472796 205140 472802
rect 205088 472738 205140 472744
rect 205100 271318 205128 472738
rect 205548 465724 205600 465730
rect 205548 465666 205600 465672
rect 205178 464400 205234 464409
rect 205178 464335 205234 464344
rect 205192 272610 205220 464335
rect 205560 378894 205588 465666
rect 205744 380526 205772 474234
rect 205928 472802 205956 493037
rect 206020 493023 206402 493051
rect 205916 472796 205968 472802
rect 205916 472738 205968 472744
rect 205824 471436 205876 471442
rect 205824 471378 205876 471384
rect 205732 380520 205784 380526
rect 205732 380462 205784 380468
rect 205836 380118 205864 471378
rect 206020 413302 206048 493023
rect 206652 491224 206704 491230
rect 206652 491166 206704 491172
rect 206560 490748 206612 490754
rect 206560 490690 206612 490696
rect 206284 472660 206336 472666
rect 206284 472602 206336 472608
rect 206192 414724 206244 414730
rect 206192 414666 206244 414672
rect 206008 413296 206060 413302
rect 206008 413238 206060 413244
rect 205914 380216 205970 380225
rect 205914 380151 205970 380160
rect 205824 380112 205876 380118
rect 205824 380054 205876 380060
rect 205730 379128 205786 379137
rect 205730 379063 205786 379072
rect 205548 378888 205600 378894
rect 205548 378830 205600 378836
rect 205560 378321 205588 378830
rect 205640 378616 205692 378622
rect 205640 378558 205692 378564
rect 205652 378350 205680 378558
rect 205744 378350 205772 379063
rect 205640 378344 205692 378350
rect 205546 378312 205602 378321
rect 205640 378286 205692 378292
rect 205732 378344 205784 378350
rect 205732 378286 205784 378292
rect 205546 378247 205602 378256
rect 205364 378072 205416 378078
rect 205364 378014 205416 378020
rect 205376 377913 205404 378014
rect 205456 378004 205508 378010
rect 205456 377946 205508 377952
rect 205362 377904 205418 377913
rect 205362 377839 205418 377848
rect 205468 377777 205496 377946
rect 205454 377768 205510 377777
rect 205454 377703 205510 377712
rect 205928 376514 205956 380151
rect 206204 378078 206232 414666
rect 206192 378072 206244 378078
rect 206192 378014 206244 378020
rect 205916 376508 205968 376514
rect 205916 376450 205968 376456
rect 205928 373994 205956 376450
rect 206204 374814 206232 378014
rect 206192 374808 206244 374814
rect 206192 374750 206244 374756
rect 205652 373966 205956 373994
rect 205180 272604 205232 272610
rect 205180 272546 205232 272552
rect 205088 271312 205140 271318
rect 205088 271254 205140 271260
rect 205652 269074 205680 373966
rect 205640 269068 205692 269074
rect 205640 269010 205692 269016
rect 205652 267734 205680 269010
rect 205560 267706 205680 267734
rect 204996 175228 205048 175234
rect 204996 175170 205048 175176
rect 204904 165096 204956 165102
rect 204904 165038 204956 165044
rect 201500 165028 201552 165034
rect 201500 164970 201552 164976
rect 205560 161430 205588 267706
rect 206296 164830 206324 472602
rect 206468 469192 206520 469198
rect 206468 469134 206520 469140
rect 206376 466064 206428 466070
rect 206376 466006 206428 466012
rect 206388 166666 206416 466006
rect 206480 271561 206508 469134
rect 206572 378010 206600 490690
rect 206664 378010 206692 491166
rect 206744 465520 206796 465526
rect 206744 465462 206796 465468
rect 206560 378004 206612 378010
rect 206560 377946 206612 377952
rect 206652 378004 206704 378010
rect 206652 377946 206704 377952
rect 206572 374950 206600 377946
rect 206756 376514 206784 465462
rect 206848 416770 206876 493037
rect 207230 493023 207428 493051
rect 207020 491496 207072 491502
rect 207020 491438 207072 491444
rect 206836 416764 206888 416770
rect 206836 416706 206888 416712
rect 206836 411528 206888 411534
rect 206836 411470 206888 411476
rect 206848 409154 206876 411470
rect 206836 409148 206888 409154
rect 206836 409090 206888 409096
rect 207032 380769 207060 491438
rect 207296 474156 207348 474162
rect 207296 474098 207348 474104
rect 207112 465792 207164 465798
rect 207112 465734 207164 465740
rect 207018 380760 207074 380769
rect 207018 380695 207074 380704
rect 207032 380361 207060 380695
rect 207018 380352 207074 380361
rect 207018 380287 207074 380296
rect 207124 380050 207152 465734
rect 207204 416764 207256 416770
rect 207204 416706 207256 416712
rect 207216 414866 207244 416706
rect 207204 414860 207256 414866
rect 207204 414802 207256 414808
rect 207112 380044 207164 380050
rect 207112 379986 207164 379992
rect 207018 379128 207074 379137
rect 207018 379063 207074 379072
rect 206836 378616 206888 378622
rect 206836 378558 206888 378564
rect 206744 376508 206796 376514
rect 206744 376450 206796 376456
rect 206560 374944 206612 374950
rect 206560 374886 206612 374892
rect 206466 271552 206522 271561
rect 206466 271487 206522 271496
rect 206848 269822 206876 378558
rect 207032 378418 207060 379063
rect 207020 378412 207072 378418
rect 207020 378354 207072 378360
rect 206928 378344 206980 378350
rect 206928 378286 206980 378292
rect 206836 269816 206888 269822
rect 206836 269758 206888 269764
rect 206940 269686 206968 378286
rect 207308 377330 207336 474098
rect 207400 464506 207428 493023
rect 207492 493023 207690 493051
rect 207768 493023 208150 493051
rect 207388 464500 207440 464506
rect 207388 464442 207440 464448
rect 207492 464370 207520 493023
rect 207768 491502 207796 493023
rect 207756 491496 207808 491502
rect 207756 491438 207808 491444
rect 207940 490884 207992 490890
rect 207940 490826 207992 490832
rect 207756 472864 207808 472870
rect 207756 472806 207808 472812
rect 207664 469872 207716 469878
rect 207664 469814 207716 469820
rect 207480 464364 207532 464370
rect 207480 464306 207532 464312
rect 207572 378412 207624 378418
rect 207572 378354 207624 378360
rect 207296 377324 207348 377330
rect 207296 377266 207348 377272
rect 207296 376440 207348 376446
rect 207296 376382 207348 376388
rect 207308 374649 207336 376382
rect 207294 374640 207350 374649
rect 207294 374575 207350 374584
rect 206928 269680 206980 269686
rect 206928 269622 206980 269628
rect 207584 268394 207612 378354
rect 207572 268388 207624 268394
rect 207572 268330 207624 268336
rect 206376 166660 206428 166666
rect 206376 166602 206428 166608
rect 207676 164898 207704 469814
rect 207768 271017 207796 472806
rect 207848 466336 207900 466342
rect 207848 466278 207900 466284
rect 207860 273290 207888 466278
rect 207952 376446 207980 490826
rect 208400 490680 208452 490686
rect 208400 490622 208452 490628
rect 208412 490385 208440 490622
rect 208398 490376 208454 490385
rect 208398 490311 208454 490320
rect 208596 489938 208624 493037
rect 208688 493023 209070 493051
rect 208584 489932 208636 489938
rect 208584 489874 208636 489880
rect 208032 467492 208084 467498
rect 208032 467434 208084 467440
rect 207940 376440 207992 376446
rect 207940 376382 207992 376388
rect 208044 375970 208072 467434
rect 208216 464500 208268 464506
rect 208216 464442 208268 464448
rect 208124 464364 208176 464370
rect 208124 464306 208176 464312
rect 208136 417450 208164 464306
rect 208228 418810 208256 464442
rect 208216 418804 208268 418810
rect 208216 418746 208268 418752
rect 208216 418056 208268 418062
rect 208216 417998 208268 418004
rect 208124 417444 208176 417450
rect 208124 417386 208176 417392
rect 208228 391950 208256 417998
rect 208688 402974 208716 493023
rect 209044 490816 209096 490822
rect 209044 490758 209096 490764
rect 208952 464772 209004 464778
rect 208952 464714 209004 464720
rect 208688 402946 208808 402974
rect 208492 400240 208544 400246
rect 208492 400182 208544 400188
rect 208216 391944 208268 391950
rect 208216 391886 208268 391892
rect 208306 379944 208362 379953
rect 208306 379879 208308 379888
rect 208360 379879 208362 379888
rect 208308 379850 208360 379856
rect 208122 378448 208178 378457
rect 208122 378383 208178 378392
rect 208032 375964 208084 375970
rect 208032 375906 208084 375912
rect 207848 273284 207900 273290
rect 207848 273226 207900 273232
rect 207754 271008 207810 271017
rect 207754 270943 207810 270952
rect 208136 270337 208164 378383
rect 208122 270328 208178 270337
rect 208122 270263 208178 270272
rect 207664 164892 207716 164898
rect 207664 164834 207716 164840
rect 206284 164824 206336 164830
rect 206284 164766 206336 164772
rect 205548 161424 205600 161430
rect 205548 161366 205600 161372
rect 208136 147626 208164 270263
rect 208320 268462 208348 379850
rect 208504 371210 208532 400182
rect 208780 379370 208808 402946
rect 208768 379364 208820 379370
rect 208768 379306 208820 379312
rect 208780 378486 208808 379306
rect 208768 378480 208820 378486
rect 208768 378422 208820 378428
rect 208964 376378 208992 464714
rect 208952 376372 209004 376378
rect 208952 376314 209004 376320
rect 208492 371204 208544 371210
rect 208492 371146 208544 371152
rect 208308 268456 208360 268462
rect 208308 268398 208360 268404
rect 208124 147620 208176 147626
rect 208124 147562 208176 147568
rect 209056 58954 209084 490758
rect 209424 490686 209452 493037
rect 209780 491496 209832 491502
rect 209780 491438 209832 491444
rect 209412 490680 209464 490686
rect 209412 490622 209464 490628
rect 209136 488300 209188 488306
rect 209136 488242 209188 488248
rect 209148 164762 209176 488242
rect 209504 479664 209556 479670
rect 209504 479606 209556 479612
rect 209226 471200 209282 471209
rect 209226 471135 209282 471144
rect 209240 166802 209268 471135
rect 209412 470008 209464 470014
rect 209412 469950 209464 469956
rect 209320 468852 209372 468858
rect 209320 468794 209372 468800
rect 209228 166796 209280 166802
rect 209228 166738 209280 166744
rect 209332 166598 209360 468794
rect 209424 178022 209452 469950
rect 209516 271182 209544 479606
rect 209792 468314 209820 491438
rect 209780 468308 209832 468314
rect 209780 468250 209832 468256
rect 209596 467356 209648 467362
rect 209596 467298 209648 467304
rect 209608 272746 209636 467298
rect 209884 379001 209912 493037
rect 210056 490680 210108 490686
rect 210056 490622 210108 490628
rect 210068 379438 210096 490622
rect 210240 471232 210292 471238
rect 210240 471174 210292 471180
rect 210056 379432 210108 379438
rect 210056 379374 210108 379380
rect 209870 378992 209926 379001
rect 209870 378927 209926 378936
rect 209686 378584 209742 378593
rect 209686 378519 209742 378528
rect 209596 272740 209648 272746
rect 209596 272682 209648 272688
rect 209504 271176 209556 271182
rect 209504 271118 209556 271124
rect 209412 178016 209464 178022
rect 209412 177958 209464 177964
rect 209320 166592 209372 166598
rect 209320 166534 209372 166540
rect 209136 164756 209188 164762
rect 209136 164698 209188 164704
rect 209044 58948 209096 58954
rect 209044 58890 209096 58896
rect 201408 58880 201460 58886
rect 201408 58822 201460 58828
rect 209700 57866 209728 378519
rect 210252 376174 210280 471174
rect 210344 379302 210372 493037
rect 210528 493023 210818 493051
rect 210528 491502 210556 493023
rect 210516 491496 210568 491502
rect 210516 491438 210568 491444
rect 210516 489252 210568 489258
rect 210516 489194 210568 489200
rect 210424 466472 210476 466478
rect 210424 466414 210476 466420
rect 210436 389366 210464 466414
rect 210424 389360 210476 389366
rect 210424 389302 210476 389308
rect 210332 379296 210384 379302
rect 210332 379238 210384 379244
rect 210330 378856 210386 378865
rect 210330 378791 210386 378800
rect 210344 378418 210372 378791
rect 210332 378412 210384 378418
rect 210332 378354 210384 378360
rect 210240 376168 210292 376174
rect 210240 376110 210292 376116
rect 210344 270502 210372 378354
rect 210436 360874 210464 389302
rect 210424 360868 210476 360874
rect 210424 360810 210476 360816
rect 210332 270496 210384 270502
rect 210332 270438 210384 270444
rect 210528 165510 210556 489194
rect 210608 476876 210660 476882
rect 210608 476818 210660 476824
rect 210516 165504 210568 165510
rect 210516 165446 210568 165452
rect 210620 164966 210648 476818
rect 210700 472728 210752 472734
rect 210700 472670 210752 472676
rect 210712 271250 210740 472670
rect 210792 470076 210844 470082
rect 210792 470018 210844 470024
rect 210700 271244 210752 271250
rect 210700 271186 210752 271192
rect 210804 271046 210832 470018
rect 210884 464568 210936 464574
rect 210884 464510 210936 464516
rect 210896 272882 210924 464510
rect 211066 379536 211122 379545
rect 211066 379471 211122 379480
rect 210976 379296 211028 379302
rect 210976 379238 211028 379244
rect 210988 378690 211016 379238
rect 210976 378684 211028 378690
rect 210976 378626 211028 378632
rect 210976 378276 211028 378282
rect 210976 378218 211028 378224
rect 210988 378185 211016 378218
rect 210974 378176 211030 378185
rect 210974 378111 211030 378120
rect 210976 378072 211028 378078
rect 210976 378014 211028 378020
rect 210884 272876 210936 272882
rect 210884 272818 210936 272824
rect 210792 271040 210844 271046
rect 210792 270982 210844 270988
rect 210884 270496 210936 270502
rect 210884 270438 210936 270444
rect 210896 270162 210924 270438
rect 210988 270366 211016 378014
rect 210976 270360 211028 270366
rect 210976 270302 211028 270308
rect 210884 270156 210936 270162
rect 210884 270098 210936 270104
rect 210792 269680 210844 269686
rect 210792 269622 210844 269628
rect 210608 164960 210660 164966
rect 210608 164902 210660 164908
rect 210804 144906 210832 269622
rect 210896 148510 210924 270098
rect 210884 148504 210936 148510
rect 210884 148446 210936 148452
rect 210792 144900 210844 144906
rect 210792 144842 210844 144848
rect 197452 57860 197504 57866
rect 197452 57802 197504 57808
rect 209688 57860 209740 57866
rect 209688 57802 209740 57808
rect 183192 57792 183244 57798
rect 183190 57760 183192 57769
rect 197360 57792 197412 57798
rect 183244 57760 183246 57769
rect 197360 57734 197412 57740
rect 183190 57695 183246 57704
rect 155958 57624 156014 57633
rect 155958 57559 156014 57568
rect 160098 57624 160154 57633
rect 160098 57559 160154 57568
rect 165618 57624 165674 57633
rect 165618 57559 165674 57568
rect 153290 56264 153346 56273
rect 153290 56199 153346 56208
rect 155972 54913 156000 57559
rect 160112 55049 160140 57559
rect 165632 55185 165660 57559
rect 211080 57526 211108 379471
rect 211172 379166 211200 493037
rect 211632 491230 211660 493037
rect 211620 491224 211672 491230
rect 211620 491166 211672 491172
rect 212092 491065 212120 493037
rect 212566 493023 212672 493051
rect 212540 491292 212592 491298
rect 212540 491234 212592 491240
rect 212078 491056 212134 491065
rect 212078 490991 212134 491000
rect 212552 490657 212580 491234
rect 212538 490648 212594 490657
rect 212538 490583 212594 490592
rect 212264 490340 212316 490346
rect 212264 490282 212316 490288
rect 211252 489932 211304 489938
rect 211252 489874 211304 489880
rect 211264 380769 211292 489874
rect 211804 486532 211856 486538
rect 211804 486474 211856 486480
rect 211620 464704 211672 464710
rect 211620 464646 211672 464652
rect 211250 380760 211306 380769
rect 211250 380695 211306 380704
rect 211528 379432 211580 379438
rect 211528 379374 211580 379380
rect 211160 379160 211212 379166
rect 211160 379102 211212 379108
rect 211540 378758 211568 379374
rect 211528 378752 211580 378758
rect 211528 378694 211580 378700
rect 211540 270502 211568 378694
rect 211632 376242 211660 464646
rect 211712 378956 211764 378962
rect 211712 378898 211764 378904
rect 211724 378214 211752 378898
rect 211712 378208 211764 378214
rect 211712 378150 211764 378156
rect 211620 376236 211672 376242
rect 211620 376178 211672 376184
rect 211724 273426 211752 378150
rect 211712 273420 211764 273426
rect 211712 273362 211764 273368
rect 211528 270496 211580 270502
rect 211528 270438 211580 270444
rect 211724 146169 211752 273362
rect 211816 165306 211844 486474
rect 211896 475516 211948 475522
rect 211896 475458 211948 475464
rect 211908 165578 211936 475458
rect 212080 471776 212132 471782
rect 212080 471718 212132 471724
rect 211988 468784 212040 468790
rect 211988 468726 212040 468732
rect 212000 166530 212028 468726
rect 212092 273494 212120 471718
rect 212172 467424 212224 467430
rect 212172 467366 212224 467372
rect 212080 273488 212132 273494
rect 212080 273430 212132 273436
rect 212184 271862 212212 467366
rect 212276 378078 212304 490282
rect 212448 465792 212500 465798
rect 212448 465734 212500 465740
rect 212356 378480 212408 378486
rect 212356 378422 212408 378428
rect 212264 378072 212316 378078
rect 212264 378014 212316 378020
rect 212172 271856 212224 271862
rect 212172 271798 212224 271804
rect 212368 270434 212396 378422
rect 212460 378185 212488 465734
rect 212644 380633 212672 493023
rect 212908 466404 212960 466410
rect 212908 466346 212960 466352
rect 212630 380624 212686 380633
rect 212630 380559 212686 380568
rect 212644 379778 212672 380559
rect 212632 379772 212684 379778
rect 212632 379714 212684 379720
rect 212446 378176 212502 378185
rect 212446 378111 212502 378120
rect 212446 378040 212502 378049
rect 212446 377975 212502 377984
rect 212356 270428 212408 270434
rect 212356 270370 212408 270376
rect 212172 268388 212224 268394
rect 212172 268330 212224 268336
rect 211988 166524 212040 166530
rect 211988 166466 212040 166472
rect 211896 165572 211948 165578
rect 211896 165514 211948 165520
rect 211804 165300 211856 165306
rect 211804 165242 211856 165248
rect 212184 148986 212212 268330
rect 212368 258074 212396 270370
rect 212276 258046 212396 258074
rect 212172 148980 212224 148986
rect 212172 148922 212224 148928
rect 211710 146160 211766 146169
rect 211710 146095 211766 146104
rect 211802 145888 211858 145897
rect 211802 145823 211858 145832
rect 211816 144906 211844 145823
rect 211804 144900 211856 144906
rect 211804 144842 211856 144848
rect 211068 57520 211120 57526
rect 211068 57462 211120 57468
rect 211816 55894 211844 144842
rect 211804 55888 211856 55894
rect 211804 55830 211856 55836
rect 212184 55185 212212 148922
rect 212276 144770 212304 258046
rect 212264 144764 212316 144770
rect 212264 144706 212316 144712
rect 212460 57730 212488 377975
rect 212920 376446 212948 466346
rect 213012 380497 213040 493037
rect 213380 491201 213408 493037
rect 213840 491298 213868 493037
rect 214012 491564 214064 491570
rect 214012 491506 214064 491512
rect 213920 491496 213972 491502
rect 213920 491438 213972 491444
rect 213828 491292 213880 491298
rect 213828 491234 213880 491240
rect 213366 491192 213422 491201
rect 213366 491127 213422 491136
rect 213276 486464 213328 486470
rect 213276 486406 213328 486412
rect 213184 475448 213236 475454
rect 213184 475390 213236 475396
rect 213092 468444 213144 468450
rect 213092 468386 213144 468392
rect 212998 380488 213054 380497
rect 212998 380423 213054 380432
rect 213012 379817 213040 380423
rect 212998 379808 213054 379817
rect 212998 379743 213054 379752
rect 212998 379400 213054 379409
rect 212998 379335 213054 379344
rect 213012 379001 213040 379335
rect 212998 378992 213054 379001
rect 212998 378927 213054 378936
rect 213000 378548 213052 378554
rect 213000 378490 213052 378496
rect 212908 376440 212960 376446
rect 212908 376382 212960 376388
rect 213012 277394 213040 378490
rect 213104 377330 213132 468386
rect 213092 377324 213144 377330
rect 213092 377266 213144 377272
rect 213092 376032 213144 376038
rect 213092 375974 213144 375980
rect 212828 277366 213040 277394
rect 212828 273358 212856 277366
rect 212816 273352 212868 273358
rect 212816 273294 212868 273300
rect 212828 149054 212856 273294
rect 212906 270192 212962 270201
rect 212906 270127 212962 270136
rect 212816 149048 212868 149054
rect 212816 148990 212868 148996
rect 212828 147694 212856 148990
rect 212920 148578 212948 270127
rect 213000 269816 213052 269822
rect 213000 269758 213052 269764
rect 212908 148572 212960 148578
rect 212908 148514 212960 148520
rect 212816 147688 212868 147694
rect 212816 147630 212868 147636
rect 213012 144838 213040 269758
rect 213104 268666 213132 375974
rect 213092 268660 213144 268666
rect 213092 268602 213144 268608
rect 213092 148368 213144 148374
rect 213092 148310 213144 148316
rect 213000 144832 213052 144838
rect 213000 144774 213052 144780
rect 212448 57724 212500 57730
rect 212448 57666 212500 57672
rect 213104 56574 213132 148310
rect 213196 57458 213224 475390
rect 213288 68950 213316 486406
rect 213368 479596 213420 479602
rect 213368 479538 213420 479544
rect 213380 165374 213408 479538
rect 213552 474224 213604 474230
rect 213552 474166 213604 474172
rect 213460 468716 213512 468722
rect 213460 468658 213512 468664
rect 213472 166394 213500 468658
rect 213564 271425 213592 474166
rect 213828 466404 213880 466410
rect 213828 466346 213880 466352
rect 213642 380760 213698 380769
rect 213642 380695 213698 380704
rect 213656 379846 213684 380695
rect 213736 380044 213788 380050
rect 213736 379986 213788 379992
rect 213644 379840 213696 379846
rect 213644 379782 213696 379788
rect 213748 379574 213776 379986
rect 213736 379568 213788 379574
rect 213656 379516 213736 379522
rect 213656 379510 213788 379516
rect 213656 379494 213776 379510
rect 213656 271930 213684 379494
rect 213736 379432 213788 379438
rect 213736 379374 213788 379380
rect 213748 378554 213776 379374
rect 213840 379273 213868 466346
rect 213826 379264 213882 379273
rect 213826 379199 213882 379208
rect 213840 379001 213868 379199
rect 213826 378992 213882 379001
rect 213826 378927 213882 378936
rect 213828 378888 213880 378894
rect 213828 378830 213880 378836
rect 213736 378548 213788 378554
rect 213736 378490 213788 378496
rect 213840 378434 213868 378830
rect 213748 378406 213868 378434
rect 213644 271924 213696 271930
rect 213644 271866 213696 271872
rect 213550 271416 213606 271425
rect 213550 271351 213606 271360
rect 213748 268870 213776 378406
rect 213826 378040 213882 378049
rect 213826 377975 213882 377984
rect 213736 268864 213788 268870
rect 213736 268806 213788 268812
rect 213748 258074 213776 268806
rect 213564 258046 213776 258074
rect 213460 166388 213512 166394
rect 213460 166330 213512 166336
rect 213368 165368 213420 165374
rect 213368 165310 213420 165316
rect 213460 148504 213512 148510
rect 213460 148446 213512 148452
rect 213368 147620 213420 147626
rect 213368 147562 213420 147568
rect 213276 68944 213328 68950
rect 213276 68886 213328 68892
rect 213184 57452 213236 57458
rect 213184 57394 213236 57400
rect 213092 56568 213144 56574
rect 213092 56510 213144 56516
rect 165618 55176 165674 55185
rect 165618 55111 165674 55120
rect 212170 55176 212226 55185
rect 212170 55111 212226 55120
rect 160098 55040 160154 55049
rect 160098 54975 160154 54984
rect 155958 54904 156014 54913
rect 155958 54839 156014 54848
rect 86960 54742 87012 54748
rect 118698 54768 118754 54777
rect 81440 54732 81492 54738
rect 118698 54703 118754 54712
rect 81440 54674 81492 54680
rect 213380 54670 213408 147562
rect 78680 54664 78732 54670
rect 78680 54606 78732 54612
rect 213368 54664 213420 54670
rect 213368 54606 213420 54612
rect 213472 54398 213500 148446
rect 213564 144906 213592 258046
rect 213644 148912 213696 148918
rect 213644 148854 213696 148860
rect 213656 148578 213684 148854
rect 213644 148572 213696 148578
rect 213644 148514 213696 148520
rect 213552 144900 213604 144906
rect 213552 144842 213604 144848
rect 213656 55826 213684 148514
rect 213736 148436 213788 148442
rect 213736 148378 213788 148384
rect 213748 147626 213776 148378
rect 213736 147620 213788 147626
rect 213736 147562 213788 147568
rect 213736 147484 213788 147490
rect 213736 147426 213788 147432
rect 213748 56438 213776 147426
rect 213840 59090 213868 377975
rect 213932 375358 213960 491438
rect 214024 376582 214052 491506
rect 214300 383654 214328 493037
rect 214392 493023 214774 493051
rect 214944 493023 215234 493051
rect 214392 491502 214420 493023
rect 214944 491570 214972 493023
rect 214932 491564 214984 491570
rect 214932 491506 214984 491512
rect 214380 491496 214432 491502
rect 214380 491438 214432 491444
rect 215300 491496 215352 491502
rect 215300 491438 215352 491444
rect 214564 485104 214616 485110
rect 214564 485046 214616 485052
rect 214472 464636 214524 464642
rect 214472 464578 214524 464584
rect 214300 383626 214420 383654
rect 214392 380089 214420 383626
rect 214378 380080 214434 380089
rect 214378 380015 214434 380024
rect 214104 379840 214156 379846
rect 214104 379782 214156 379788
rect 214116 378894 214144 379782
rect 214104 378888 214156 378894
rect 214104 378830 214156 378836
rect 214392 376650 214420 380015
rect 214380 376644 214432 376650
rect 214380 376586 214432 376592
rect 214012 376576 214064 376582
rect 214012 376518 214064 376524
rect 214024 375834 214052 376518
rect 214012 375828 214064 375834
rect 214012 375770 214064 375776
rect 213920 375352 213972 375358
rect 213920 375294 213972 375300
rect 213932 374338 213960 375294
rect 213920 374332 213972 374338
rect 213920 374274 213972 374280
rect 214102 271824 214158 271833
rect 214102 271759 214158 271768
rect 213828 59084 213880 59090
rect 213828 59026 213880 59032
rect 214116 57186 214144 271759
rect 214288 269952 214340 269958
rect 214288 269894 214340 269900
rect 214300 164218 214328 269894
rect 214392 268598 214420 376586
rect 214484 376582 214512 464578
rect 214472 376576 214524 376582
rect 214472 376518 214524 376524
rect 214472 357672 214524 357678
rect 214472 357614 214524 357620
rect 214484 270201 214512 357614
rect 214470 270192 214526 270201
rect 214470 270127 214526 270136
rect 214472 268728 214524 268734
rect 214472 268670 214524 268676
rect 214380 268592 214432 268598
rect 214380 268534 214432 268540
rect 214484 268462 214512 268670
rect 214472 268456 214524 268462
rect 214472 268398 214524 268404
rect 214288 164212 214340 164218
rect 214288 164154 214340 164160
rect 214484 151814 214512 268398
rect 214576 164694 214604 485046
rect 214840 483676 214892 483682
rect 214840 483618 214892 483624
rect 214748 467220 214800 467226
rect 214748 467162 214800 467168
rect 214656 465928 214708 465934
rect 214656 465870 214708 465876
rect 214668 165238 214696 465870
rect 214760 166326 214788 467162
rect 214852 271386 214880 483618
rect 214932 471980 214984 471986
rect 214932 471922 214984 471928
rect 214944 376310 214972 471922
rect 215208 469940 215260 469946
rect 215208 469882 215260 469888
rect 215114 376680 215170 376689
rect 215114 376615 215170 376624
rect 215022 376544 215078 376553
rect 215022 376479 215078 376488
rect 214932 376304 214984 376310
rect 214932 376246 214984 376252
rect 214932 375352 214984 375358
rect 214932 375294 214984 375300
rect 214944 374746 214972 375294
rect 214932 374740 214984 374746
rect 214932 374682 214984 374688
rect 214840 271380 214892 271386
rect 214840 271322 214892 271328
rect 214840 270360 214892 270366
rect 214840 270302 214892 270308
rect 214852 269890 214880 270302
rect 214944 269958 214972 374682
rect 214932 269952 214984 269958
rect 214932 269894 214984 269900
rect 214840 269884 214892 269890
rect 214840 269826 214892 269832
rect 214748 166320 214800 166326
rect 214748 166262 214800 166268
rect 214656 165232 214708 165238
rect 214656 165174 214708 165180
rect 214564 164688 214616 164694
rect 214564 164630 214616 164636
rect 214656 162580 214708 162586
rect 214656 162522 214708 162528
rect 214300 151786 214512 151814
rect 214194 146296 214250 146305
rect 214194 146231 214250 146240
rect 214104 57180 214156 57186
rect 214104 57122 214156 57128
rect 213736 56432 213788 56438
rect 213736 56374 213788 56380
rect 213644 55820 213696 55826
rect 213644 55762 213696 55768
rect 214208 54466 214236 146231
rect 214300 145518 214328 151786
rect 214380 145852 214432 145858
rect 214380 145794 214432 145800
rect 214288 145512 214340 145518
rect 214288 145454 214340 145460
rect 214300 55146 214328 145454
rect 214392 56030 214420 145794
rect 214564 145580 214616 145586
rect 214564 145522 214616 145528
rect 214576 69018 214604 145522
rect 214564 69012 214616 69018
rect 214564 68954 214616 68960
rect 214668 59498 214696 162522
rect 214748 161900 214800 161906
rect 214748 161842 214800 161848
rect 214760 62014 214788 161842
rect 214852 146305 214880 269826
rect 214944 269550 214972 269894
rect 214932 269544 214984 269550
rect 214932 269486 214984 269492
rect 214838 146296 214894 146305
rect 214838 146231 214894 146240
rect 214838 146160 214894 146169
rect 214838 146095 214894 146104
rect 214852 145625 214880 146095
rect 214838 145616 214894 145625
rect 214838 145551 214894 145560
rect 214748 62008 214800 62014
rect 214748 61950 214800 61956
rect 214656 59492 214708 59498
rect 214656 59434 214708 59440
rect 214748 59356 214800 59362
rect 214748 59298 214800 59304
rect 214760 57934 214788 59298
rect 214748 57928 214800 57934
rect 214748 57870 214800 57876
rect 214380 56024 214432 56030
rect 214380 55966 214432 55972
rect 214288 55140 214340 55146
rect 214288 55082 214340 55088
rect 214852 54534 214880 145551
rect 214932 62008 214984 62014
rect 214932 61950 214984 61956
rect 214944 59158 214972 61950
rect 214932 59152 214984 59158
rect 214932 59094 214984 59100
rect 215036 57798 215064 376479
rect 215024 57792 215076 57798
rect 215024 57734 215076 57740
rect 215128 57390 215156 376615
rect 215220 270910 215248 469882
rect 215312 383654 215340 491438
rect 215312 383626 215432 383654
rect 215298 380352 215354 380361
rect 215298 380287 215354 380296
rect 215312 379982 215340 380287
rect 215300 379976 215352 379982
rect 215300 379918 215352 379924
rect 215404 377913 215432 383626
rect 215390 377904 215446 377913
rect 215390 377839 215446 377848
rect 215588 375358 215616 493037
rect 215944 489184 215996 489190
rect 215944 489126 215996 489132
rect 215852 471912 215904 471918
rect 215852 471854 215904 471860
rect 215668 379704 215720 379710
rect 215668 379646 215720 379652
rect 215680 377262 215708 379646
rect 215668 377256 215720 377262
rect 215668 377198 215720 377204
rect 215864 375766 215892 471854
rect 215852 375760 215904 375766
rect 215852 375702 215904 375708
rect 215576 375352 215628 375358
rect 215576 375294 215628 375300
rect 215852 374876 215904 374882
rect 215852 374818 215904 374824
rect 215864 374338 215892 374818
rect 215852 374332 215904 374338
rect 215852 374274 215904 374280
rect 215668 271924 215720 271930
rect 215668 271866 215720 271872
rect 215208 270904 215260 270910
rect 215208 270846 215260 270852
rect 215208 270088 215260 270094
rect 215208 270030 215260 270036
rect 215220 145858 215248 270030
rect 215208 145852 215260 145858
rect 215208 145794 215260 145800
rect 215220 145382 215248 145794
rect 215680 145450 215708 271866
rect 215864 268530 215892 374274
rect 215852 268524 215904 268530
rect 215852 268466 215904 268472
rect 215956 165034 215984 489126
rect 216048 379710 216076 493037
rect 216232 493023 216522 493051
rect 216232 491502 216260 493023
rect 216220 491496 216272 491502
rect 216220 491438 216272 491444
rect 216128 471844 216180 471850
rect 216128 471786 216180 471792
rect 216036 379704 216088 379710
rect 216036 379646 216088 379652
rect 216036 374808 216088 374814
rect 216036 374750 216088 374756
rect 216048 251870 216076 374750
rect 216140 272814 216168 471786
rect 216772 471708 216824 471714
rect 216772 471650 216824 471656
rect 216220 467288 216272 467294
rect 216220 467230 216272 467236
rect 216128 272808 216180 272814
rect 216128 272750 216180 272756
rect 216232 271697 216260 467230
rect 216312 466132 216364 466138
rect 216312 466074 216364 466080
rect 216218 271688 216274 271697
rect 216218 271623 216274 271632
rect 216324 271522 216352 466074
rect 216784 422294 216812 471650
rect 216692 422266 216812 422294
rect 216692 415290 216720 422266
rect 216864 418804 216916 418810
rect 216864 418746 216916 418752
rect 216770 417888 216826 417897
rect 216770 417823 216826 417832
rect 216784 417450 216812 417823
rect 216772 417444 216824 417450
rect 216772 417386 216824 417392
rect 216876 416945 216904 418746
rect 216862 416936 216918 416945
rect 216862 416871 216918 416880
rect 216508 415262 216720 415290
rect 216404 379976 216456 379982
rect 216404 379918 216456 379924
rect 216312 271516 216364 271522
rect 216312 271458 216364 271464
rect 216416 268802 216444 379918
rect 216508 271454 216536 415262
rect 216864 414860 216916 414866
rect 216864 414802 216916 414808
rect 216876 414769 216904 414802
rect 216862 414760 216918 414769
rect 216968 414730 216996 493037
rect 217428 490890 217456 493037
rect 217416 490884 217468 490890
rect 217416 490826 217468 490832
rect 217796 490754 217824 493037
rect 218152 491224 218204 491230
rect 218152 491166 218204 491172
rect 217784 490748 217836 490754
rect 217784 490690 217836 490696
rect 217416 490612 217468 490618
rect 217416 490554 217468 490560
rect 217324 483744 217376 483750
rect 217324 483686 217376 483692
rect 216862 414695 216918 414704
rect 216956 414724 217008 414730
rect 216678 413808 216734 413817
rect 216678 413743 216734 413752
rect 216692 413302 216720 413743
rect 216680 413296 216732 413302
rect 216680 413238 216732 413244
rect 216692 407658 216720 413238
rect 216770 409184 216826 409193
rect 216770 409119 216772 409128
rect 216824 409119 216826 409128
rect 216772 409090 216824 409096
rect 216680 407652 216732 407658
rect 216680 407594 216732 407600
rect 216876 407538 216904 414695
rect 216956 414666 217008 414672
rect 217336 412634 217364 483686
rect 217244 412606 217364 412634
rect 217244 410961 217272 412606
rect 217230 410952 217286 410961
rect 217230 410887 217286 410896
rect 216956 409148 217008 409154
rect 216956 409090 217008 409096
rect 216692 407510 216904 407538
rect 216692 389450 216720 407510
rect 216772 407448 216824 407454
rect 216772 407390 216824 407396
rect 216600 389422 216720 389450
rect 216600 389178 216628 389422
rect 216680 389360 216732 389366
rect 216678 389328 216680 389337
rect 216732 389328 216734 389337
rect 216678 389263 216734 389272
rect 216600 389150 216720 389178
rect 216692 380798 216720 389150
rect 216784 380866 216812 407390
rect 216968 393314 216996 409090
rect 216876 393286 216996 393314
rect 216772 380860 216824 380866
rect 216772 380802 216824 380808
rect 216680 380792 216732 380798
rect 216680 380734 216732 380740
rect 216692 379642 216720 380734
rect 216680 379636 216732 379642
rect 216680 379578 216732 379584
rect 216586 378040 216642 378049
rect 216586 377975 216642 377984
rect 216496 271448 216548 271454
rect 216496 271390 216548 271396
rect 216496 269204 216548 269210
rect 216496 269146 216548 269152
rect 216404 268796 216456 268802
rect 216404 268738 216456 268744
rect 216416 258074 216444 268738
rect 216324 258046 216444 258074
rect 216128 252068 216180 252074
rect 216128 252010 216180 252016
rect 216036 251864 216088 251870
rect 216036 251806 216088 251812
rect 215944 165028 215996 165034
rect 215944 164970 215996 164976
rect 215760 164212 215812 164218
rect 215760 164154 215812 164160
rect 215772 163674 215800 164154
rect 215760 163668 215812 163674
rect 215760 163610 215812 163616
rect 215668 145444 215720 145450
rect 215668 145386 215720 145392
rect 215208 145376 215260 145382
rect 215208 145318 215260 145324
rect 215680 143750 215708 145386
rect 215668 143744 215720 143750
rect 215668 143686 215720 143692
rect 215208 69012 215260 69018
rect 215208 68954 215260 68960
rect 215220 68406 215248 68954
rect 215208 68400 215260 68406
rect 215208 68342 215260 68348
rect 215220 59362 215248 68342
rect 215772 59430 215800 163610
rect 216140 162790 216168 252010
rect 216220 252000 216272 252006
rect 216220 251942 216272 251948
rect 216128 162784 216180 162790
rect 216128 162726 216180 162732
rect 215852 146328 215904 146334
rect 215852 146270 215904 146276
rect 215864 96626 215892 146270
rect 215944 144832 215996 144838
rect 215944 144774 215996 144780
rect 215852 96620 215904 96626
rect 215852 96562 215904 96568
rect 215760 59424 215812 59430
rect 215760 59366 215812 59372
rect 215208 59356 215260 59362
rect 215208 59298 215260 59304
rect 215116 57384 215168 57390
rect 215116 57326 215168 57332
rect 215956 56370 215984 144774
rect 216036 144764 216088 144770
rect 216036 144706 216088 144712
rect 215944 56364 215996 56370
rect 215944 56306 215996 56312
rect 216048 55962 216076 144706
rect 216140 59566 216168 162726
rect 216232 162586 216260 251942
rect 216220 162580 216272 162586
rect 216220 162522 216272 162528
rect 216324 147674 216352 258046
rect 216232 147646 216352 147674
rect 216232 145722 216260 147646
rect 216508 146062 216536 269146
rect 216496 146056 216548 146062
rect 216496 145998 216548 146004
rect 216508 145840 216536 145998
rect 216324 145812 216536 145840
rect 216220 145716 216272 145722
rect 216220 145658 216272 145664
rect 216232 138014 216260 145658
rect 216324 144650 216352 145812
rect 216402 145752 216458 145761
rect 216402 145687 216458 145696
rect 216416 144838 216444 145687
rect 216496 145580 216548 145586
rect 216496 145522 216548 145528
rect 216404 144832 216456 144838
rect 216404 144774 216456 144780
rect 216508 144770 216536 145522
rect 216496 144764 216548 144770
rect 216496 144706 216548 144712
rect 216324 144622 216444 144650
rect 216232 137986 216352 138014
rect 216128 59560 216180 59566
rect 216128 59502 216180 59508
rect 216036 55956 216088 55962
rect 216036 55898 216088 55904
rect 216324 54602 216352 137986
rect 216416 54874 216444 144622
rect 216496 143744 216548 143750
rect 216496 143686 216548 143692
rect 216404 54868 216456 54874
rect 216404 54810 216456 54816
rect 216312 54596 216364 54602
rect 216312 54538 216364 54544
rect 214840 54528 214892 54534
rect 214840 54470 214892 54476
rect 214196 54460 214248 54466
rect 214196 54402 214248 54408
rect 213460 54392 213512 54398
rect 213460 54334 213512 54340
rect 216508 54330 216536 143686
rect 216600 57594 216628 377975
rect 216680 375284 216732 375290
rect 216680 375226 216732 375232
rect 216692 374649 216720 375226
rect 216678 374640 216734 374649
rect 216678 374575 216734 374584
rect 216784 373994 216812 380802
rect 216876 380662 216904 393286
rect 216956 391944 217008 391950
rect 216956 391886 217008 391892
rect 216968 390969 216996 391886
rect 216954 390960 217010 390969
rect 216954 390895 217010 390904
rect 216956 389156 217008 389162
rect 216956 389098 217008 389104
rect 216968 389065 216996 389098
rect 216954 389056 217010 389065
rect 216954 388991 217010 389000
rect 217244 383654 217272 410887
rect 217152 383626 217272 383654
rect 217152 380730 217180 383626
rect 217140 380724 217192 380730
rect 217140 380666 217192 380672
rect 216864 380656 216916 380662
rect 216864 380598 216916 380604
rect 216876 379574 216904 380598
rect 216864 379568 216916 379574
rect 216864 379510 216916 379516
rect 217048 377256 217100 377262
rect 217048 377198 217100 377204
rect 217060 376990 217088 377198
rect 217048 376984 217100 376990
rect 217048 376926 217100 376932
rect 216784 373966 216996 373994
rect 216968 307737 216996 373966
rect 216954 307728 217010 307737
rect 216954 307663 217010 307672
rect 217060 305017 217088 376926
rect 217046 305008 217102 305017
rect 217046 304943 217102 304952
rect 217152 303929 217180 380666
rect 217324 379704 217376 379710
rect 217322 379672 217324 379681
rect 217376 379672 217378 379681
rect 217322 379607 217378 379616
rect 217324 379568 217376 379574
rect 217324 379510 217376 379516
rect 217232 358284 217284 358290
rect 217232 358226 217284 358232
rect 217138 303920 217194 303929
rect 217138 303855 217194 303864
rect 217046 302152 217102 302161
rect 217046 302087 217102 302096
rect 216680 284300 216732 284306
rect 216680 284242 216732 284248
rect 216692 284073 216720 284242
rect 216678 284064 216734 284073
rect 216678 283999 216734 284008
rect 216680 282872 216732 282878
rect 216680 282814 216732 282820
rect 216692 282441 216720 282814
rect 216772 282804 216824 282810
rect 216772 282746 216824 282752
rect 216678 282432 216734 282441
rect 216678 282367 216734 282376
rect 216784 282169 216812 282746
rect 216770 282160 216826 282169
rect 216770 282095 216826 282104
rect 216956 270496 217008 270502
rect 216956 270438 217008 270444
rect 216968 269754 216996 270438
rect 216956 269748 217008 269754
rect 216956 269690 217008 269696
rect 216862 203008 216918 203017
rect 216862 202943 216918 202952
rect 216680 178016 216732 178022
rect 216680 177958 216732 177964
rect 216692 177041 216720 177958
rect 216678 177032 216734 177041
rect 216678 176967 216734 176976
rect 216680 175976 216732 175982
rect 216680 175918 216732 175924
rect 216692 175409 216720 175918
rect 216678 175400 216734 175409
rect 216678 175335 216734 175344
rect 216680 175228 216732 175234
rect 216680 175170 216732 175176
rect 216692 175137 216720 175170
rect 216678 175128 216734 175137
rect 216678 175063 216734 175072
rect 216678 162752 216734 162761
rect 216678 162687 216734 162696
rect 216692 161906 216720 162687
rect 216680 161900 216732 161906
rect 216680 161842 216732 161848
rect 216876 95985 216904 202943
rect 216968 161474 216996 269690
rect 217060 195265 217088 302087
rect 217244 270230 217272 358226
rect 217336 302161 217364 379510
rect 217428 378146 217456 490554
rect 217692 472796 217744 472802
rect 217692 472738 217744 472744
rect 217508 468988 217560 468994
rect 217508 468930 217560 468936
rect 217416 378140 217468 378146
rect 217416 378082 217468 378088
rect 217520 375902 217548 468930
rect 217600 468920 217652 468926
rect 217600 468862 217652 468868
rect 217612 380934 217640 468862
rect 217704 412049 217732 472738
rect 217968 469056 218020 469062
rect 217968 468998 218020 469004
rect 217782 417888 217838 417897
rect 217782 417823 217838 417832
rect 217690 412040 217746 412049
rect 217690 411975 217746 411984
rect 217600 380928 217652 380934
rect 217600 380870 217652 380876
rect 217600 379636 217652 379642
rect 217600 379578 217652 379584
rect 217508 375896 217560 375902
rect 217508 375838 217560 375844
rect 217416 375828 217468 375834
rect 217416 375770 217468 375776
rect 217428 375737 217456 375770
rect 217414 375728 217470 375737
rect 217414 375663 217470 375672
rect 217506 310856 217562 310865
rect 217506 310791 217562 310800
rect 217414 310040 217470 310049
rect 217414 309975 217470 309984
rect 217322 302152 217378 302161
rect 217322 302087 217378 302096
rect 217232 270224 217284 270230
rect 217232 270166 217284 270172
rect 217322 270056 217378 270065
rect 217140 270020 217192 270026
rect 217322 269991 217324 270000
rect 217140 269962 217192 269968
rect 217376 269991 217378 270000
rect 217324 269962 217376 269968
rect 217046 195256 217102 195265
rect 217046 195191 217102 195200
rect 217152 163742 217180 269962
rect 217232 269000 217284 269006
rect 217232 268942 217284 268948
rect 217140 163736 217192 163742
rect 217140 163678 217192 163684
rect 217244 162858 217272 268942
rect 217428 203017 217456 309975
rect 217520 203969 217548 310791
rect 217612 307873 217640 379578
rect 217704 377262 217732 411975
rect 217692 377256 217744 377262
rect 217692 377198 217744 377204
rect 217796 310865 217824 417823
rect 217874 416936 217930 416945
rect 217874 416871 217930 416880
rect 217782 310856 217838 310865
rect 217782 310791 217838 310800
rect 217888 310049 217916 416871
rect 217980 409902 218008 468998
rect 217968 409896 218020 409902
rect 217968 409838 218020 409844
rect 217966 379808 218022 379817
rect 217966 379743 218022 379752
rect 217980 379710 218008 379743
rect 217968 379704 218020 379710
rect 217968 379646 218020 379652
rect 217874 310040 217930 310049
rect 217874 309975 217930 309984
rect 217598 307864 217654 307873
rect 217598 307799 217654 307808
rect 217506 203960 217562 203969
rect 217506 203895 217562 203904
rect 217414 203008 217470 203017
rect 217414 202943 217470 202952
rect 217414 198792 217470 198801
rect 217414 198727 217470 198736
rect 217232 162852 217284 162858
rect 217232 162794 217284 162800
rect 216968 161446 217272 161474
rect 217244 145790 217272 161446
rect 217232 145784 217284 145790
rect 217232 145726 217284 145732
rect 217140 145104 217192 145110
rect 217140 145046 217192 145052
rect 216862 95976 216918 95985
rect 216862 95911 216918 95920
rect 216772 68944 216824 68950
rect 216772 68886 216824 68892
rect 216680 68400 216732 68406
rect 216678 68368 216680 68377
rect 216732 68368 216734 68377
rect 216678 68303 216734 68312
rect 216784 68105 216812 68886
rect 216770 68096 216826 68105
rect 216770 68031 216826 68040
rect 216588 57588 216640 57594
rect 216588 57530 216640 57536
rect 217152 56166 217180 145046
rect 217140 56160 217192 56166
rect 217140 56102 217192 56108
rect 217244 54738 217272 145726
rect 217428 92857 217456 198727
rect 217520 96937 217548 203895
rect 217612 200841 217640 307799
rect 217690 307728 217746 307737
rect 217690 307663 217746 307672
rect 217704 306785 217732 307663
rect 217690 306776 217746 306785
rect 217690 306711 217746 306720
rect 217598 200832 217654 200841
rect 217598 200767 217654 200776
rect 217506 96928 217562 96937
rect 217506 96863 217562 96872
rect 217508 96620 217560 96626
rect 217508 96562 217560 96568
rect 217414 92848 217470 92857
rect 217414 92783 217470 92792
rect 217520 56506 217548 96562
rect 217612 93809 217640 200767
rect 217704 199889 217732 306711
rect 217874 305008 217930 305017
rect 217874 304943 217930 304952
rect 217782 303920 217838 303929
rect 217782 303855 217838 303864
rect 217690 199880 217746 199889
rect 217690 199815 217746 199824
rect 217704 198801 217732 199815
rect 217690 198792 217746 198801
rect 217690 198727 217746 198736
rect 217796 197033 217824 303855
rect 217888 198121 217916 304943
rect 217980 269006 218008 379646
rect 218164 379302 218192 491166
rect 218256 379438 218284 493037
rect 218716 490006 218744 493037
rect 219176 490482 219204 493037
rect 219256 491292 219308 491298
rect 219256 491234 219308 491240
rect 219164 490476 219216 490482
rect 219164 490418 219216 490424
rect 218704 490000 218756 490006
rect 218704 489942 218756 489948
rect 218704 487824 218756 487830
rect 218704 487766 218756 487772
rect 218612 409896 218664 409902
rect 218612 409838 218664 409844
rect 218244 379432 218296 379438
rect 218244 379374 218296 379380
rect 218152 379296 218204 379302
rect 218152 379238 218204 379244
rect 218256 378282 218284 379374
rect 218336 378752 218388 378758
rect 218336 378694 218388 378700
rect 218348 378282 218376 378694
rect 218244 378276 218296 378282
rect 218244 378218 218296 378224
rect 218336 378276 218388 378282
rect 218336 378218 218388 378224
rect 218624 376106 218652 409838
rect 218612 376100 218664 376106
rect 218612 376042 218664 376048
rect 218520 358760 218572 358766
rect 218520 358702 218572 358708
rect 218532 269346 218560 358702
rect 218612 358488 218664 358494
rect 218612 358430 218664 358436
rect 218520 269340 218572 269346
rect 218520 269282 218572 269288
rect 218624 269278 218652 358430
rect 218612 269272 218664 269278
rect 218612 269214 218664 269220
rect 217968 269000 218020 269006
rect 217968 268942 218020 268948
rect 217968 252544 218020 252550
rect 217966 252512 217968 252521
rect 218020 252512 218022 252521
rect 217966 252447 218022 252456
rect 218428 252476 218480 252482
rect 218428 252418 218480 252424
rect 217874 198112 217930 198121
rect 217874 198047 217930 198056
rect 217782 197024 217838 197033
rect 217782 196959 217838 196968
rect 217690 195256 217746 195265
rect 217690 195191 217746 195200
rect 217598 93800 217654 93809
rect 217598 93735 217654 93744
rect 217704 88233 217732 195191
rect 217796 90001 217824 196959
rect 217888 91089 217916 198047
rect 217968 162852 218020 162858
rect 217968 162794 218020 162800
rect 217980 161498 218008 162794
rect 217968 161492 218020 161498
rect 217968 161434 218020 161440
rect 217874 91080 217930 91089
rect 217874 91015 217930 91024
rect 217782 89992 217838 90001
rect 217782 89927 217838 89936
rect 217690 88224 217746 88233
rect 217690 88159 217746 88168
rect 217980 59702 218008 161434
rect 218440 146169 218468 252418
rect 218612 251932 218664 251938
rect 218612 251874 218664 251880
rect 218520 251864 218572 251870
rect 218520 251806 218572 251812
rect 218532 162994 218560 251806
rect 218520 162988 218572 162994
rect 218520 162930 218572 162936
rect 218624 162654 218652 251874
rect 218612 162648 218664 162654
rect 218610 162616 218612 162625
rect 218664 162616 218666 162625
rect 218610 162551 218666 162560
rect 218426 146160 218482 146169
rect 218426 146095 218482 146104
rect 218440 144945 218468 146095
rect 218520 145648 218572 145654
rect 218520 145590 218572 145596
rect 218426 144936 218482 144945
rect 218532 144906 218560 145590
rect 218612 145036 218664 145042
rect 218612 144978 218664 144984
rect 218426 144871 218482 144880
rect 218520 144900 218572 144906
rect 218520 144842 218572 144848
rect 217968 59696 218020 59702
rect 217968 59638 218020 59644
rect 217508 56500 217560 56506
rect 217508 56442 217560 56448
rect 218532 55214 218560 144842
rect 218624 56098 218652 144978
rect 218716 57254 218744 487766
rect 218978 468616 219034 468625
rect 218978 468551 219034 468560
rect 218794 468480 218850 468489
rect 218794 468415 218850 468424
rect 218808 57322 218836 468415
rect 218888 467152 218940 467158
rect 218888 467094 218940 467100
rect 218900 165170 218928 467094
rect 218888 165164 218940 165170
rect 218888 165106 218940 165112
rect 218886 163568 218942 163577
rect 218886 163503 218888 163512
rect 218940 163503 218942 163512
rect 218888 163474 218940 163480
rect 218886 162752 218942 162761
rect 218886 162687 218888 162696
rect 218940 162687 218942 162696
rect 218888 162658 218940 162664
rect 218888 144968 218940 144974
rect 218888 144910 218940 144916
rect 218796 57316 218848 57322
rect 218796 57258 218848 57264
rect 218704 57248 218756 57254
rect 218704 57190 218756 57196
rect 218612 56092 218664 56098
rect 218612 56034 218664 56040
rect 218520 55208 218572 55214
rect 218520 55150 218572 55156
rect 218900 54942 218928 144910
rect 218992 57662 219020 468551
rect 219164 465996 219216 466002
rect 219164 465938 219216 465944
rect 219070 465896 219126 465905
rect 219070 465831 219126 465840
rect 219084 165442 219112 465831
rect 219176 270978 219204 465938
rect 219268 379642 219296 491234
rect 219256 379636 219308 379642
rect 219256 379578 219308 379584
rect 219440 379636 219492 379642
rect 219440 379578 219492 379584
rect 219346 379536 219402 379545
rect 219346 379471 219402 379480
rect 219254 377904 219310 377913
rect 219254 377839 219310 377848
rect 219268 377194 219296 377839
rect 219256 377188 219308 377194
rect 219256 377130 219308 377136
rect 219164 270972 219216 270978
rect 219164 270914 219216 270920
rect 219164 269136 219216 269142
rect 219164 269078 219216 269084
rect 219072 165436 219124 165442
rect 219072 165378 219124 165384
rect 219072 163736 219124 163742
rect 219072 163678 219124 163684
rect 219084 59634 219112 163678
rect 219176 145858 219204 269078
rect 219268 252482 219296 377130
rect 219256 252476 219308 252482
rect 219256 252418 219308 252424
rect 219256 163532 219308 163538
rect 219256 163474 219308 163480
rect 219164 145852 219216 145858
rect 219164 145794 219216 145800
rect 219072 59628 219124 59634
rect 219072 59570 219124 59576
rect 219070 59528 219126 59537
rect 219070 59463 219126 59472
rect 219084 58682 219112 59463
rect 219072 58676 219124 58682
rect 219072 58618 219124 58624
rect 218980 57656 219032 57662
rect 218980 57598 219032 57604
rect 218888 54936 218940 54942
rect 218888 54878 218940 54884
rect 219176 54806 219204 145794
rect 219268 55078 219296 163474
rect 219360 58818 219388 379471
rect 219452 376038 219480 379578
rect 219544 379506 219572 493037
rect 219900 491496 219952 491502
rect 219900 491438 219952 491444
rect 219624 490000 219676 490006
rect 219624 489942 219676 489948
rect 219532 379500 219584 379506
rect 219532 379442 219584 379448
rect 219532 378752 219584 378758
rect 219532 378694 219584 378700
rect 219440 376032 219492 376038
rect 219440 375974 219492 375980
rect 219440 375692 219492 375698
rect 219440 375634 219492 375640
rect 219452 270094 219480 375634
rect 219544 373994 219572 378694
rect 219636 378622 219664 489942
rect 219808 382968 219860 382974
rect 219808 382910 219860 382916
rect 219716 379772 219768 379778
rect 219716 379714 219768 379720
rect 219624 378616 219676 378622
rect 219624 378558 219676 378564
rect 219544 373966 219664 373994
rect 219532 271788 219584 271794
rect 219532 271730 219584 271736
rect 219544 271114 219572 271730
rect 219532 271108 219584 271114
rect 219532 271050 219584 271056
rect 219440 270088 219492 270094
rect 219440 270030 219492 270036
rect 219440 269340 219492 269346
rect 219440 269282 219492 269288
rect 219452 156534 219480 269282
rect 219544 164218 219572 271050
rect 219636 270366 219664 373966
rect 219624 270360 219676 270366
rect 219624 270302 219676 270308
rect 219728 268938 219756 379714
rect 219820 376650 219848 382910
rect 219912 379030 219940 491438
rect 220004 379137 220032 493037
rect 220096 493023 220478 493051
rect 220096 491502 220124 493023
rect 220084 491496 220136 491502
rect 220084 491438 220136 491444
rect 220924 465730 220952 493037
rect 221384 466410 221412 493037
rect 221372 466404 221424 466410
rect 221372 466346 221424 466352
rect 221752 465798 221780 493037
rect 222212 489190 222240 493037
rect 222200 489184 222252 489190
rect 222200 489126 222252 489132
rect 222672 472734 222700 493037
rect 223132 490618 223160 493037
rect 223592 490686 223620 493037
rect 223580 490680 223632 490686
rect 223580 490622 223632 490628
rect 223120 490612 223172 490618
rect 223120 490554 223172 490560
rect 223960 481001 223988 493037
rect 223946 480992 224002 481001
rect 223946 480927 224002 480936
rect 222660 472728 222712 472734
rect 222660 472670 222712 472676
rect 221740 465792 221792 465798
rect 224420 465769 224448 493037
rect 224880 491201 224908 493037
rect 224866 491192 224922 491201
rect 224866 491127 224922 491136
rect 225340 490754 225368 493037
rect 225328 490748 225380 490754
rect 225328 490690 225380 490696
rect 225708 490657 225736 493037
rect 226168 490793 226196 493037
rect 226154 490784 226210 490793
rect 226154 490719 226210 490728
rect 225694 490648 225750 490657
rect 225694 490583 225750 490592
rect 226628 490521 226656 493037
rect 226614 490512 226670 490521
rect 226614 490447 226670 490456
rect 227088 472802 227116 493037
rect 227076 472796 227128 472802
rect 227076 472738 227128 472744
rect 227548 472666 227576 493037
rect 227916 479602 227944 493037
rect 228376 483721 228404 493037
rect 228836 487801 228864 493037
rect 228822 487792 228878 487801
rect 228822 487727 228878 487736
rect 229296 486441 229324 493037
rect 229282 486432 229338 486441
rect 229282 486367 229338 486376
rect 229756 485081 229784 493037
rect 229742 485072 229798 485081
rect 229742 485007 229798 485016
rect 228362 483712 228418 483721
rect 228362 483647 228418 483656
rect 227904 479596 227956 479602
rect 227904 479538 227956 479544
rect 230124 474065 230152 493037
rect 230584 490793 230612 493037
rect 230570 490784 230626 490793
rect 230570 490719 230626 490728
rect 231044 475425 231072 493037
rect 231504 490929 231532 493037
rect 231490 490920 231546 490929
rect 231490 490855 231546 490864
rect 231872 483750 231900 493037
rect 232332 490521 232360 493037
rect 232318 490512 232374 490521
rect 232318 490447 232374 490456
rect 231860 483744 231912 483750
rect 231860 483686 231912 483692
rect 232792 476814 232820 493037
rect 233252 490822 233280 493037
rect 233240 490816 233292 490822
rect 233240 490758 233292 490764
rect 232780 476808 232832 476814
rect 232780 476750 232832 476756
rect 231030 475416 231086 475425
rect 231030 475351 231086 475360
rect 230110 474056 230166 474065
rect 230110 473991 230166 474000
rect 227536 472660 227588 472666
rect 227536 472602 227588 472608
rect 233712 472569 233740 493037
rect 234080 490657 234108 493037
rect 234066 490648 234122 490657
rect 234066 490583 234122 490592
rect 234540 476785 234568 493037
rect 235000 491201 235028 493037
rect 234986 491192 235042 491201
rect 234986 491127 235042 491136
rect 235460 482361 235488 493037
rect 235446 482352 235502 482361
rect 235446 482287 235502 482296
rect 235920 479505 235948 493037
rect 236288 491065 236316 493037
rect 236274 491056 236330 491065
rect 236274 490991 236330 491000
rect 236748 487830 236776 493037
rect 236736 487824 236788 487830
rect 236736 487766 236788 487772
rect 235906 479496 235962 479505
rect 235906 479431 235962 479440
rect 234526 476776 234582 476785
rect 234526 476711 234582 476720
rect 237208 474094 237236 493037
rect 237668 490890 237696 493037
rect 237656 490884 237708 490890
rect 237656 490826 237708 490832
rect 238128 479670 238156 493037
rect 238496 483682 238524 493037
rect 238956 490958 238984 493037
rect 239416 491026 239444 493037
rect 239404 491020 239456 491026
rect 239404 490962 239456 490968
rect 238944 490952 238996 490958
rect 238944 490894 238996 490900
rect 238484 483676 238536 483682
rect 238484 483618 238536 483624
rect 239876 482322 239904 493037
rect 239864 482316 239916 482322
rect 239864 482258 239916 482264
rect 238116 479664 238168 479670
rect 238116 479606 238168 479612
rect 237196 474088 237248 474094
rect 237196 474030 237248 474036
rect 233698 472560 233754 472569
rect 233698 472495 233754 472504
rect 240244 469878 240272 493037
rect 240704 491094 240732 493037
rect 240692 491088 240744 491094
rect 240692 491030 240744 491036
rect 240232 469872 240284 469878
rect 240232 469814 240284 469820
rect 221740 465734 221792 465740
rect 224406 465760 224462 465769
rect 220912 465724 220964 465730
rect 241164 465730 241192 493037
rect 241624 472870 241652 493037
rect 242084 489258 242112 493037
rect 242072 489252 242124 489258
rect 242072 489194 242124 489200
rect 242452 486538 242480 493037
rect 242440 486532 242492 486538
rect 242440 486474 242492 486480
rect 242912 485110 242940 493037
rect 242900 485104 242952 485110
rect 242900 485046 242952 485052
rect 243372 483818 243400 493037
rect 243360 483812 243412 483818
rect 243360 483754 243412 483760
rect 241612 472864 241664 472870
rect 241612 472806 241664 472812
rect 243832 466002 243860 493037
rect 243820 465996 243872 466002
rect 243820 465938 243872 465944
rect 244292 465866 244320 493037
rect 244660 476882 244688 493037
rect 245120 482390 245148 493037
rect 245108 482384 245160 482390
rect 245108 482326 245160 482332
rect 244648 476876 244700 476882
rect 244648 476818 244700 476824
rect 245580 475386 245608 493037
rect 246040 478242 246068 493037
rect 246028 478236 246080 478242
rect 246028 478178 246080 478184
rect 245568 475380 245620 475386
rect 245568 475322 245620 475328
rect 244280 465860 244332 465866
rect 244280 465802 244332 465808
rect 246408 465798 246436 493037
rect 246868 487898 246896 493037
rect 247328 489161 247356 493037
rect 247314 489152 247370 489161
rect 247314 489087 247370 489096
rect 246856 487892 246908 487898
rect 246856 487834 246908 487840
rect 247788 486470 247816 493037
rect 247776 486464 247828 486470
rect 247776 486406 247828 486412
rect 248248 474026 248276 493037
rect 248616 491162 248644 493037
rect 248604 491156 248656 491162
rect 248604 491098 248656 491104
rect 248236 474020 248288 474026
rect 248236 473962 248288 473968
rect 249076 467158 249104 493037
rect 249536 467362 249564 493037
rect 249524 467356 249576 467362
rect 249524 467298 249576 467304
rect 249996 467294 250024 493037
rect 249984 467288 250036 467294
rect 249984 467230 250036 467236
rect 250456 467226 250484 493037
rect 250824 470014 250852 493037
rect 250812 470008 250864 470014
rect 250812 469950 250864 469956
rect 251284 469946 251312 493037
rect 251272 469940 251324 469946
rect 251272 469882 251324 469888
rect 251744 467430 251772 493037
rect 252204 467498 252232 493037
rect 252572 475561 252600 493037
rect 253032 482458 253060 493037
rect 253020 482452 253072 482458
rect 253020 482394 253072 482400
rect 253492 481137 253520 493037
rect 253478 481128 253534 481137
rect 253478 481063 253534 481072
rect 252558 475552 252614 475561
rect 253952 475522 253980 493037
rect 254412 479738 254440 493037
rect 254400 479732 254452 479738
rect 254400 479674 254452 479680
rect 252558 475487 252614 475496
rect 253940 475516 253992 475522
rect 253940 475458 253992 475464
rect 254780 468518 254808 493037
rect 255240 468586 255268 493037
rect 255700 478145 255728 493037
rect 256160 478446 256188 493037
rect 256148 478440 256200 478446
rect 256148 478382 256200 478388
rect 256620 478378 256648 493037
rect 256988 487966 257016 493037
rect 256976 487960 257028 487966
rect 256976 487902 257028 487908
rect 256608 478372 256660 478378
rect 256608 478314 256660 478320
rect 255686 478136 255742 478145
rect 255686 478071 255742 478080
rect 255228 468580 255280 468586
rect 255228 468522 255280 468528
rect 254768 468512 254820 468518
rect 254768 468454 254820 468460
rect 252192 467492 252244 467498
rect 252192 467434 252244 467440
rect 251732 467424 251784 467430
rect 251732 467366 251784 467372
rect 250444 467220 250496 467226
rect 250444 467162 250496 467168
rect 249064 467152 249116 467158
rect 249064 467094 249116 467100
rect 257448 466138 257476 493037
rect 257908 489326 257936 493037
rect 257896 489320 257948 489326
rect 257896 489262 257948 489268
rect 257436 466132 257488 466138
rect 257436 466074 257488 466080
rect 258368 466070 258396 493037
rect 258828 480962 258856 493037
rect 258816 480956 258868 480962
rect 258816 480898 258868 480904
rect 259196 474162 259224 493037
rect 259656 476950 259684 493037
rect 260116 478310 260144 493037
rect 260576 483886 260604 493037
rect 260944 486606 260972 493037
rect 260932 486600 260984 486606
rect 260932 486542 260984 486548
rect 261404 485178 261432 493037
rect 261392 485172 261444 485178
rect 261392 485114 261444 485120
rect 260564 483880 260616 483886
rect 260564 483822 260616 483828
rect 260104 478304 260156 478310
rect 260104 478246 260156 478252
rect 259644 476944 259696 476950
rect 259644 476886 259696 476892
rect 259184 474156 259236 474162
rect 259184 474098 259236 474104
rect 261864 472938 261892 493037
rect 261852 472932 261904 472938
rect 261852 472874 261904 472880
rect 262324 467634 262352 493037
rect 262312 467628 262364 467634
rect 262312 467570 262364 467576
rect 258356 466064 258408 466070
rect 258356 466006 258408 466012
rect 262784 465934 262812 493037
rect 263152 466274 263180 493037
rect 263140 466268 263192 466274
rect 263140 466210 263192 466216
rect 263612 466206 263640 493037
rect 264072 473278 264100 493037
rect 264060 473272 264112 473278
rect 264060 473214 264112 473220
rect 264532 473210 264560 493037
rect 264520 473204 264572 473210
rect 264520 473146 264572 473152
rect 264992 473006 265020 493037
rect 265360 475454 265388 493037
rect 265348 475448 265400 475454
rect 265348 475390 265400 475396
rect 265820 473142 265848 493037
rect 266280 475658 266308 493037
rect 266268 475652 266320 475658
rect 266268 475594 266320 475600
rect 265808 473136 265860 473142
rect 265808 473078 265860 473084
rect 264980 473000 265032 473006
rect 264980 472942 265032 472948
rect 266740 469062 266768 493037
rect 266728 469056 266780 469062
rect 266728 468998 266780 469004
rect 267108 468994 267136 493037
rect 267568 473074 267596 493037
rect 267556 473068 267608 473074
rect 267556 473010 267608 473016
rect 267096 468988 267148 468994
rect 267096 468930 267148 468936
rect 268028 468654 268056 493037
rect 268488 483954 268516 493037
rect 268948 484022 268976 493037
rect 268936 484016 268988 484022
rect 268936 483958 268988 483964
rect 268476 483948 268528 483954
rect 268476 483890 268528 483896
rect 269316 469198 269344 493037
rect 269776 484226 269804 493037
rect 270236 484294 270264 493037
rect 270224 484288 270276 484294
rect 270224 484230 270276 484236
rect 269764 484220 269816 484226
rect 269764 484162 269816 484168
rect 269304 469192 269356 469198
rect 269304 469134 269356 469140
rect 268016 468648 268068 468654
rect 268016 468590 268068 468596
rect 270696 467566 270724 493037
rect 271156 471306 271184 493037
rect 271524 471374 271552 493037
rect 271512 471368 271564 471374
rect 271512 471310 271564 471316
rect 271144 471300 271196 471306
rect 271144 471242 271196 471248
rect 271984 468722 272012 493037
rect 272444 468790 272472 493037
rect 272904 475590 272932 493037
rect 273272 478514 273300 493037
rect 273732 478582 273760 493037
rect 273720 478576 273772 478582
rect 273720 478518 273772 478524
rect 273260 478508 273312 478514
rect 273260 478450 273312 478456
rect 272892 475584 272944 475590
rect 272892 475526 272944 475532
rect 272432 468784 272484 468790
rect 272432 468726 272484 468732
rect 271972 468716 272024 468722
rect 271972 468658 272024 468664
rect 270684 467560 270736 467566
rect 270684 467502 270736 467508
rect 263600 466200 263652 466206
rect 263600 466142 263652 466148
rect 262772 465928 262824 465934
rect 262772 465870 262824 465876
rect 246396 465792 246448 465798
rect 246396 465734 246448 465740
rect 224406 465695 224462 465704
rect 241152 465724 241204 465730
rect 220912 465666 220964 465672
rect 241152 465666 241204 465672
rect 274192 465662 274220 493037
rect 274652 481098 274680 493037
rect 274640 481092 274692 481098
rect 274640 481034 274692 481040
rect 275112 481030 275140 493037
rect 275100 481024 275152 481030
rect 275100 480966 275152 480972
rect 275480 468858 275508 493037
rect 275468 468852 275520 468858
rect 275468 468794 275520 468800
rect 275940 466342 275968 493037
rect 276400 468489 276428 493037
rect 276386 468480 276442 468489
rect 276386 468415 276442 468424
rect 275928 466336 275980 466342
rect 275928 466278 275980 466284
rect 274180 465656 274232 465662
rect 274180 465598 274232 465604
rect 276860 464370 276888 493037
rect 277320 469130 277348 493037
rect 277688 475726 277716 493037
rect 278148 478650 278176 493037
rect 278608 478718 278636 493037
rect 279068 481302 279096 493037
rect 279056 481296 279108 481302
rect 279056 481238 279108 481244
rect 279528 481234 279556 493037
rect 279516 481228 279568 481234
rect 279516 481170 279568 481176
rect 279896 481166 279924 493037
rect 279884 481160 279936 481166
rect 279884 481102 279936 481108
rect 278596 478712 278648 478718
rect 278596 478654 278648 478660
rect 278136 478644 278188 478650
rect 278136 478586 278188 478592
rect 277676 475720 277728 475726
rect 277676 475662 277728 475668
rect 277308 469124 277360 469130
rect 277308 469066 277360 469072
rect 280356 466410 280384 493037
rect 280816 484158 280844 493037
rect 280804 484152 280856 484158
rect 280804 484094 280856 484100
rect 281276 484090 281304 493037
rect 281264 484084 281316 484090
rect 281264 484026 281316 484032
rect 281644 470422 281672 493037
rect 281632 470416 281684 470422
rect 281632 470358 281684 470364
rect 282104 470082 282132 493037
rect 282564 471442 282592 493037
rect 282552 471436 282604 471442
rect 282552 471378 282604 471384
rect 283024 470490 283052 493037
rect 283484 470558 283512 493037
rect 283852 489394 283880 493037
rect 283840 489388 283892 489394
rect 283840 489330 283892 489336
rect 284312 485246 284340 493037
rect 284300 485240 284352 485246
rect 284300 485182 284352 485188
rect 283472 470552 283524 470558
rect 283472 470494 283524 470500
rect 283012 470484 283064 470490
rect 283012 470426 283064 470432
rect 284772 470150 284800 493037
rect 284760 470144 284812 470150
rect 284760 470086 284812 470092
rect 282092 470076 282144 470082
rect 282092 470018 282144 470024
rect 285232 468926 285260 493037
rect 285692 475794 285720 493037
rect 285680 475788 285732 475794
rect 285680 475730 285732 475736
rect 286060 471782 286088 493037
rect 286048 471776 286100 471782
rect 286048 471718 286100 471724
rect 286520 471578 286548 493037
rect 286508 471572 286560 471578
rect 286508 471514 286560 471520
rect 286980 471510 287008 493037
rect 287440 471646 287468 493037
rect 287808 474230 287836 493037
rect 287796 474224 287848 474230
rect 287796 474166 287848 474172
rect 287428 471640 287480 471646
rect 287428 471582 287480 471588
rect 286968 471504 287020 471510
rect 286968 471446 287020 471452
rect 285220 468920 285272 468926
rect 285220 468862 285272 468868
rect 288268 467702 288296 493037
rect 288256 467696 288308 467702
rect 288256 467638 288308 467644
rect 280344 466404 280396 466410
rect 280344 466346 280396 466352
rect 288728 464438 288756 493037
rect 289188 478786 289216 493037
rect 289648 481370 289676 493037
rect 290016 491230 290044 493037
rect 290004 491224 290056 491230
rect 290004 491166 290056 491172
rect 289636 481364 289688 481370
rect 289636 481306 289688 481312
rect 289176 478780 289228 478786
rect 289176 478722 289228 478728
rect 290476 468382 290504 493037
rect 290936 475862 290964 493037
rect 291396 478854 291424 493037
rect 291856 481438 291884 493037
rect 292224 484362 292252 493037
rect 292212 484356 292264 484362
rect 292212 484298 292264 484304
rect 292684 481506 292712 493037
rect 292672 481500 292724 481506
rect 292672 481442 292724 481448
rect 291844 481432 291896 481438
rect 291844 481374 291896 481380
rect 291384 478848 291436 478854
rect 291384 478790 291436 478796
rect 290924 475856 290976 475862
rect 290924 475798 290976 475804
rect 293144 470286 293172 493037
rect 293604 471714 293632 493037
rect 293592 471708 293644 471714
rect 293592 471650 293644 471656
rect 293132 470280 293184 470286
rect 293132 470222 293184 470228
rect 293972 470218 294000 493037
rect 293960 470212 294012 470218
rect 293960 470154 294012 470160
rect 290464 468376 290516 468382
rect 290464 468318 290516 468324
rect 294432 464506 294460 493037
rect 294892 471850 294920 493037
rect 294880 471844 294932 471850
rect 294880 471786 294932 471792
rect 295352 471481 295380 493037
rect 295338 471472 295394 471481
rect 295338 471407 295394 471416
rect 295812 469810 295840 493037
rect 296180 471209 296208 493037
rect 296166 471200 296222 471209
rect 296166 471135 296222 471144
rect 295800 469804 295852 469810
rect 295800 469746 295852 469752
rect 296640 467838 296668 493037
rect 296628 467832 296680 467838
rect 296628 467774 296680 467780
rect 297100 465594 297128 493037
rect 297560 471345 297588 493037
rect 297546 471336 297602 471345
rect 297546 471271 297602 471280
rect 298020 470354 298048 493037
rect 298008 470348 298060 470354
rect 298008 470290 298060 470296
rect 298388 465905 298416 493037
rect 298848 468450 298876 493037
rect 298836 468444 298888 468450
rect 298836 468386 298888 468392
rect 299308 467770 299336 493037
rect 299768 471918 299796 493068
rect 309796 479534 309824 629274
rect 309888 558278 309916 638930
rect 311176 568002 311204 648110
rect 316776 648100 316828 648106
rect 316776 648042 316828 648048
rect 313924 647488 313976 647494
rect 313924 647430 313976 647436
rect 312544 643136 312596 643142
rect 312544 643078 312596 643084
rect 311256 610020 311308 610026
rect 311256 609962 311308 609968
rect 311164 567996 311216 568002
rect 311164 567938 311216 567944
rect 309876 558272 309928 558278
rect 309876 558214 309928 558220
rect 311268 556850 311296 609962
rect 312556 566710 312584 643078
rect 312636 619676 312688 619682
rect 312636 619618 312688 619624
rect 312544 566704 312596 566710
rect 312544 566646 312596 566652
rect 312648 558346 312676 619618
rect 313936 572150 313964 647430
rect 316682 647320 316738 647329
rect 316682 647255 316738 647264
rect 314108 645040 314160 645046
rect 314108 644982 314160 644988
rect 314016 644836 314068 644842
rect 314016 644778 314068 644784
rect 314028 578882 314056 644778
rect 314016 578876 314068 578882
rect 314016 578818 314068 578824
rect 314120 578746 314148 644982
rect 314200 615528 314252 615534
rect 314200 615470 314252 615476
rect 314108 578740 314160 578746
rect 314108 578682 314160 578688
rect 313924 572144 313976 572150
rect 313924 572086 313976 572092
rect 314212 566642 314240 615470
rect 314200 566636 314252 566642
rect 314200 566578 314252 566584
rect 316696 559706 316724 647255
rect 316788 565282 316816 648042
rect 323768 648032 323820 648038
rect 323768 647974 323820 647980
rect 322388 647964 322440 647970
rect 322388 647906 322440 647912
rect 322296 647896 322348 647902
rect 322296 647838 322348 647844
rect 318156 647760 318208 647766
rect 318156 647702 318208 647708
rect 316868 646196 316920 646202
rect 316868 646138 316920 646144
rect 316880 579562 316908 646138
rect 318064 644972 318116 644978
rect 318064 644914 318116 644920
rect 316960 644700 317012 644706
rect 316960 644642 317012 644648
rect 316868 579556 316920 579562
rect 316868 579498 316920 579504
rect 316972 579426 317000 644642
rect 317052 644632 317104 644638
rect 317052 644574 317104 644580
rect 317064 579494 317092 644574
rect 317144 590708 317196 590714
rect 317144 590650 317196 590656
rect 317052 579488 317104 579494
rect 317052 579430 317104 579436
rect 316960 579420 317012 579426
rect 316960 579362 317012 579368
rect 317156 570858 317184 590650
rect 317144 570852 317196 570858
rect 317144 570794 317196 570800
rect 316776 565276 316828 565282
rect 316776 565218 316828 565224
rect 316684 559700 316736 559706
rect 316684 559642 316736 559648
rect 312636 558340 312688 558346
rect 312636 558282 312688 558288
rect 316776 557932 316828 557938
rect 316776 557874 316828 557880
rect 311256 556844 311308 556850
rect 311256 556786 311308 556792
rect 316684 556640 316736 556646
rect 316684 556582 316736 556588
rect 316696 529786 316724 556582
rect 316788 531010 316816 557874
rect 316868 556708 316920 556714
rect 316868 556650 316920 556656
rect 316776 531004 316828 531010
rect 316776 530946 316828 530952
rect 316880 530874 316908 556650
rect 318076 555490 318104 644914
rect 318168 563922 318196 647702
rect 320916 647692 320968 647698
rect 320916 647634 320968 647640
rect 320824 647420 320876 647426
rect 320824 647362 320876 647368
rect 319444 646332 319496 646338
rect 319444 646274 319496 646280
rect 319456 579358 319484 646274
rect 319536 646128 319588 646134
rect 319536 646070 319588 646076
rect 319444 579352 319496 579358
rect 319444 579294 319496 579300
rect 319548 578814 319576 646070
rect 319628 644768 319680 644774
rect 319628 644710 319680 644716
rect 319640 579630 319668 644710
rect 319628 579624 319680 579630
rect 319628 579566 319680 579572
rect 319536 578808 319588 578814
rect 319536 578750 319588 578756
rect 318156 563916 318208 563922
rect 318156 563858 318208 563864
rect 320836 563854 320864 647362
rect 320928 573510 320956 647634
rect 322204 647352 322256 647358
rect 322204 647294 322256 647300
rect 321008 643748 321060 643754
rect 321008 643690 321060 643696
rect 321020 582321 321048 643690
rect 321558 643648 321614 643657
rect 321558 643583 321614 643592
rect 321572 643142 321600 643583
rect 321560 643136 321612 643142
rect 321560 643078 321612 643084
rect 321558 639024 321614 639033
rect 321558 638959 321560 638968
rect 321612 638959 321614 638968
rect 321560 638930 321612 638936
rect 321558 634128 321614 634137
rect 321558 634063 321614 634072
rect 321572 633486 321600 634063
rect 321560 633480 321612 633486
rect 321560 633422 321612 633428
rect 321558 629504 321614 629513
rect 321558 629439 321614 629448
rect 321572 629338 321600 629439
rect 321560 629332 321612 629338
rect 321560 629274 321612 629280
rect 321558 625288 321614 625297
rect 321558 625223 321614 625232
rect 321572 625190 321600 625223
rect 321560 625184 321612 625190
rect 321560 625126 321612 625132
rect 321558 619984 321614 619993
rect 321558 619919 321614 619928
rect 321572 619682 321600 619919
rect 321560 619676 321612 619682
rect 321560 619618 321612 619624
rect 321558 615632 321614 615641
rect 321558 615567 321614 615576
rect 321572 615534 321600 615567
rect 321560 615528 321612 615534
rect 321560 615470 321612 615476
rect 321558 610328 321614 610337
rect 321558 610263 321614 610272
rect 321572 610026 321600 610263
rect 321560 610020 321612 610026
rect 321560 609962 321612 609968
rect 321558 600808 321614 600817
rect 321558 600743 321614 600752
rect 321572 600370 321600 600743
rect 321560 600364 321612 600370
rect 321560 600306 321612 600312
rect 321558 596456 321614 596465
rect 321558 596391 321614 596400
rect 321572 596222 321600 596391
rect 321560 596216 321612 596222
rect 321560 596158 321612 596164
rect 321558 591288 321614 591297
rect 321558 591223 321614 591232
rect 321572 590714 321600 591223
rect 321560 590708 321612 590714
rect 321560 590650 321612 590656
rect 321098 585848 321154 585857
rect 321098 585783 321154 585792
rect 321006 582312 321062 582321
rect 321006 582247 321062 582256
rect 320916 573504 320968 573510
rect 320916 573446 320968 573452
rect 320824 563848 320876 563854
rect 320824 563790 320876 563796
rect 321112 559638 321140 585783
rect 321834 576872 321890 576881
rect 321834 576807 321890 576816
rect 321848 574802 321876 576807
rect 321836 574796 321888 574802
rect 321836 574738 321888 574744
rect 321558 571704 321614 571713
rect 321558 571639 321614 571648
rect 321572 571402 321600 571639
rect 321560 571396 321612 571402
rect 321560 571338 321612 571344
rect 322216 569362 322244 647294
rect 322308 575006 322336 647838
rect 322400 577590 322428 647906
rect 323584 647828 323636 647834
rect 323584 647770 323636 647776
rect 322572 646468 322624 646474
rect 322572 646410 322624 646416
rect 322480 646400 322532 646406
rect 322480 646342 322532 646348
rect 322492 579290 322520 646342
rect 322480 579284 322532 579290
rect 322480 579226 322532 579232
rect 322584 579222 322612 646410
rect 322664 645108 322716 645114
rect 322664 645050 322716 645056
rect 322676 609278 322704 645050
rect 322664 609272 322716 609278
rect 322664 609214 322716 609220
rect 322572 579216 322624 579222
rect 322572 579158 322624 579164
rect 322388 577584 322440 577590
rect 322388 577526 322440 577532
rect 322296 575000 322348 575006
rect 322296 574942 322348 574948
rect 322204 569356 322256 569362
rect 322204 569298 322256 569304
rect 321558 567352 321614 567361
rect 321558 567287 321614 567296
rect 321572 567254 321600 567287
rect 321560 567248 321612 567254
rect 321560 567190 321612 567196
rect 321560 563032 321612 563038
rect 321560 562974 321612 562980
rect 321572 562873 321600 562974
rect 321558 562864 321614 562873
rect 321558 562799 321614 562808
rect 323596 561066 323624 647770
rect 323676 647284 323728 647290
rect 323676 647226 323728 647232
rect 323688 569294 323716 647226
rect 323780 570790 323808 647974
rect 324240 606801 324268 649266
rect 337568 648168 337620 648174
rect 337568 648110 337620 648116
rect 324872 647624 324924 647630
rect 324872 647566 324924 647572
rect 324780 647556 324832 647562
rect 324780 647498 324832 647504
rect 324226 606792 324282 606801
rect 324226 606727 324282 606736
rect 324792 577522 324820 647498
rect 324780 577516 324832 577522
rect 324780 577458 324832 577464
rect 323860 576156 323912 576162
rect 323860 576098 323912 576104
rect 323768 570784 323820 570790
rect 323768 570726 323820 570732
rect 323676 569288 323728 569294
rect 323676 569230 323728 569236
rect 323584 561060 323636 561066
rect 323584 561002 323636 561008
rect 321100 559632 321152 559638
rect 321100 559574 321152 559580
rect 319444 557864 319496 557870
rect 319444 557806 319496 557812
rect 321558 557832 321614 557841
rect 318156 556232 318208 556238
rect 318156 556174 318208 556180
rect 318064 555484 318116 555490
rect 318064 555426 318116 555432
rect 316958 553752 317014 553761
rect 316958 553687 317014 553696
rect 316868 530868 316920 530874
rect 316868 530810 316920 530816
rect 316972 529922 317000 553687
rect 318168 532030 318196 556174
rect 318156 532024 318208 532030
rect 318156 531966 318208 531972
rect 316960 529916 317012 529922
rect 316960 529858 317012 529864
rect 316684 529780 316736 529786
rect 316684 529722 316736 529728
rect 319456 529650 319484 557806
rect 321558 557767 321614 557776
rect 322204 557796 322256 557802
rect 321572 557734 321600 557767
rect 322204 557738 322256 557744
rect 321560 557728 321612 557734
rect 321560 557670 321612 557676
rect 319720 557660 319772 557666
rect 319720 557602 319772 557608
rect 319536 553648 319588 553654
rect 319536 553590 319588 553596
rect 319444 529644 319496 529650
rect 319444 529586 319496 529592
rect 319548 529582 319576 553590
rect 319626 553480 319682 553489
rect 319626 553415 319682 553424
rect 319640 529854 319668 553415
rect 319732 533798 319760 557602
rect 320824 556436 320876 556442
rect 320824 556378 320876 556384
rect 319810 553616 319866 553625
rect 319810 553551 319866 553560
rect 319720 533792 319772 533798
rect 319720 533734 319772 533740
rect 319628 529848 319680 529854
rect 319628 529790 319680 529796
rect 319824 529718 319852 553551
rect 320836 532098 320864 556378
rect 321652 554260 321704 554266
rect 321652 554202 321704 554208
rect 321560 553376 321612 553382
rect 321558 553344 321560 553353
rect 321612 553344 321614 553353
rect 321558 553279 321614 553288
rect 321664 549001 321692 554202
rect 321650 548992 321706 549001
rect 321650 548927 321706 548936
rect 321560 543720 321612 543726
rect 321558 543688 321560 543697
rect 321612 543688 321614 543697
rect 321558 543623 321614 543632
rect 321560 539572 321612 539578
rect 321560 539514 321612 539520
rect 321572 539345 321600 539514
rect 321558 539336 321614 539345
rect 321558 539271 321614 539280
rect 320824 532092 320876 532098
rect 320824 532034 320876 532040
rect 319812 529712 319864 529718
rect 319812 529654 319864 529660
rect 319536 529576 319588 529582
rect 319536 529518 319588 529524
rect 322216 529514 322244 557738
rect 322296 557592 322348 557598
rect 322296 557534 322348 557540
rect 322308 533458 322336 557534
rect 323676 556504 323728 556510
rect 323676 556446 323728 556452
rect 323584 556300 323636 556306
rect 323584 556242 323636 556248
rect 322386 555248 322442 555257
rect 322386 555183 322442 555192
rect 322296 533452 322348 533458
rect 322296 533394 322348 533400
rect 322400 531214 322428 555183
rect 322480 555144 322532 555150
rect 322480 555086 322532 555092
rect 322388 531208 322440 531214
rect 322388 531150 322440 531156
rect 322492 531146 322520 555086
rect 322664 555076 322716 555082
rect 322664 555018 322716 555024
rect 322572 553580 322624 553586
rect 322572 553522 322624 553528
rect 322584 532642 322612 553522
rect 322676 533730 322704 555018
rect 322756 553104 322808 553110
rect 322756 553046 322808 553052
rect 322664 533724 322716 533730
rect 322664 533666 322716 533672
rect 322572 532636 322624 532642
rect 322572 532578 322624 532584
rect 322768 532545 322796 553046
rect 322754 532536 322810 532545
rect 322754 532471 322810 532480
rect 323596 532438 323624 556242
rect 323584 532432 323636 532438
rect 323584 532374 323636 532380
rect 323688 532370 323716 556446
rect 323768 555620 323820 555626
rect 323768 555562 323820 555568
rect 323780 533662 323808 555562
rect 323768 533656 323820 533662
rect 323768 533598 323820 533604
rect 323872 532409 323900 576098
rect 324884 567934 324912 647566
rect 328552 647284 328604 647290
rect 328552 647226 328604 647232
rect 328564 644994 328592 647226
rect 333058 646232 333114 646241
rect 333058 646167 333114 646176
rect 333072 644994 333100 646167
rect 337580 644994 337608 648110
rect 342260 648100 342312 648106
rect 342260 648042 342312 648048
rect 342272 644994 342300 648042
rect 401692 648032 401744 648038
rect 401692 647974 401744 647980
rect 346584 647964 346636 647970
rect 346584 647906 346636 647912
rect 346596 644994 346624 647906
rect 355600 647896 355652 647902
rect 355600 647838 355652 647844
rect 351090 646096 351146 646105
rect 351090 646031 351146 646040
rect 351104 644994 351132 646031
rect 355612 644994 355640 647838
rect 369124 647828 369176 647834
rect 369124 647770 369176 647776
rect 364616 647760 364668 647766
rect 364616 647702 364668 647708
rect 360200 646264 360252 646270
rect 360200 646206 360252 646212
rect 360212 644994 360240 646206
rect 364628 644994 364656 647702
rect 369136 644994 369164 647770
rect 374000 647692 374052 647698
rect 374000 647634 374052 647640
rect 374012 644994 374040 647634
rect 378140 647624 378192 647630
rect 378140 647566 378192 647572
rect 328564 644966 328900 644994
rect 333072 644966 333408 644994
rect 337580 644966 337916 644994
rect 342272 644966 342424 644994
rect 346596 644966 346932 644994
rect 351104 644966 351440 644994
rect 355612 644966 355948 644994
rect 360212 644966 360456 644994
rect 364628 644966 364964 644994
rect 369136 644966 369472 644994
rect 373980 644966 374040 644994
rect 378152 644994 378180 647566
rect 387800 647556 387852 647562
rect 387800 647498 387852 647504
rect 383660 647488 383712 647494
rect 383660 647430 383712 647436
rect 383672 644994 383700 647430
rect 378152 644966 378488 644994
rect 383640 644966 383700 644994
rect 387812 644994 387840 647498
rect 392308 647420 392360 647426
rect 392308 647362 392360 647368
rect 391940 647284 391992 647290
rect 391940 647226 391992 647232
rect 391952 646542 391980 647226
rect 391940 646536 391992 646542
rect 391940 646478 391992 646484
rect 392320 644994 392348 647362
rect 396816 647284 396868 647290
rect 396816 647226 396868 647232
rect 396828 644994 396856 647226
rect 387812 644966 388148 644994
rect 392320 644966 392656 644994
rect 396828 644966 397164 644994
rect 401704 644858 401732 647974
rect 405844 644994 405872 651986
rect 423862 647320 423918 647329
rect 419540 647284 419592 647290
rect 423862 647255 423918 647264
rect 419540 647226 419592 647232
rect 414848 645992 414900 645998
rect 410338 645960 410394 645969
rect 414848 645934 414900 645940
rect 410338 645895 410394 645904
rect 410352 644994 410380 645895
rect 414860 644994 414888 645934
rect 419552 645930 419580 647226
rect 419540 645924 419592 645930
rect 419540 645866 419592 645872
rect 419552 644994 419580 645866
rect 423876 644994 423904 647255
rect 428292 644994 428320 654106
rect 432880 647352 432932 647358
rect 432880 647294 432932 647300
rect 432892 644994 432920 647294
rect 433340 646060 433392 646066
rect 433340 646002 433392 646008
rect 405844 644966 406180 644994
rect 410352 644966 410688 644994
rect 414860 644966 415196 644994
rect 419552 644966 419704 644994
rect 423876 644966 424212 644994
rect 428292 644966 428720 644994
rect 432892 644966 433228 644994
rect 401672 644830 401732 644858
rect 433352 630873 433380 646002
rect 433338 630864 433394 630873
rect 433338 630799 433394 630808
rect 433338 611416 433394 611425
rect 433338 611351 433394 611360
rect 324872 567928 324924 567934
rect 324872 567870 324924 567876
rect 324872 556368 324924 556374
rect 324872 556310 324924 556316
rect 324688 555688 324740 555694
rect 324688 555630 324740 555636
rect 323950 555520 324006 555529
rect 323950 555455 324006 555464
rect 323964 533594 323992 555455
rect 324136 555416 324188 555422
rect 324136 555358 324188 555364
rect 324044 554192 324096 554198
rect 324044 554134 324096 554140
rect 323952 533588 324004 533594
rect 323952 533530 324004 533536
rect 324056 532710 324084 554134
rect 324148 535430 324176 555358
rect 324320 554056 324372 554062
rect 324320 553998 324372 554004
rect 324136 535424 324188 535430
rect 324136 535366 324188 535372
rect 324332 534614 324360 553998
rect 324596 553920 324648 553926
rect 324596 553862 324648 553868
rect 324320 534608 324372 534614
rect 324320 534550 324372 534556
rect 324044 532704 324096 532710
rect 324044 532646 324096 532652
rect 323858 532400 323914 532409
rect 323676 532364 323728 532370
rect 323858 532335 323914 532344
rect 323676 532306 323728 532312
rect 324608 531826 324636 553862
rect 324700 533526 324728 555630
rect 324780 553716 324832 553722
rect 324780 553658 324832 553664
rect 324688 533520 324740 533526
rect 324688 533462 324740 533468
rect 324792 532574 324820 553658
rect 324780 532568 324832 532574
rect 324780 532510 324832 532516
rect 324884 532234 324912 556310
rect 325148 534608 325200 534614
rect 325036 534556 325148 534562
rect 325036 534550 325200 534556
rect 325036 534534 325188 534550
rect 329544 534126 329788 534154
rect 334052 534126 334112 534154
rect 324872 532228 324924 532234
rect 324872 532170 324924 532176
rect 324596 531820 324648 531826
rect 324596 531762 324648 531768
rect 322480 531140 322532 531146
rect 322480 531082 322532 531088
rect 322204 529508 322256 529514
rect 322204 529450 322256 529456
rect 329760 529446 329788 534126
rect 334084 532574 334112 534126
rect 338224 534126 338560 534154
rect 342732 534126 343068 534154
rect 347240 534126 347576 534154
rect 351932 534126 352084 534154
rect 356256 534126 356592 534154
rect 360764 534126 361100 534154
rect 365272 534126 365608 534154
rect 369872 534126 370116 534154
rect 374288 534126 374624 534154
rect 379532 534126 379776 534154
rect 383672 534126 384284 534154
rect 388456 534126 388792 534154
rect 393300 534126 393360 534154
rect 338224 532710 338252 534126
rect 338212 532704 338264 532710
rect 338212 532646 338264 532652
rect 334072 532568 334124 532574
rect 334072 532510 334124 532516
rect 342732 532409 342760 534126
rect 342718 532400 342774 532409
rect 342718 532335 342774 532344
rect 347240 531962 347268 534126
rect 351932 532030 351960 534126
rect 356256 532914 356284 534126
rect 356244 532908 356296 532914
rect 356244 532850 356296 532856
rect 360764 532545 360792 534126
rect 360750 532536 360806 532545
rect 360750 532471 360806 532480
rect 365272 532166 365300 534126
rect 369872 532302 369900 534126
rect 374288 532846 374316 534126
rect 374276 532840 374328 532846
rect 374276 532782 374328 532788
rect 369860 532296 369912 532302
rect 369860 532238 369912 532244
rect 365260 532160 365312 532166
rect 365260 532102 365312 532108
rect 379532 532098 379560 534126
rect 379520 532092 379572 532098
rect 379520 532034 379572 532040
rect 351920 532024 351972 532030
rect 351920 531966 351972 531972
rect 347228 531956 347280 531962
rect 347228 531898 347280 531904
rect 329748 529440 329800 529446
rect 329748 529382 329800 529388
rect 363604 527876 363656 527882
rect 363604 527818 363656 527824
rect 356980 491224 357032 491230
rect 356980 491166 357032 491172
rect 356796 491088 356848 491094
rect 356796 491030 356848 491036
rect 356704 491020 356756 491026
rect 356704 490962 356756 490968
rect 309784 479528 309836 479534
rect 309784 479470 309836 479476
rect 299756 471912 299808 471918
rect 299756 471854 299808 471860
rect 299296 467764 299348 467770
rect 299296 467706 299348 467712
rect 338488 466608 338540 466614
rect 338486 466576 338488 466585
rect 338540 466576 338542 466585
rect 338486 466511 338542 466520
rect 339774 466576 339830 466585
rect 339774 466511 339776 466520
rect 339828 466511 339830 466520
rect 350998 466576 351054 466585
rect 350998 466511 351054 466520
rect 339776 466482 339828 466488
rect 351012 466478 351040 466511
rect 351000 466472 351052 466478
rect 351000 466414 351052 466420
rect 298374 465896 298430 465905
rect 298374 465831 298430 465840
rect 297088 465588 297140 465594
rect 297088 465530 297140 465536
rect 294420 464500 294472 464506
rect 294420 464442 294472 464448
rect 288716 464432 288768 464438
rect 288716 464374 288768 464380
rect 276848 464364 276900 464370
rect 276848 464306 276900 464312
rect 248236 380928 248288 380934
rect 248236 380870 248288 380876
rect 248248 380769 248276 380870
rect 235998 380760 236054 380769
rect 235998 380695 236054 380704
rect 237102 380760 237158 380769
rect 237102 380695 237158 380704
rect 243082 380760 243138 380769
rect 243082 380695 243138 380704
rect 248234 380760 248290 380769
rect 248234 380695 248290 380704
rect 254490 380760 254546 380769
rect 254490 380695 254546 380704
rect 255870 380760 255926 380769
rect 255870 380695 255926 380704
rect 313462 380760 313518 380769
rect 313462 380695 313518 380704
rect 220726 380352 220782 380361
rect 220726 380287 220782 380296
rect 220740 379409 220768 380287
rect 236012 380050 236040 380695
rect 236000 380044 236052 380050
rect 236000 379986 236052 379992
rect 237116 379914 237144 380695
rect 243096 379982 243124 380695
rect 244278 380488 244334 380497
rect 244278 380423 244334 380432
rect 243084 379976 243136 379982
rect 243084 379918 243136 379924
rect 237104 379908 237156 379914
rect 237104 379850 237156 379856
rect 239772 379908 239824 379914
rect 239772 379850 239824 379856
rect 220082 379400 220138 379409
rect 220726 379400 220782 379409
rect 220082 379335 220138 379344
rect 220452 379364 220504 379370
rect 219990 379128 220046 379137
rect 219990 379063 220046 379072
rect 219900 379024 219952 379030
rect 219900 378966 219952 378972
rect 219992 378684 220044 378690
rect 219992 378626 220044 378632
rect 219808 376644 219860 376650
rect 219808 376586 219860 376592
rect 219808 374944 219860 374950
rect 219808 374886 219860 374892
rect 219820 271794 219848 374886
rect 220004 272490 220032 378626
rect 220096 375698 220124 379335
rect 220726 379335 220782 379344
rect 239586 379400 239642 379409
rect 239586 379335 239642 379344
rect 220452 379306 220504 379312
rect 220464 378622 220492 379306
rect 221004 379296 221056 379302
rect 221004 379238 221056 379244
rect 222016 379296 222068 379302
rect 222016 379238 222068 379244
rect 238206 379264 238262 379273
rect 220820 379092 220872 379098
rect 220820 379034 220872 379040
rect 220728 379024 220780 379030
rect 220728 378966 220780 378972
rect 220636 378820 220688 378826
rect 220636 378762 220688 378768
rect 220648 378690 220676 378762
rect 220636 378684 220688 378690
rect 220636 378626 220688 378632
rect 220452 378616 220504 378622
rect 220740 378593 220768 378966
rect 220452 378558 220504 378564
rect 220726 378584 220782 378593
rect 220726 378519 220782 378528
rect 220084 375692 220136 375698
rect 220084 375634 220136 375640
rect 220636 374944 220688 374950
rect 220636 374886 220688 374892
rect 220648 374746 220676 374886
rect 220636 374740 220688 374746
rect 220636 374682 220688 374688
rect 220832 358766 220860 379034
rect 220910 378720 220966 378729
rect 220910 378655 220966 378664
rect 220820 358760 220872 358766
rect 220820 358702 220872 358708
rect 220924 357678 220952 378655
rect 221016 358290 221044 379238
rect 221464 379160 221516 379166
rect 221464 379102 221516 379108
rect 221476 378690 221504 379102
rect 221096 378684 221148 378690
rect 221096 378626 221148 378632
rect 221464 378684 221516 378690
rect 221464 378626 221516 378632
rect 221108 358494 221136 378626
rect 222028 378622 222056 379238
rect 238206 379199 238262 379208
rect 222108 379092 222160 379098
rect 222108 379034 222160 379040
rect 222016 378616 222068 378622
rect 222016 378558 222068 378564
rect 222120 378554 222148 379034
rect 222108 378548 222160 378554
rect 222108 378490 222160 378496
rect 238220 378350 238248 379199
rect 239600 378418 239628 379335
rect 239588 378412 239640 378418
rect 239588 378354 239640 378360
rect 238208 378344 238260 378350
rect 238208 378286 238260 378292
rect 239784 375834 239812 379850
rect 244292 379846 244320 380423
rect 244280 379840 244332 379846
rect 244280 379782 244332 379788
rect 254504 379778 254532 380695
rect 254492 379772 254544 379778
rect 254492 379714 254544 379720
rect 255884 379710 255912 380695
rect 258078 380624 258134 380633
rect 258078 380559 258134 380568
rect 261758 380624 261814 380633
rect 261758 380559 261814 380568
rect 270958 380624 271014 380633
rect 270958 380559 271014 380568
rect 255872 379704 255924 379710
rect 255872 379646 255924 379652
rect 258092 379642 258120 380559
rect 261772 379914 261800 380559
rect 261760 379908 261812 379914
rect 261760 379850 261812 379856
rect 258080 379636 258132 379642
rect 258080 379578 258132 379584
rect 263876 379568 263928 379574
rect 263876 379510 263928 379516
rect 263888 379409 263916 379510
rect 269764 379432 269816 379438
rect 244922 379400 244978 379409
rect 244922 379335 244978 379344
rect 246210 379400 246266 379409
rect 246210 379335 246266 379344
rect 248602 379400 248658 379409
rect 248602 379335 248658 379344
rect 250074 379400 250130 379409
rect 250074 379335 250130 379344
rect 251178 379400 251234 379409
rect 251178 379335 251234 379344
rect 252282 379400 252338 379409
rect 252282 379335 252338 379344
rect 253386 379400 253442 379409
rect 253386 379335 253442 379344
rect 263874 379400 263930 379409
rect 263874 379335 263930 379344
rect 264978 379400 265034 379409
rect 264978 379335 265034 379344
rect 268290 379400 268346 379409
rect 268290 379335 268346 379344
rect 269762 379400 269764 379409
rect 269816 379400 269818 379409
rect 269762 379335 269818 379344
rect 244936 378486 244964 379335
rect 244924 378480 244976 378486
rect 244924 378422 244976 378428
rect 246224 378282 246252 379335
rect 248616 378826 248644 379335
rect 248604 378820 248656 378826
rect 248604 378762 248656 378768
rect 250088 378758 250116 379335
rect 250626 378856 250682 378865
rect 250626 378791 250682 378800
rect 250076 378752 250128 378758
rect 250076 378694 250128 378700
rect 246212 378276 246264 378282
rect 246212 378218 246264 378224
rect 250640 375970 250668 378791
rect 251192 378690 251220 379335
rect 251180 378684 251232 378690
rect 251180 378626 251232 378632
rect 252296 378622 252324 379335
rect 253202 378856 253258 378865
rect 253202 378791 253258 378800
rect 252284 378616 252336 378622
rect 252284 378558 252336 378564
rect 253216 378457 253244 378791
rect 253400 378554 253428 379335
rect 258354 378584 258410 378593
rect 253388 378548 253440 378554
rect 258354 378519 258410 378528
rect 260562 378584 260618 378593
rect 260562 378519 260618 378528
rect 260930 378584 260986 378593
rect 262770 378584 262826 378593
rect 260930 378519 260986 378528
rect 262220 378548 262272 378554
rect 253388 378490 253440 378496
rect 253202 378448 253258 378457
rect 253202 378383 253258 378392
rect 253386 378448 253442 378457
rect 253386 378383 253442 378392
rect 255962 378448 256018 378457
rect 255962 378383 256018 378392
rect 250628 375964 250680 375970
rect 250628 375906 250680 375912
rect 253400 375902 253428 378383
rect 253388 375896 253440 375902
rect 253388 375838 253440 375844
rect 239772 375828 239824 375834
rect 239772 375770 239824 375776
rect 255976 375766 256004 378383
rect 258368 376174 258396 378519
rect 258356 376168 258408 376174
rect 258356 376110 258408 376116
rect 255964 375760 256016 375766
rect 255964 375702 256016 375708
rect 260576 374882 260604 378519
rect 260944 376242 260972 378519
rect 262770 378519 262826 378528
rect 263598 378584 263654 378593
rect 263598 378519 263654 378528
rect 262220 378490 262272 378496
rect 260932 376236 260984 376242
rect 260932 376178 260984 376184
rect 260564 374876 260616 374882
rect 260564 374818 260616 374824
rect 262232 374814 262260 378490
rect 262784 375358 262812 378519
rect 263612 376378 263640 378519
rect 263876 378276 263928 378282
rect 263876 378218 263928 378224
rect 263600 376372 263652 376378
rect 263600 376314 263652 376320
rect 262772 375352 262824 375358
rect 262772 375294 262824 375300
rect 263888 375290 263916 378218
rect 264992 377262 265020 379335
rect 268304 378894 268332 379335
rect 266452 378888 266504 378894
rect 266452 378830 266504 378836
rect 268292 378888 268344 378894
rect 268292 378830 268344 378836
rect 265898 378584 265954 378593
rect 265898 378519 265954 378528
rect 266358 378584 266414 378593
rect 266358 378519 266360 378528
rect 264980 377256 265032 377262
rect 264980 377198 265032 377204
rect 265912 376106 265940 378519
rect 266412 378519 266414 378528
rect 266360 378490 266412 378496
rect 265900 376100 265952 376106
rect 265900 376042 265952 376048
rect 263876 375284 263928 375290
rect 263876 375226 263928 375232
rect 262220 374808 262272 374814
rect 262220 374750 262272 374756
rect 266464 374746 266492 378830
rect 267554 378584 267610 378593
rect 267554 378519 267610 378528
rect 268014 378584 268070 378593
rect 268014 378519 268070 378528
rect 267568 378282 267596 378519
rect 267556 378276 267608 378282
rect 267556 378218 267608 378224
rect 268028 376310 268056 378519
rect 270972 377330 271000 380559
rect 291844 380384 291896 380390
rect 291844 380326 291896 380332
rect 291856 379506 291884 380326
rect 298008 380316 298060 380322
rect 298008 380258 298060 380264
rect 273260 379500 273312 379506
rect 273260 379442 273312 379448
rect 291844 379500 291896 379506
rect 291844 379442 291896 379448
rect 273272 379409 273300 379442
rect 298020 379438 298048 380258
rect 313476 380254 313504 380695
rect 315854 380624 315910 380633
rect 315854 380559 315910 380568
rect 313464 380248 313516 380254
rect 313464 380190 313516 380196
rect 315868 380186 315896 380559
rect 315856 380180 315908 380186
rect 315856 380122 315908 380128
rect 320916 379500 320968 379506
rect 320916 379442 320968 379448
rect 298008 379432 298060 379438
rect 271050 379400 271106 379409
rect 271050 379335 271052 379344
rect 271104 379335 271106 379344
rect 272154 379400 272210 379409
rect 272154 379335 272210 379344
rect 273258 379400 273314 379409
rect 273258 379335 273314 379344
rect 275742 379400 275798 379409
rect 275742 379335 275798 379344
rect 285954 379400 286010 379409
rect 285954 379335 286010 379344
rect 287702 379400 287758 379409
rect 287702 379335 287758 379344
rect 290186 379400 290242 379409
rect 290186 379335 290242 379344
rect 293314 379400 293370 379409
rect 293314 379335 293370 379344
rect 295890 379400 295946 379409
rect 305828 379432 305880 379438
rect 298008 379374 298060 379380
rect 298098 379400 298154 379409
rect 295890 379335 295946 379344
rect 298098 379335 298154 379344
rect 305826 379400 305828 379409
rect 320928 379409 320956 379442
rect 305880 379400 305882 379409
rect 305826 379335 305882 379344
rect 307850 379400 307906 379409
rect 307850 379335 307906 379344
rect 310978 379400 311034 379409
rect 310978 379335 311034 379344
rect 317786 379400 317842 379409
rect 317786 379335 317842 379344
rect 320914 379400 320970 379409
rect 320914 379335 320970 379344
rect 325882 379400 325938 379409
rect 325882 379335 325938 379344
rect 271052 379306 271104 379312
rect 272168 378214 272196 379335
rect 273442 378992 273498 379001
rect 273442 378927 273498 378936
rect 272156 378208 272208 378214
rect 272156 378150 272208 378156
rect 273260 378208 273312 378214
rect 273260 378150 273312 378156
rect 273272 377874 273300 378150
rect 273260 377868 273312 377874
rect 273260 377810 273312 377816
rect 270960 377324 271012 377330
rect 270960 377266 271012 377272
rect 273456 376446 273484 378927
rect 274638 378448 274694 378457
rect 274638 378383 274694 378392
rect 274652 378282 274680 378383
rect 275756 378282 275784 379335
rect 276110 379264 276166 379273
rect 276110 379199 276166 379208
rect 277030 379264 277086 379273
rect 277030 379199 277086 379208
rect 278410 379264 278466 379273
rect 278410 379199 278466 379208
rect 280802 379264 280858 379273
rect 280802 379199 280858 379208
rect 283102 379264 283158 379273
rect 283102 379199 283158 379208
rect 276020 378480 276072 378486
rect 276020 378422 276072 378428
rect 276032 378321 276060 378422
rect 276018 378312 276074 378321
rect 274640 378276 274692 378282
rect 274640 378218 274692 378224
rect 275744 378276 275796 378282
rect 276018 378247 276074 378256
rect 275744 378218 275796 378224
rect 276124 376582 276152 379199
rect 277044 378486 277072 379199
rect 277306 378992 277362 379001
rect 277306 378927 277362 378936
rect 277032 378480 277084 378486
rect 277032 378422 277084 378428
rect 276112 376576 276164 376582
rect 276112 376518 276164 376524
rect 273444 376440 273496 376446
rect 273444 376382 273496 376388
rect 268016 376304 268068 376310
rect 268016 376246 268068 376252
rect 266452 374740 266504 374746
rect 266452 374682 266504 374688
rect 277320 359582 277348 378927
rect 278424 377398 278452 379199
rect 280068 378548 280120 378554
rect 280068 378490 280120 378496
rect 280080 378185 280108 378490
rect 280066 378176 280122 378185
rect 280066 378111 280122 378120
rect 280816 377466 280844 379199
rect 280804 377460 280856 377466
rect 280804 377402 280856 377408
rect 278412 377392 278464 377398
rect 278412 377334 278464 377340
rect 283116 376514 283144 379199
rect 285968 378214 285996 379335
rect 285956 378208 286008 378214
rect 285956 378150 286008 378156
rect 287716 377534 287744 379335
rect 290200 377602 290228 379335
rect 293328 377670 293356 379335
rect 295904 377738 295932 379335
rect 298112 377806 298140 379335
rect 300858 379264 300914 379273
rect 300858 379199 300914 379208
rect 298100 377800 298152 377806
rect 298100 377742 298152 377748
rect 295892 377732 295944 377738
rect 295892 377674 295944 377680
rect 293316 377664 293368 377670
rect 293316 377606 293368 377612
rect 290188 377596 290240 377602
rect 290188 377538 290240 377544
rect 287704 377528 287756 377534
rect 287704 377470 287756 377476
rect 300872 376718 300900 379199
rect 302514 378992 302570 379001
rect 302514 378927 302570 378936
rect 300860 376712 300912 376718
rect 300860 376654 300912 376660
rect 302528 376650 302556 378927
rect 307864 377942 307892 379335
rect 310992 378146 311020 379335
rect 310980 378140 311032 378146
rect 310980 378082 311032 378088
rect 317800 378010 317828 379335
rect 325896 378078 325924 379335
rect 343454 379128 343510 379137
rect 343454 379063 343510 379072
rect 343468 378622 343496 379063
rect 343546 378992 343602 379001
rect 343546 378927 343602 378936
rect 343560 378758 343588 378927
rect 343548 378752 343600 378758
rect 343548 378694 343600 378700
rect 342904 378616 342956 378622
rect 342904 378558 342956 378564
rect 343456 378616 343508 378622
rect 343456 378558 343508 378564
rect 325884 378072 325936 378078
rect 325884 378014 325936 378020
rect 317788 378004 317840 378010
rect 317788 377946 317840 377952
rect 307852 377936 307904 377942
rect 307852 377878 307904 377884
rect 302516 376644 302568 376650
rect 302516 376586 302568 376592
rect 283104 376508 283156 376514
rect 283104 376450 283156 376456
rect 342916 367810 342944 378558
rect 342904 367804 342956 367810
rect 342904 367746 342956 367752
rect 277308 359576 277360 359582
rect 277308 359518 277360 359524
rect 343560 358970 343588 378694
rect 356612 378276 356664 378282
rect 356612 378218 356664 378224
rect 351736 359508 351788 359514
rect 351736 359450 351788 359456
rect 342260 358964 342312 358970
rect 342260 358906 342312 358912
rect 343548 358964 343600 358970
rect 343548 358906 343600 358912
rect 339776 358896 339828 358902
rect 338486 358864 338542 358873
rect 338486 358799 338488 358808
rect 338540 358799 338542 358808
rect 339774 358864 339776 358873
rect 339828 358864 339830 358873
rect 339774 358799 339830 358808
rect 338488 358770 338540 358776
rect 221096 358488 221148 358494
rect 221096 358430 221148 358436
rect 221004 358284 221056 358290
rect 221004 358226 221056 358232
rect 342272 358086 342300 358906
rect 351748 358873 351776 359450
rect 351734 358864 351790 358873
rect 351734 358799 351790 358808
rect 342260 358080 342312 358086
rect 342260 358022 342312 358028
rect 220912 357672 220964 357678
rect 220912 357614 220964 357620
rect 250718 273592 250774 273601
rect 250718 273527 250774 273536
rect 272246 273592 272302 273601
rect 272246 273527 272302 273536
rect 280894 273592 280950 273601
rect 280894 273527 280950 273536
rect 250732 273494 250760 273527
rect 250720 273488 250772 273494
rect 250720 273430 250772 273436
rect 272260 273426 272288 273527
rect 273258 273456 273314 273465
rect 272248 273420 272300 273426
rect 273258 273391 273314 273400
rect 272248 273362 272300 273368
rect 273272 273358 273300 273391
rect 273260 273352 273312 273358
rect 273260 273294 273312 273300
rect 280908 273290 280936 273527
rect 280896 273284 280948 273290
rect 280896 273226 280948 273232
rect 283380 272876 283432 272882
rect 283380 272818 283432 272824
rect 283392 272785 283420 272818
rect 295892 272808 295944 272814
rect 283378 272776 283434 272785
rect 283378 272711 283434 272720
rect 288162 272776 288218 272785
rect 288162 272711 288218 272720
rect 290922 272776 290978 272785
rect 290922 272711 290924 272720
rect 288176 272678 288204 272711
rect 290976 272711 290978 272720
rect 295890 272776 295892 272785
rect 295944 272776 295946 272785
rect 295890 272711 295946 272720
rect 290924 272682 290976 272688
rect 288164 272672 288216 272678
rect 288164 272614 288216 272620
rect 298466 272640 298522 272649
rect 298466 272575 298468 272584
rect 298520 272575 298522 272584
rect 300858 272640 300914 272649
rect 300858 272575 300914 272584
rect 298468 272546 298520 272552
rect 300872 272542 300900 272575
rect 300860 272536 300912 272542
rect 220004 272462 220216 272490
rect 300860 272478 300912 272484
rect 219808 271788 219860 271794
rect 219808 271730 219860 271736
rect 220188 270298 220216 272462
rect 235998 272232 236054 272241
rect 235998 272167 236054 272176
rect 236012 271930 236040 272167
rect 236000 271924 236052 271930
rect 236000 271866 236052 271872
rect 307760 271856 307812 271862
rect 255318 271824 255374 271833
rect 223580 271788 223632 271794
rect 255318 271759 255374 271768
rect 263598 271824 263654 271833
rect 263598 271759 263654 271768
rect 264978 271824 265034 271833
rect 264978 271759 265034 271768
rect 268014 271824 268070 271833
rect 268014 271759 268070 271768
rect 270498 271824 270554 271833
rect 270498 271759 270554 271768
rect 273258 271824 273314 271833
rect 273258 271759 273314 271768
rect 275926 271824 275982 271833
rect 275926 271759 275982 271768
rect 276110 271824 276166 271833
rect 276110 271759 276166 271768
rect 277214 271824 277270 271833
rect 277214 271759 277270 271768
rect 278686 271824 278742 271833
rect 278686 271759 278742 271768
rect 302238 271824 302294 271833
rect 302238 271759 302240 271768
rect 223580 271730 223632 271736
rect 223592 271386 223620 271730
rect 223580 271380 223632 271386
rect 223580 271322 223632 271328
rect 224224 271380 224276 271386
rect 224224 271322 224276 271328
rect 224236 270910 224264 271322
rect 255332 271318 255360 271759
rect 263612 271590 263640 271759
rect 264992 271658 265020 271759
rect 264980 271652 265032 271658
rect 264980 271594 265032 271600
rect 263600 271584 263652 271590
rect 263600 271526 263652 271532
rect 268028 271386 268056 271759
rect 270512 271726 270540 271759
rect 270500 271720 270552 271726
rect 270500 271662 270552 271668
rect 273272 271454 273300 271759
rect 273260 271448 273312 271454
rect 273260 271390 273312 271396
rect 268016 271380 268068 271386
rect 268016 271322 268068 271328
rect 255320 271312 255372 271318
rect 255320 271254 255372 271260
rect 258262 271280 258318 271289
rect 258262 271215 258318 271224
rect 260838 271280 260894 271289
rect 260838 271215 260840 271224
rect 258276 271182 258304 271215
rect 260892 271215 260894 271224
rect 260840 271186 260892 271192
rect 275940 271182 275968 271759
rect 276124 271522 276152 271759
rect 276112 271516 276164 271522
rect 276112 271458 276164 271464
rect 277228 271318 277256 271759
rect 278700 271386 278728 271759
rect 302292 271759 302294 271768
rect 307758 271824 307760 271833
rect 307812 271824 307814 271833
rect 307758 271759 307814 271768
rect 302240 271730 302292 271736
rect 343546 271688 343602 271697
rect 343546 271623 343602 271632
rect 343560 271590 343588 271623
rect 343548 271584 343600 271590
rect 343454 271552 343510 271561
rect 343548 271526 343600 271532
rect 343454 271487 343510 271496
rect 343468 271454 343496 271487
rect 343456 271448 343508 271454
rect 343456 271390 343508 271396
rect 278688 271380 278740 271386
rect 278688 271322 278740 271328
rect 277216 271312 277268 271318
rect 277216 271254 277268 271260
rect 280066 271280 280122 271289
rect 280066 271215 280068 271224
rect 280120 271215 280122 271224
rect 280068 271186 280120 271192
rect 258264 271176 258316 271182
rect 239126 271144 239182 271153
rect 239126 271079 239182 271088
rect 247038 271144 247094 271153
rect 247038 271079 247094 271088
rect 252558 271144 252614 271153
rect 275928 271176 275980 271182
rect 258264 271118 258316 271124
rect 260838 271144 260894 271153
rect 252558 271079 252614 271088
rect 260838 271079 260894 271088
rect 266358 271144 266414 271153
rect 266358 271079 266414 271088
rect 268106 271144 268162 271153
rect 268106 271079 268108 271088
rect 224224 270904 224276 270910
rect 224224 270846 224276 270852
rect 235998 270600 236054 270609
rect 235998 270535 236054 270544
rect 237378 270600 237434 270609
rect 237378 270535 237434 270544
rect 224224 270496 224276 270502
rect 224224 270438 224276 270444
rect 220452 270360 220504 270366
rect 220452 270302 220504 270308
rect 220176 270292 220228 270298
rect 220176 270234 220228 270240
rect 219900 270224 219952 270230
rect 219900 270166 219952 270172
rect 219808 269272 219860 269278
rect 219808 269214 219860 269220
rect 219716 268932 219768 268938
rect 219716 268874 219768 268880
rect 219622 167104 219678 167113
rect 219622 167039 219678 167048
rect 219532 164212 219584 164218
rect 219532 164154 219584 164160
rect 219532 162988 219584 162994
rect 219532 162930 219584 162936
rect 219440 156528 219492 156534
rect 219440 156470 219492 156476
rect 219440 156392 219492 156398
rect 219440 156334 219492 156340
rect 219452 59226 219480 156334
rect 219440 59220 219492 59226
rect 219440 59162 219492 59168
rect 219348 58812 219400 58818
rect 219348 58754 219400 58760
rect 219346 58576 219402 58585
rect 219346 58511 219402 58520
rect 219360 58002 219388 58511
rect 219348 57996 219400 58002
rect 219348 57938 219400 57944
rect 219544 56234 219572 162930
rect 219636 58750 219664 167039
rect 219728 146266 219756 268874
rect 219820 156670 219848 269214
rect 219808 156664 219860 156670
rect 219808 156606 219860 156612
rect 219808 156528 219860 156534
rect 219808 156470 219860 156476
rect 219716 146260 219768 146266
rect 219716 146202 219768 146208
rect 219624 58744 219676 58750
rect 219624 58686 219676 58692
rect 219532 56228 219584 56234
rect 219532 56170 219584 56176
rect 219256 55072 219308 55078
rect 219256 55014 219308 55020
rect 219728 55010 219756 146202
rect 219820 146198 219848 156470
rect 219808 146192 219860 146198
rect 219808 146134 219860 146140
rect 219820 145042 219848 146134
rect 219912 145926 219940 270166
rect 220188 269210 220216 270234
rect 220176 269204 220228 269210
rect 220176 269146 220228 269152
rect 220464 269142 220492 270302
rect 220544 270088 220596 270094
rect 220544 270030 220596 270036
rect 220636 270088 220688 270094
rect 220636 270030 220688 270036
rect 220556 269618 220584 270030
rect 220544 269612 220596 269618
rect 220544 269554 220596 269560
rect 220648 269278 220676 270030
rect 220728 270020 220780 270026
rect 220728 269962 220780 269968
rect 220740 269346 220768 269962
rect 224236 269550 224264 270438
rect 224224 269544 224276 269550
rect 224224 269486 224276 269492
rect 220728 269340 220780 269346
rect 220728 269282 220780 269288
rect 220636 269272 220688 269278
rect 220636 269214 220688 269220
rect 220452 269136 220504 269142
rect 220452 269078 220504 269084
rect 236012 268734 236040 270535
rect 237392 269686 237420 270535
rect 239140 270162 239168 271079
rect 247052 270978 247080 271079
rect 252572 271046 252600 271079
rect 252560 271040 252612 271046
rect 252560 270982 252612 270988
rect 247040 270972 247092 270978
rect 247040 270914 247092 270920
rect 252558 270872 252614 270881
rect 252558 270807 252614 270816
rect 244278 270736 244334 270745
rect 244278 270671 244334 270680
rect 251270 270736 251326 270745
rect 251270 270671 251326 270680
rect 242898 270600 242954 270609
rect 242898 270535 242954 270544
rect 239128 270156 239180 270162
rect 239128 270098 239180 270104
rect 237380 269680 237432 269686
rect 237380 269622 237432 269628
rect 242912 268802 242940 270535
rect 244292 270434 244320 270671
rect 244370 270600 244426 270609
rect 244370 270535 244426 270544
rect 245658 270600 245714 270609
rect 245658 270535 245714 270544
rect 247038 270600 247094 270609
rect 247038 270535 247094 270544
rect 248510 270600 248566 270609
rect 248510 270535 248566 270544
rect 249798 270600 249854 270609
rect 249798 270535 249854 270544
rect 251178 270600 251234 270609
rect 251178 270535 251234 270544
rect 244280 270428 244332 270434
rect 244280 270370 244332 270376
rect 244384 268870 244412 270535
rect 245672 269754 245700 270535
rect 245660 269748 245712 269754
rect 245660 269690 245712 269696
rect 247052 269618 247080 270535
rect 248524 270298 248552 270535
rect 249812 270366 249840 270535
rect 249800 270360 249852 270366
rect 249800 270302 249852 270308
rect 248512 270292 248564 270298
rect 248512 270234 248564 270240
rect 251192 270094 251220 270535
rect 251284 270230 251312 270671
rect 251272 270224 251324 270230
rect 251272 270166 251324 270172
rect 251180 270088 251232 270094
rect 251180 270030 251232 270036
rect 252572 270026 252600 270807
rect 259550 270736 259606 270745
rect 259550 270671 259606 270680
rect 253938 270600 253994 270609
rect 253938 270535 253994 270544
rect 255318 270600 255374 270609
rect 255318 270535 255374 270544
rect 256698 270600 256754 270609
rect 256698 270535 256754 270544
rect 258078 270600 258134 270609
rect 258078 270535 258134 270544
rect 259458 270600 259514 270609
rect 259458 270535 259514 270544
rect 252560 270020 252612 270026
rect 252560 269962 252612 269968
rect 247040 269612 247092 269618
rect 247040 269554 247092 269560
rect 253952 268938 253980 270535
rect 255332 269006 255360 270535
rect 256712 269074 256740 270535
rect 256700 269068 256752 269074
rect 256700 269010 256752 269016
rect 255320 269000 255372 269006
rect 255320 268942 255372 268948
rect 253940 268932 253992 268938
rect 253940 268874 253992 268880
rect 244372 268864 244424 268870
rect 244372 268806 244424 268812
rect 242900 268796 242952 268802
rect 242900 268738 242952 268744
rect 236000 268728 236052 268734
rect 236000 268670 236052 268676
rect 258092 268666 258120 270535
rect 233240 268660 233292 268666
rect 233240 268602 233292 268608
rect 258080 268660 258132 268666
rect 258080 268602 258132 268608
rect 231860 268592 231912 268598
rect 231860 268534 231912 268540
rect 230480 268524 230532 268530
rect 230480 268466 230532 268472
rect 230388 268456 230440 268462
rect 229098 268424 229154 268433
rect 229098 268359 229154 268368
rect 230386 268424 230388 268433
rect 230440 268424 230442 268433
rect 230386 268359 230442 268368
rect 229112 252074 229140 268359
rect 229100 252068 229152 252074
rect 229100 252010 229152 252016
rect 230492 252006 230520 268466
rect 230480 252000 230532 252006
rect 230480 251942 230532 251948
rect 231872 251841 231900 268534
rect 233252 251938 233280 268602
rect 259472 268598 259500 270535
rect 259460 268592 259512 268598
rect 259460 268534 259512 268540
rect 259564 268530 259592 270671
rect 259552 268524 259604 268530
rect 259552 268466 259604 268472
rect 260852 268462 260880 271079
rect 266372 270910 266400 271079
rect 268160 271079 268162 271088
rect 270498 271144 270554 271153
rect 275928 271118 275980 271124
rect 270498 271079 270554 271088
rect 268108 271050 268160 271056
rect 264244 270904 264296 270910
rect 266360 270904 266412 270910
rect 264244 270846 264296 270852
rect 264978 270872 265034 270881
rect 262218 270600 262274 270609
rect 262218 270535 262274 270544
rect 263598 270600 263654 270609
rect 263598 270535 263654 270544
rect 262232 270502 262260 270535
rect 262220 270496 262272 270502
rect 262220 270438 262272 270444
rect 263612 269958 263640 270535
rect 263600 269952 263652 269958
rect 263600 269894 263652 269900
rect 260840 268456 260892 268462
rect 260840 268398 260892 268404
rect 233240 251932 233292 251938
rect 233240 251874 233292 251880
rect 264256 251870 264284 270846
rect 266360 270846 266412 270852
rect 264978 270807 265034 270816
rect 264992 252482 265020 270807
rect 265622 270736 265678 270745
rect 265622 270671 265678 270680
rect 265636 252550 265664 270671
rect 269118 270600 269174 270609
rect 268844 270564 268896 270570
rect 269118 270535 269174 270544
rect 268844 270506 268896 270512
rect 268856 268394 268884 270506
rect 269132 269890 269160 270535
rect 269120 269884 269172 269890
rect 269120 269826 269172 269832
rect 270512 269822 270540 271079
rect 273258 270600 273314 270609
rect 273258 270535 273260 270544
rect 273312 270535 273314 270544
rect 273260 270506 273312 270512
rect 270500 269816 270552 269822
rect 270500 269758 270552 269764
rect 268844 268388 268896 268394
rect 268844 268330 268896 268336
rect 343468 267734 343496 271390
rect 356624 271182 356652 378218
rect 356612 271176 356664 271182
rect 356612 271118 356664 271124
rect 343468 267706 343588 267734
rect 340788 253904 340840 253910
rect 340788 253846 340840 253852
rect 340800 253473 340828 253846
rect 340786 253464 340842 253473
rect 340786 253399 340842 253408
rect 339408 253292 339460 253298
rect 339408 253234 339460 253240
rect 339420 253065 339448 253234
rect 339406 253056 339462 253065
rect 339406 252991 339462 253000
rect 265624 252544 265676 252550
rect 265624 252486 265676 252492
rect 264980 252476 265032 252482
rect 264980 252418 265032 252424
rect 343560 251870 343588 267706
rect 351828 253224 351880 253230
rect 351826 253192 351828 253201
rect 351880 253192 351882 253201
rect 351826 253127 351882 253136
rect 264244 251864 264296 251870
rect 231858 251832 231914 251841
rect 264244 251806 264296 251812
rect 343548 251864 343600 251870
rect 343548 251806 343600 251812
rect 231858 251767 231914 251776
rect 356716 166870 356744 490962
rect 253572 166864 253624 166870
rect 356704 166864 356756 166870
rect 253572 166806 253624 166812
rect 298466 166832 298522 166841
rect 253584 166569 253612 166806
rect 270868 166796 270920 166802
rect 298466 166767 298522 166776
rect 303526 166832 303582 166841
rect 356704 166806 356756 166812
rect 356808 166802 356836 491030
rect 356888 478440 356940 478446
rect 356888 478382 356940 478388
rect 356900 272950 356928 478382
rect 356992 380798 357020 491166
rect 361120 491156 361172 491162
rect 361120 491098 361172 491104
rect 358268 490952 358320 490958
rect 358268 490894 358320 490900
rect 358176 490748 358228 490754
rect 358176 490690 358228 490696
rect 357072 484288 357124 484294
rect 357072 484230 357124 484236
rect 356980 380792 357032 380798
rect 356980 380734 357032 380740
rect 356980 378480 357032 378486
rect 356980 378422 357032 378428
rect 356992 287054 357020 378422
rect 357084 376310 357112 484230
rect 357992 481500 358044 481506
rect 357992 481442 358044 481448
rect 357164 478712 357216 478718
rect 357164 478654 357216 478660
rect 357176 376718 357204 478654
rect 357256 469804 357308 469810
rect 357256 469746 357308 469752
rect 357164 376712 357216 376718
rect 357164 376654 357216 376660
rect 357072 376304 357124 376310
rect 357072 376246 357124 376252
rect 357268 374814 357296 469746
rect 357900 464364 357952 464370
rect 357900 464306 357952 464312
rect 357912 377942 357940 464306
rect 358004 380662 358032 481442
rect 358084 475788 358136 475794
rect 358084 475730 358136 475736
rect 358096 417450 358124 475730
rect 358084 417444 358136 417450
rect 358084 417386 358136 417392
rect 358084 389224 358136 389230
rect 358084 389166 358136 389172
rect 357992 380656 358044 380662
rect 357992 380598 358044 380604
rect 357900 377936 357952 377942
rect 357900 377878 357952 377884
rect 357256 374808 357308 374814
rect 357256 374750 357308 374756
rect 357440 359576 357492 359582
rect 357440 359518 357492 359524
rect 357348 358896 357400 358902
rect 357348 358838 357400 358844
rect 356992 287026 357204 287054
rect 356888 272944 356940 272950
rect 356888 272886 356940 272892
rect 357072 271584 357124 271590
rect 357072 271526 357124 271532
rect 356888 271176 356940 271182
rect 356888 271118 356940 271124
rect 303526 166767 303582 166776
rect 356796 166796 356848 166802
rect 270868 166738 270920 166744
rect 265900 166728 265952 166734
rect 265900 166670 265952 166676
rect 265912 166569 265940 166670
rect 270880 166569 270908 166738
rect 288254 166696 288310 166705
rect 288254 166631 288256 166640
rect 288308 166631 288310 166640
rect 295890 166696 295946 166705
rect 295890 166631 295946 166640
rect 288256 166602 288308 166608
rect 253570 166560 253626 166569
rect 253570 166495 253626 166504
rect 265898 166560 265954 166569
rect 265898 166495 265954 166504
rect 270866 166560 270922 166569
rect 270866 166495 270922 166504
rect 295904 166462 295932 166631
rect 298480 166598 298508 166767
rect 298468 166592 298520 166598
rect 298468 166534 298520 166540
rect 303540 166530 303568 166767
rect 356796 166738 356848 166744
rect 308494 166696 308550 166705
rect 308494 166631 308550 166640
rect 315854 166696 315910 166705
rect 315854 166631 315910 166640
rect 303528 166524 303580 166530
rect 303528 166466 303580 166472
rect 295892 166456 295944 166462
rect 295892 166398 295944 166404
rect 308508 166394 308536 166631
rect 308496 166388 308548 166394
rect 308496 166330 308548 166336
rect 315868 166326 315896 166631
rect 315856 166320 315908 166326
rect 315856 166262 315908 166268
rect 236090 165608 236146 165617
rect 236090 165543 236146 165552
rect 238758 165608 238814 165617
rect 238758 165543 238814 165552
rect 242898 165608 242954 165617
rect 242898 165543 242954 165552
rect 247130 165608 247186 165617
rect 247130 165543 247186 165552
rect 258170 165608 258226 165617
rect 258170 165543 258226 165552
rect 260838 165608 260894 165617
rect 260838 165543 260894 165552
rect 273442 165608 273498 165617
rect 273442 165543 273498 165552
rect 276018 165608 276074 165617
rect 276018 165543 276074 165552
rect 278410 165608 278466 165617
rect 278410 165543 278466 165552
rect 280802 165608 280858 165617
rect 280802 165543 280858 165552
rect 285954 165608 286010 165617
rect 285954 165543 286010 165552
rect 293314 165608 293370 165617
rect 293314 165543 293370 165552
rect 300858 165608 300914 165617
rect 300858 165543 300914 165552
rect 310978 165608 311034 165617
rect 310978 165543 310980 165552
rect 235998 164248 236054 164257
rect 219992 164212 220044 164218
rect 235998 164183 236054 164192
rect 219992 164154 220044 164160
rect 219900 145920 219952 145926
rect 219900 145862 219952 145868
rect 219808 145036 219860 145042
rect 219808 144978 219860 144984
rect 219912 144974 219940 145862
rect 219900 144968 219952 144974
rect 219900 144910 219952 144916
rect 220004 56302 220032 164154
rect 220728 163600 220780 163606
rect 220728 163542 220780 163548
rect 220740 162994 220768 163542
rect 220728 162988 220780 162994
rect 220728 162930 220780 162936
rect 220176 162172 220228 162178
rect 220176 162114 220228 162120
rect 220188 161430 220216 162114
rect 235264 161492 235316 161498
rect 235264 161434 235316 161440
rect 220176 161424 220228 161430
rect 220176 161366 220228 161372
rect 220084 156664 220136 156670
rect 220084 156606 220136 156612
rect 220096 145994 220124 156606
rect 220188 156398 220216 161366
rect 220176 156392 220228 156398
rect 220176 156334 220228 156340
rect 235276 146198 235304 161434
rect 235264 146192 235316 146198
rect 235264 146134 235316 146140
rect 220084 145988 220136 145994
rect 220084 145930 220136 145936
rect 220096 145110 220124 145930
rect 236012 145518 236040 164183
rect 236000 145512 236052 145518
rect 236000 145454 236052 145460
rect 236104 145450 236132 165543
rect 237378 164248 237434 164257
rect 237378 164183 237434 164192
rect 237392 145897 237420 164183
rect 238772 148510 238800 165543
rect 240138 164248 240194 164257
rect 240138 164183 240194 164192
rect 241518 164248 241574 164257
rect 241518 164183 241574 164192
rect 240152 148918 240180 164183
rect 240140 148912 240192 148918
rect 240140 148854 240192 148860
rect 238760 148504 238812 148510
rect 238760 148446 238812 148452
rect 241532 148442 241560 164183
rect 241520 148436 241572 148442
rect 241520 148378 241572 148384
rect 237378 145888 237434 145897
rect 237378 145823 237434 145832
rect 242912 145722 242940 165543
rect 247038 164928 247094 164937
rect 247038 164863 247094 164872
rect 247052 164694 247080 164863
rect 247040 164688 247092 164694
rect 247040 164630 247092 164636
rect 244370 164384 244426 164393
rect 244370 164319 244426 164328
rect 244278 164248 244334 164257
rect 244278 164183 244334 164192
rect 242900 145716 242952 145722
rect 242900 145658 242952 145664
rect 244292 145586 244320 164183
rect 244384 145654 244412 164319
rect 245658 164248 245714 164257
rect 245658 164183 245714 164192
rect 245672 145790 245700 164183
rect 245660 145784 245712 145790
rect 245660 145726 245712 145732
rect 244372 145648 244424 145654
rect 244372 145590 244424 145596
rect 244280 145580 244332 145586
rect 244280 145522 244332 145528
rect 236092 145444 236144 145450
rect 236092 145386 236144 145392
rect 247144 145382 247172 165543
rect 249798 164928 249854 164937
rect 249798 164863 249854 164872
rect 255318 164928 255374 164937
rect 255318 164863 255374 164872
rect 258078 164928 258134 164937
rect 258078 164863 258080 164872
rect 249812 164762 249840 164863
rect 255332 164830 255360 164863
rect 258132 164863 258134 164872
rect 258080 164834 258132 164840
rect 255320 164824 255372 164830
rect 255320 164766 255372 164772
rect 249800 164756 249852 164762
rect 249800 164698 249852 164704
rect 251270 164384 251326 164393
rect 251270 164319 251326 164328
rect 256698 164384 256754 164393
rect 256698 164319 256754 164328
rect 248418 164248 248474 164257
rect 248418 164183 248474 164192
rect 249890 164248 249946 164257
rect 249890 164183 249946 164192
rect 251178 164248 251234 164257
rect 251178 164183 251234 164192
rect 248432 146062 248460 164183
rect 248420 146056 248472 146062
rect 248420 145998 248472 146004
rect 249904 145858 249932 164183
rect 251192 145994 251220 164183
rect 251180 145988 251232 145994
rect 251180 145930 251232 145936
rect 251284 145926 251312 164319
rect 252558 164248 252614 164257
rect 252558 164183 252614 164192
rect 253938 164248 253994 164257
rect 253938 164183 253994 164192
rect 255410 164248 255466 164257
rect 255410 164183 255466 164192
rect 252572 146130 252600 164183
rect 253952 146266 253980 164183
rect 253940 146260 253992 146266
rect 253940 146202 253992 146208
rect 255424 146198 255452 164183
rect 256712 162178 256740 164319
rect 258184 162654 258212 165543
rect 259550 164384 259606 164393
rect 259550 164319 259606 164328
rect 259458 164248 259514 164257
rect 259458 164183 259514 164192
rect 259472 162722 259500 164183
rect 259564 162790 259592 164319
rect 260852 162858 260880 165543
rect 263598 165200 263654 165209
rect 263598 165135 263654 165144
rect 266266 165200 266322 165209
rect 271878 165200 271934 165209
rect 266322 165158 266400 165186
rect 266266 165135 266322 165144
rect 263612 165102 263640 165135
rect 263600 165096 263652 165102
rect 263600 165038 263652 165044
rect 262218 164248 262274 164257
rect 262218 164183 262274 164192
rect 263782 164248 263838 164257
rect 263782 164183 263838 164192
rect 262232 163674 262260 164183
rect 263796 163742 263824 164183
rect 263784 163736 263836 163742
rect 263784 163678 263836 163684
rect 262220 163668 262272 163674
rect 262220 163610 262272 163616
rect 260840 162852 260892 162858
rect 260840 162794 260892 162800
rect 259552 162784 259604 162790
rect 259552 162726 259604 162732
rect 259460 162716 259512 162722
rect 259460 162658 259512 162664
rect 258172 162648 258224 162654
rect 258172 162590 258224 162596
rect 256700 162172 256752 162178
rect 256700 162114 256752 162120
rect 266372 157334 266400 165158
rect 271878 165135 271934 165144
rect 267738 165064 267794 165073
rect 267738 164999 267794 165008
rect 267752 164966 267780 164999
rect 267740 164960 267792 164966
rect 267740 164902 267792 164908
rect 266542 164384 266598 164393
rect 266542 164319 266598 164328
rect 266450 164248 266506 164257
rect 266450 164183 266506 164192
rect 266464 163606 266492 164183
rect 266452 163600 266504 163606
rect 266452 163542 266504 163548
rect 266556 163538 266584 164319
rect 269764 164280 269816 164286
rect 267738 164248 267794 164257
rect 267738 164183 267740 164192
rect 267792 164183 267794 164192
rect 269118 164248 269174 164257
rect 269764 164222 269816 164228
rect 270498 164248 270554 164257
rect 269118 164183 269174 164192
rect 267740 164154 267792 164160
rect 266544 163532 266596 163538
rect 266544 163474 266596 163480
rect 266372 157306 266584 157334
rect 255412 146192 255464 146198
rect 266556 146169 266584 157306
rect 269132 146305 269160 164183
rect 269776 148986 269804 164222
rect 270498 164183 270554 164192
rect 269764 148980 269816 148986
rect 269764 148922 269816 148928
rect 269118 146296 269174 146305
rect 269118 146231 269174 146240
rect 255412 146134 255464 146140
rect 266542 146160 266598 146169
rect 252560 146124 252612 146130
rect 266542 146095 266598 146104
rect 252560 146066 252612 146072
rect 251272 145920 251324 145926
rect 251272 145862 251324 145868
rect 249892 145852 249944 145858
rect 249892 145794 249944 145800
rect 270512 145761 270540 164183
rect 270498 145752 270554 145761
rect 270498 145687 270554 145696
rect 271892 145625 271920 165135
rect 273456 165034 273484 165543
rect 276032 165306 276060 165543
rect 276020 165300 276072 165306
rect 276020 165242 276072 165248
rect 278424 165238 278452 165543
rect 278412 165232 278464 165238
rect 275282 165200 275338 165209
rect 278412 165174 278464 165180
rect 280066 165200 280122 165209
rect 275282 165135 275338 165144
rect 280816 165170 280844 165543
rect 285968 165374 285996 165543
rect 293328 165510 293356 165543
rect 293316 165504 293368 165510
rect 293316 165446 293368 165452
rect 300872 165442 300900 165543
rect 311032 165543 311034 165552
rect 325882 165608 325938 165617
rect 325882 165543 325938 165552
rect 343270 165608 343326 165617
rect 343270 165543 343272 165552
rect 310980 165514 311032 165520
rect 300860 165436 300912 165442
rect 300860 165378 300912 165384
rect 285956 165368 286008 165374
rect 285956 165310 286008 165316
rect 280066 165135 280122 165144
rect 280804 165164 280856 165170
rect 273444 165028 273496 165034
rect 273444 164970 273496 164976
rect 273810 164384 273866 164393
rect 273810 164319 273866 164328
rect 273824 164286 273852 164319
rect 273812 164280 273864 164286
rect 273812 164222 273864 164228
rect 274546 164248 274602 164257
rect 274602 164206 274680 164234
rect 274546 164183 274602 164192
rect 274652 149054 274680 164206
rect 275296 149054 275324 165135
rect 276662 164248 276718 164257
rect 276662 164183 276718 164192
rect 277398 164248 277454 164257
rect 277398 164183 277454 164192
rect 274640 149048 274692 149054
rect 274640 148990 274692 148996
rect 274732 149048 274784 149054
rect 274732 148990 274784 148996
rect 275284 149048 275336 149054
rect 276676 149025 276704 164183
rect 275284 148990 275336 148996
rect 276018 149016 276074 149025
rect 274744 148374 274772 148990
rect 276018 148951 276074 148960
rect 276662 149016 276718 149025
rect 276662 148951 276718 148960
rect 274732 148368 274784 148374
rect 276032 148345 276060 148951
rect 274732 148310 274784 148316
rect 276018 148336 276074 148345
rect 276018 148271 276074 148280
rect 277412 146334 277440 164183
rect 277400 146328 277452 146334
rect 277400 146270 277452 146276
rect 280080 145654 280108 165135
rect 280804 165106 280856 165112
rect 325896 164121 325924 165543
rect 343324 165543 343326 165552
rect 343272 165514 343324 165520
rect 343546 164928 343602 164937
rect 343546 164863 343548 164872
rect 343600 164863 343602 164872
rect 343548 164834 343600 164840
rect 325882 164112 325938 164121
rect 325882 164047 325938 164056
rect 338488 146192 338540 146198
rect 338488 146134 338540 146140
rect 280068 145648 280120 145654
rect 271878 145616 271934 145625
rect 280068 145590 280120 145596
rect 271878 145551 271934 145560
rect 247132 145376 247184 145382
rect 247132 145318 247184 145324
rect 220084 145104 220136 145110
rect 220084 145046 220136 145052
rect 338500 144945 338528 146134
rect 340236 146124 340288 146130
rect 340236 146066 340288 146072
rect 340248 144945 340276 146066
rect 343560 145722 343588 164834
rect 356900 149054 356928 271118
rect 357084 165578 357112 271526
rect 357176 271318 357204 287026
rect 357164 271312 357216 271318
rect 357164 271254 357216 271260
rect 357072 165572 357124 165578
rect 357072 165514 357124 165520
rect 356888 149048 356940 149054
rect 357176 149025 357204 271254
rect 357360 253978 357388 358838
rect 357452 271386 357480 359518
rect 358096 359514 358124 389166
rect 358084 359508 358136 359514
rect 358084 359450 358136 359456
rect 358096 281518 358124 359450
rect 358084 281512 358136 281518
rect 358084 281454 358136 281460
rect 357440 271380 357492 271386
rect 357440 271322 357492 271328
rect 357348 253972 357400 253978
rect 357348 253914 357400 253920
rect 356888 148990 356940 148996
rect 357162 149016 357218 149025
rect 357162 148951 357218 148960
rect 357452 146266 357480 271322
rect 357532 254040 357584 254046
rect 357532 253982 357584 253988
rect 357544 253298 357572 253982
rect 357624 253972 357676 253978
rect 357624 253914 357676 253920
rect 357532 253292 357584 253298
rect 357532 253234 357584 253240
rect 357532 165572 357584 165578
rect 357532 165514 357584 165520
rect 357440 146260 357492 146266
rect 357440 146202 357492 146208
rect 343548 145716 343600 145722
rect 343548 145658 343600 145664
rect 356612 145716 356664 145722
rect 356612 145658 356664 145664
rect 351644 145580 351696 145586
rect 351644 145522 351696 145528
rect 351656 144945 351684 145522
rect 338486 144936 338542 144945
rect 338486 144871 338542 144880
rect 340234 144936 340290 144945
rect 340234 144871 340290 144880
rect 351642 144936 351698 144945
rect 351642 144871 351698 144880
rect 255870 59800 255926 59809
rect 255870 59735 255926 59744
rect 260654 59800 260710 59809
rect 260654 59735 260710 59744
rect 261758 59800 261814 59809
rect 261758 59735 261814 59744
rect 262862 59800 262918 59809
rect 262862 59735 262918 59744
rect 263874 59800 263930 59809
rect 263874 59735 263930 59744
rect 255884 59702 255912 59735
rect 255872 59696 255924 59702
rect 255872 59638 255924 59644
rect 256974 59664 257030 59673
rect 256974 59599 257030 59608
rect 256988 59226 257016 59599
rect 260668 59498 260696 59735
rect 261772 59566 261800 59735
rect 261760 59560 261812 59566
rect 261760 59502 261812 59508
rect 260656 59492 260708 59498
rect 260656 59434 260708 59440
rect 262876 59430 262904 59735
rect 263888 59634 263916 59735
rect 308494 59664 308550 59673
rect 263876 59628 263928 59634
rect 308494 59599 308550 59608
rect 263876 59570 263928 59576
rect 262864 59424 262916 59430
rect 259458 59392 259514 59401
rect 262864 59366 262916 59372
rect 259458 59327 259514 59336
rect 256976 59220 257028 59226
rect 256976 59162 257028 59168
rect 259472 59158 259500 59327
rect 295890 59256 295946 59265
rect 295890 59191 295946 59200
rect 298466 59256 298522 59265
rect 298466 59191 298522 59200
rect 303434 59256 303490 59265
rect 303434 59191 303490 59200
rect 259460 59152 259512 59158
rect 259460 59094 259512 59100
rect 295904 59022 295932 59191
rect 298480 59090 298508 59191
rect 298468 59084 298520 59090
rect 298468 59026 298520 59032
rect 295892 59016 295944 59022
rect 295892 58958 295944 58964
rect 303448 58886 303476 59191
rect 308508 58954 308536 59599
rect 308496 58948 308548 58954
rect 308496 58890 308548 58896
rect 303436 58880 303488 58886
rect 303436 58822 303488 58828
rect 222934 58576 222990 58585
rect 222934 58511 222990 58520
rect 222948 58313 222976 58511
rect 222934 58304 222990 58313
rect 222934 58239 222990 58248
rect 343180 57928 343232 57934
rect 236090 57896 236146 57905
rect 236090 57831 236146 57840
rect 238114 57896 238170 57905
rect 238114 57831 238170 57840
rect 238758 57896 238814 57905
rect 238758 57831 238814 57840
rect 240506 57896 240562 57905
rect 240506 57831 240562 57840
rect 241518 57896 241574 57905
rect 241518 57831 241574 57840
rect 242898 57896 242954 57905
rect 242898 57831 242954 57840
rect 244370 57896 244426 57905
rect 244370 57831 244426 57840
rect 245290 57896 245346 57905
rect 245290 57831 245346 57840
rect 245658 57896 245714 57905
rect 245658 57831 245714 57840
rect 247682 57896 247738 57905
rect 247682 57831 247738 57840
rect 248142 57896 248198 57905
rect 248142 57831 248198 57840
rect 248418 57896 248474 57905
rect 248418 57831 248474 57840
rect 249798 57896 249854 57905
rect 249798 57831 249854 57840
rect 251178 57896 251234 57905
rect 251178 57831 251234 57840
rect 251362 57896 251418 57905
rect 251362 57831 251418 57840
rect 253386 57896 253442 57905
rect 253386 57831 253442 57840
rect 253938 57896 253994 57905
rect 253938 57831 253994 57840
rect 271234 57896 271290 57905
rect 271234 57831 271290 57840
rect 271878 57896 271934 57905
rect 271878 57831 271934 57840
rect 273258 57896 273314 57905
rect 273258 57831 273314 57840
rect 275650 57896 275706 57905
rect 275650 57831 275706 57840
rect 278042 57896 278098 57905
rect 278042 57831 278098 57840
rect 279054 57896 279110 57905
rect 279054 57831 279110 57840
rect 287610 57896 287666 57905
rect 287610 57831 287666 57840
rect 293314 57896 293370 57905
rect 293314 57831 293370 57840
rect 300858 57896 300914 57905
rect 300858 57831 300914 57840
rect 305826 57896 305882 57905
rect 305826 57831 305882 57840
rect 310978 57896 311034 57905
rect 310978 57831 311034 57840
rect 313370 57896 313426 57905
rect 313370 57831 313426 57840
rect 315026 57896 315082 57905
rect 315026 57831 315082 57840
rect 318246 57896 318302 57905
rect 318246 57831 318302 57840
rect 325882 57896 325938 57905
rect 325882 57831 325884 57840
rect 235998 56944 236054 56953
rect 235998 56879 236054 56888
rect 219992 56296 220044 56302
rect 219992 56238 220044 56244
rect 236012 55146 236040 56879
rect 236000 55140 236052 55146
rect 236000 55082 236052 55088
rect 219716 55004 219768 55010
rect 219716 54946 219768 54952
rect 219164 54800 219216 54806
rect 219164 54742 219216 54748
rect 217232 54732 217284 54738
rect 217232 54674 217284 54680
rect 236104 54330 236132 57831
rect 238128 55894 238156 57831
rect 238116 55888 238168 55894
rect 238116 55830 238168 55836
rect 238772 54398 238800 57831
rect 240520 55826 240548 57831
rect 240508 55820 240560 55826
rect 240508 55762 240560 55768
rect 241532 54670 241560 57831
rect 241520 54664 241572 54670
rect 241520 54606 241572 54612
rect 242912 54602 242940 57831
rect 244384 55214 244412 57831
rect 245304 55962 245332 57831
rect 245292 55956 245344 55962
rect 245292 55898 245344 55904
rect 244372 55208 244424 55214
rect 244372 55150 244424 55156
rect 245672 54738 245700 57831
rect 247696 56030 247724 57831
rect 248156 57254 248184 57831
rect 248144 57248 248196 57254
rect 248144 57190 248196 57196
rect 247684 56024 247736 56030
rect 247684 55966 247736 55972
rect 248432 54874 248460 57831
rect 248420 54868 248472 54874
rect 248420 54810 248472 54816
rect 249812 54806 249840 57831
rect 251192 56166 251220 57831
rect 251180 56160 251232 56166
rect 251180 56102 251232 56108
rect 251376 54942 251404 57831
rect 253400 56098 253428 57831
rect 253388 56092 253440 56098
rect 253388 56034 253440 56040
rect 253952 55010 253980 57831
rect 263598 57760 263654 57769
rect 263598 57695 263654 57704
rect 265438 57760 265494 57769
rect 265438 57695 265494 57704
rect 266450 57760 266506 57769
rect 266450 57695 266506 57704
rect 268198 57760 268254 57769
rect 268198 57695 268254 57704
rect 268658 57760 268714 57769
rect 268658 57695 268714 57704
rect 269118 57760 269174 57769
rect 269118 57695 269174 57704
rect 263612 57322 263640 57695
rect 263600 57316 263652 57322
rect 263600 57258 263652 57264
rect 265452 56137 265480 57695
rect 266358 57352 266414 57361
rect 266358 57287 266414 57296
rect 266372 56234 266400 57287
rect 266360 56228 266412 56234
rect 266360 56170 266412 56176
rect 265438 56128 265494 56137
rect 265438 56063 265494 56072
rect 266464 55078 266492 57695
rect 268212 57458 268240 57695
rect 268200 57452 268252 57458
rect 268200 57394 268252 57400
rect 268672 56302 268700 57695
rect 268660 56296 268712 56302
rect 268660 56238 268712 56244
rect 266452 55072 266504 55078
rect 266452 55014 266504 55020
rect 253940 55004 253992 55010
rect 253940 54946 253992 54952
rect 251364 54936 251416 54942
rect 251364 54878 251416 54884
rect 249800 54800 249852 54806
rect 249800 54742 249852 54748
rect 245660 54732 245712 54738
rect 245660 54674 245712 54680
rect 242900 54596 242952 54602
rect 242900 54538 242952 54544
rect 269132 54466 269160 57695
rect 271248 56370 271276 57831
rect 271236 56364 271288 56370
rect 271236 56306 271288 56312
rect 271892 54534 271920 57831
rect 273272 56438 273300 57831
rect 273350 57760 273406 57769
rect 273350 57695 273406 57704
rect 273260 56432 273312 56438
rect 273260 56374 273312 56380
rect 273364 55185 273392 57695
rect 275664 56574 275692 57831
rect 276018 57760 276074 57769
rect 276018 57695 276074 57704
rect 275652 56568 275704 56574
rect 275652 56510 275704 56516
rect 273350 55176 273406 55185
rect 273350 55111 273406 55120
rect 276032 55049 276060 57695
rect 278056 56506 278084 57831
rect 279068 57458 279096 57831
rect 279056 57452 279108 57458
rect 279056 57394 279108 57400
rect 287624 57390 287652 57831
rect 293328 57526 293356 57831
rect 300872 57594 300900 57831
rect 305840 57662 305868 57831
rect 310992 57730 311020 57831
rect 313384 57798 313412 57831
rect 313372 57792 313424 57798
rect 313372 57734 313424 57740
rect 310980 57724 311032 57730
rect 310980 57666 311032 57672
rect 305828 57656 305880 57662
rect 305828 57598 305880 57604
rect 300860 57588 300912 57594
rect 300860 57530 300912 57536
rect 293316 57520 293368 57526
rect 293316 57462 293368 57468
rect 287612 57384 287664 57390
rect 287612 57326 287664 57332
rect 278044 56500 278096 56506
rect 278044 56442 278096 56448
rect 315040 56273 315068 57831
rect 318260 57186 318288 57831
rect 325936 57831 325938 57840
rect 343178 57896 343180 57905
rect 343232 57896 343234 57905
rect 343178 57831 343234 57840
rect 343454 57896 343510 57905
rect 356624 57866 356652 145658
rect 356704 145648 356756 145654
rect 356704 145590 356756 145596
rect 343454 57831 343456 57840
rect 325884 57802 325936 57808
rect 343508 57831 343510 57840
rect 356612 57860 356664 57866
rect 343456 57802 343508 57808
rect 356612 57802 356664 57808
rect 356716 57458 356744 145590
rect 357544 57934 357572 165514
rect 357636 146130 357664 253914
rect 357716 253292 357768 253298
rect 357716 253234 357768 253240
rect 357728 146198 357756 253234
rect 357716 146192 357768 146198
rect 357716 146134 357768 146140
rect 357624 146124 357676 146130
rect 357624 146066 357676 146072
rect 358084 68196 358136 68202
rect 358084 68138 358136 68144
rect 358096 59362 358124 68138
rect 358084 59356 358136 59362
rect 358084 59298 358136 59304
rect 358188 58954 358216 490690
rect 358280 166938 358308 490894
rect 360936 490680 360988 490686
rect 360936 490622 360988 490628
rect 359740 489388 359792 489394
rect 359740 489330 359792 489336
rect 358728 484220 358780 484226
rect 358728 484162 358780 484168
rect 358452 478372 358504 478378
rect 358452 478314 358504 478320
rect 358360 465996 358412 466002
rect 358360 465938 358412 465944
rect 358268 166932 358320 166938
rect 358268 166874 358320 166880
rect 358372 165442 358400 465938
rect 358464 273290 358492 478314
rect 358544 475652 358596 475658
rect 358544 475594 358596 475600
rect 358452 273284 358504 273290
rect 358452 273226 358504 273232
rect 358556 273193 358584 475594
rect 358636 469056 358688 469062
rect 358636 468998 358688 469004
rect 358648 284306 358676 468998
rect 358740 380934 358768 484162
rect 359648 470416 359700 470422
rect 359648 470358 359700 470364
rect 359464 469192 359516 469198
rect 359464 469134 359516 469140
rect 358820 466472 358872 466478
rect 358820 466414 358872 466420
rect 358832 390522 358860 466414
rect 358912 465112 358964 465118
rect 358912 465054 358964 465060
rect 358924 460934 358952 465054
rect 358924 460906 359412 460934
rect 359384 460193 359412 460906
rect 359370 460184 359426 460193
rect 359370 460119 359426 460128
rect 359094 400344 359150 400353
rect 359094 400279 359150 400288
rect 359002 398168 359058 398177
rect 359002 398103 359058 398112
rect 358820 390516 358872 390522
rect 358820 390458 358872 390464
rect 358832 389230 358860 390458
rect 358820 389224 358872 389230
rect 358820 389166 358872 389172
rect 358728 380928 358780 380934
rect 358728 380870 358780 380876
rect 358820 378616 358872 378622
rect 358820 378558 358872 378564
rect 358636 284300 358688 284306
rect 358636 284242 358688 284248
rect 358542 273184 358598 273193
rect 358542 273119 358598 273128
rect 358832 271454 358860 378558
rect 359016 374746 359044 398103
rect 359004 374740 359056 374746
rect 359004 374682 359056 374688
rect 359108 371210 359136 400279
rect 359280 378616 359332 378622
rect 359280 378558 359332 378564
rect 359292 378282 359320 378558
rect 359280 378276 359332 378282
rect 359280 378218 359332 378224
rect 359096 371204 359148 371210
rect 359096 371146 359148 371152
rect 359108 369238 359136 371146
rect 359096 369232 359148 369238
rect 359096 369174 359148 369180
rect 358912 369164 358964 369170
rect 358912 369106 358964 369112
rect 358924 291009 358952 369106
rect 359188 363520 359240 363526
rect 359188 363462 359240 363468
rect 359096 358964 359148 358970
rect 359096 358906 359148 358912
rect 358910 291000 358966 291009
rect 358910 290935 358966 290944
rect 358820 271448 358872 271454
rect 358820 271390 358872 271396
rect 358820 271312 358872 271318
rect 358820 271254 358872 271260
rect 358728 176180 358780 176186
rect 358728 176122 358780 176128
rect 358360 165436 358412 165442
rect 358360 165378 358412 165384
rect 358740 146266 358768 176122
rect 358728 146260 358780 146266
rect 358728 146202 358780 146208
rect 358740 145586 358768 146202
rect 358832 145654 358860 271254
rect 358924 183569 358952 290935
rect 359108 271930 359136 358906
rect 359200 288833 359228 363462
rect 359280 361616 359332 361622
rect 359280 361558 359332 361564
rect 359186 288824 359242 288833
rect 359186 288759 359242 288768
rect 359096 271924 359148 271930
rect 359096 271866 359148 271872
rect 359002 245712 359058 245721
rect 359002 245647 359058 245656
rect 358910 183560 358966 183569
rect 358910 183495 358966 183504
rect 358820 145648 358872 145654
rect 358820 145590 358872 145596
rect 358728 145580 358780 145586
rect 358728 145522 358780 145528
rect 358740 68338 358768 145522
rect 359016 139369 359044 245647
rect 359200 181937 359228 288759
rect 359292 288425 359320 361558
rect 359384 354674 359412 460119
rect 359476 376174 359504 469134
rect 359556 468988 359608 468994
rect 359556 468930 359608 468936
rect 359568 389162 359596 468930
rect 359660 391950 359688 470358
rect 359752 411942 359780 489330
rect 359832 485240 359884 485246
rect 359832 485182 359884 485188
rect 359844 413302 359872 485182
rect 360844 481296 360896 481302
rect 360844 481238 360896 481244
rect 360752 478780 360804 478786
rect 360752 478722 360804 478728
rect 360660 478576 360712 478582
rect 360660 478518 360712 478524
rect 360016 470552 360068 470558
rect 360016 470494 360068 470500
rect 359924 470484 359976 470490
rect 359924 470426 359976 470432
rect 359832 413296 359884 413302
rect 359832 413238 359884 413244
rect 359740 411936 359792 411942
rect 359740 411878 359792 411884
rect 359936 409154 359964 470426
rect 360028 410582 360056 470494
rect 360568 467832 360620 467838
rect 360568 467774 360620 467780
rect 360016 410576 360068 410582
rect 360016 410518 360068 410524
rect 359924 409148 359976 409154
rect 359924 409090 359976 409096
rect 359738 396808 359794 396817
rect 359738 396743 359794 396752
rect 359648 391944 359700 391950
rect 359648 391886 359700 391892
rect 359556 389156 359608 389162
rect 359556 389098 359608 389104
rect 359464 376168 359516 376174
rect 359464 376110 359516 376116
rect 359648 374740 359700 374746
rect 359648 374682 359700 374688
rect 359464 372632 359516 372638
rect 359464 372574 359516 372580
rect 359476 362234 359504 372574
rect 359556 369232 359608 369238
rect 359556 369174 359608 369180
rect 359464 362228 359516 362234
rect 359464 362170 359516 362176
rect 359476 361622 359504 362170
rect 359464 361616 359516 361622
rect 359464 361558 359516 361564
rect 359384 354646 359504 354674
rect 359476 353161 359504 354646
rect 359462 353152 359518 353161
rect 359462 353087 359518 353096
rect 359370 292768 359426 292777
rect 359370 292703 359426 292712
rect 359278 288416 359334 288425
rect 359278 288351 359334 288360
rect 359384 190454 359412 292703
rect 359476 245721 359504 353087
rect 359568 292777 359596 369174
rect 359660 365022 359688 374682
rect 359752 370530 359780 396743
rect 359922 395312 359978 395321
rect 359922 395247 359978 395256
rect 359830 394088 359886 394097
rect 359830 394023 359886 394032
rect 359844 373318 359872 394023
rect 359936 376038 359964 395247
rect 360580 380594 360608 467774
rect 360568 380588 360620 380594
rect 360568 380530 360620 380536
rect 360672 380254 360700 478518
rect 360660 380248 360712 380254
rect 360660 380190 360712 380196
rect 360764 378894 360792 478722
rect 360752 378888 360804 378894
rect 360752 378830 360804 378836
rect 360016 378548 360068 378554
rect 360016 378490 360068 378496
rect 359924 376032 359976 376038
rect 359924 375974 359976 375980
rect 359832 373312 359884 373318
rect 359832 373254 359884 373260
rect 359844 372638 359872 373254
rect 359832 372632 359884 372638
rect 359832 372574 359884 372580
rect 359740 370524 359792 370530
rect 359740 370466 359792 370472
rect 359752 369170 359780 370466
rect 359740 369164 359792 369170
rect 359740 369106 359792 369112
rect 359648 365016 359700 365022
rect 359648 364958 359700 364964
rect 359554 292768 359610 292777
rect 359554 292703 359610 292712
rect 359660 291825 359688 364958
rect 359936 363526 359964 375974
rect 359924 363520 359976 363526
rect 359924 363462 359976 363468
rect 359646 291816 359702 291825
rect 359646 291751 359702 291760
rect 359554 288416 359610 288425
rect 359554 288351 359610 288360
rect 359568 287609 359596 288351
rect 359554 287600 359610 287609
rect 359554 287535 359610 287544
rect 359462 245712 359518 245721
rect 359462 245647 359518 245656
rect 359384 190426 359504 190454
rect 359476 186425 359504 190426
rect 359462 186416 359518 186425
rect 359462 186351 359518 186360
rect 359278 184920 359334 184929
rect 359278 184855 359334 184864
rect 359186 181928 359242 181937
rect 359186 181863 359242 181872
rect 359094 179480 359150 179489
rect 359094 179415 359150 179424
rect 359002 139360 359058 139369
rect 359002 139295 359058 139304
rect 359108 74089 359136 179415
rect 359200 75449 359228 181863
rect 359292 78305 359320 184855
rect 359370 183560 359426 183569
rect 359370 183495 359426 183504
rect 359278 78296 359334 78305
rect 359278 78231 359334 78240
rect 359384 76945 359412 183495
rect 359476 79937 359504 186351
rect 359568 180713 359596 287535
rect 359660 184929 359688 291751
rect 360028 271318 360056 378490
rect 360856 378146 360884 481238
rect 360844 378140 360896 378146
rect 360844 378082 360896 378088
rect 360292 359304 360344 359310
rect 360292 359246 360344 359252
rect 360304 358834 360332 359246
rect 360292 358828 360344 358834
rect 360292 358770 360344 358776
rect 360200 281512 360252 281518
rect 360200 281454 360252 281460
rect 360016 271312 360068 271318
rect 360016 271254 360068 271260
rect 360212 253230 360240 281454
rect 360304 254046 360332 358770
rect 360292 254040 360344 254046
rect 360292 253982 360344 253988
rect 360200 253224 360252 253230
rect 360200 253166 360252 253172
rect 359646 184920 359702 184929
rect 359646 184855 359702 184864
rect 359554 180704 359610 180713
rect 359554 180639 359610 180648
rect 359568 179489 359596 180639
rect 359554 179480 359610 179489
rect 359554 179415 359610 179424
rect 360212 176662 360240 253166
rect 360292 251864 360344 251870
rect 360292 251806 360344 251812
rect 360200 176656 360252 176662
rect 360200 176598 360252 176604
rect 360212 176186 360240 176598
rect 360200 176180 360252 176186
rect 360200 176122 360252 176128
rect 360304 164898 360332 251806
rect 360292 164892 360344 164898
rect 360292 164834 360344 164840
rect 359462 79928 359518 79937
rect 359462 79863 359518 79872
rect 359370 76936 359426 76945
rect 359370 76871 359426 76880
rect 359186 75440 359242 75449
rect 359186 75375 359242 75384
rect 359094 74080 359150 74089
rect 359094 74015 359150 74024
rect 358728 68332 358780 68338
rect 358728 68274 358780 68280
rect 358740 68202 358768 68274
rect 358728 68196 358780 68202
rect 358728 68138 358780 68144
rect 360948 59430 360976 490622
rect 361028 489252 361080 489258
rect 361028 489194 361080 489200
rect 361040 165102 361068 489194
rect 361132 166462 361160 491098
rect 362684 478848 362736 478854
rect 362684 478790 362736 478796
rect 362500 478304 362552 478310
rect 362500 478246 362552 478252
rect 361396 475856 361448 475862
rect 361396 475798 361448 475804
rect 361212 475516 361264 475522
rect 361212 475458 361264 475464
rect 361224 273494 361252 475458
rect 361304 467492 361356 467498
rect 361304 467434 361356 467440
rect 361316 282878 361344 467434
rect 361408 374814 361436 475798
rect 362316 475380 362368 475386
rect 362316 475322 362368 475328
rect 362224 472796 362276 472802
rect 362224 472738 362276 472744
rect 361580 466608 361632 466614
rect 361580 466550 361632 466556
rect 361486 379536 361542 379545
rect 361486 379471 361542 379480
rect 361396 374808 361448 374814
rect 361396 374750 361448 374756
rect 361304 282872 361356 282878
rect 361304 282814 361356 282820
rect 361212 273488 361264 273494
rect 361212 273430 361264 273436
rect 361120 166456 361172 166462
rect 361120 166398 361172 166404
rect 361028 165096 361080 165102
rect 361028 165038 361080 165044
rect 360936 59424 360988 59430
rect 360936 59366 360988 59372
rect 358176 58948 358228 58954
rect 358176 58890 358228 58896
rect 361500 57934 361528 379471
rect 361592 359310 361620 466550
rect 362132 465656 362184 465662
rect 362132 465598 362184 465604
rect 362144 380186 362172 465598
rect 362132 380180 362184 380186
rect 362132 380122 362184 380128
rect 361580 359304 361632 359310
rect 361580 359246 361632 359252
rect 357532 57928 357584 57934
rect 357532 57870 357584 57876
rect 361488 57928 361540 57934
rect 361488 57870 361540 57876
rect 362236 57526 362264 472738
rect 362328 165578 362356 475322
rect 362408 474088 362460 474094
rect 362408 474030 362460 474036
rect 362420 175234 362448 474030
rect 362512 271726 362540 478246
rect 362592 473272 362644 473278
rect 362592 473214 362644 473220
rect 362604 272542 362632 473214
rect 362696 374882 362724 478790
rect 362776 478644 362828 478650
rect 362776 478586 362828 478592
rect 362788 376446 362816 478586
rect 363512 468376 363564 468382
rect 363512 468318 363564 468324
rect 362960 466540 363012 466546
rect 362960 466482 363012 466488
rect 362868 465588 362920 465594
rect 362868 465530 362920 465536
rect 362776 376440 362828 376446
rect 362776 376382 362828 376388
rect 362684 374876 362736 374882
rect 362684 374818 362736 374824
rect 362880 374678 362908 465530
rect 362868 374672 362920 374678
rect 362868 374614 362920 374620
rect 362972 358902 363000 466482
rect 363524 377466 363552 468318
rect 363512 377460 363564 377466
rect 363512 377402 363564 377408
rect 362960 358896 363012 358902
rect 362960 358838 363012 358844
rect 362592 272536 362644 272542
rect 362592 272478 362644 272484
rect 362500 271720 362552 271726
rect 362500 271662 362552 271668
rect 362408 175228 362460 175234
rect 362408 175170 362460 175176
rect 362316 165572 362368 165578
rect 362316 165514 362368 165520
rect 362224 57520 362276 57526
rect 362224 57462 362276 57468
rect 356704 57452 356756 57458
rect 356704 57394 356756 57400
rect 318248 57180 318300 57186
rect 318248 57122 318300 57128
rect 315026 56264 315082 56273
rect 315026 56199 315082 56208
rect 276018 55040 276074 55049
rect 276018 54975 276074 54984
rect 271880 54528 271932 54534
rect 271880 54470 271932 54476
rect 269120 54460 269172 54466
rect 269120 54402 269172 54408
rect 238760 54392 238812 54398
rect 238760 54334 238812 54340
rect 216496 54324 216548 54330
rect 216496 54266 216548 54272
rect 236092 54324 236144 54330
rect 236092 54266 236144 54272
rect 143538 4040 143594 4049
rect 143538 3975 143594 3984
rect 136454 3904 136510 3913
rect 136454 3839 136510 3848
rect 132958 3496 133014 3505
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 57244 3460 57296 3466
rect 57244 3402 57296 3408
rect 125876 3460 125928 3466
rect 132958 3431 133014 3440
rect 125876 3402 125928 3408
rect 584 480 612 3402
rect 125888 480 125916 3402
rect 129370 3360 129426 3369
rect 129370 3295 129426 3304
rect 129384 480 129412 3295
rect 132972 480 133000 3431
rect 136468 480 136496 3839
rect 140042 3768 140098 3777
rect 140042 3703 140098 3712
rect 140056 480 140084 3703
rect 143552 480 143580 3975
rect 150622 3632 150678 3641
rect 150622 3567 150678 3576
rect 147128 3528 147180 3534
rect 147128 3470 147180 3476
rect 147140 480 147168 3470
rect 150636 480 150664 3567
rect 363616 3534 363644 527818
rect 383672 491978 383700 534126
rect 388456 532234 388484 534126
rect 393332 532506 393360 534126
rect 397472 534126 397808 534154
rect 401980 534126 402316 534154
rect 406488 534126 406824 534154
rect 411332 534126 411392 534154
rect 393320 532500 393372 532506
rect 393320 532442 393372 532448
rect 388444 532228 388496 532234
rect 388444 532170 388496 532176
rect 397472 529145 397500 534126
rect 401980 532370 402008 534126
rect 406488 532438 406516 534126
rect 406476 532432 406528 532438
rect 406476 532374 406528 532380
rect 401968 532364 402020 532370
rect 401968 532306 402020 532312
rect 411364 531894 411392 534126
rect 415504 534126 415840 534154
rect 420012 534126 420348 534154
rect 424520 534126 424856 534154
rect 429212 534126 429364 534154
rect 411352 531888 411404 531894
rect 411352 531830 411404 531836
rect 415504 531826 415532 534126
rect 420012 532778 420040 534126
rect 420000 532772 420052 532778
rect 420000 532714 420052 532720
rect 424520 532642 424548 534126
rect 429212 532681 429240 534126
rect 433352 533798 433380 611351
rect 433430 601760 433486 601769
rect 433430 601695 433486 601704
rect 433444 535106 433472 601695
rect 433522 586800 433578 586809
rect 433522 586735 433578 586744
rect 433536 535378 433564 586735
rect 433614 572656 433670 572665
rect 433614 572591 433670 572600
rect 433628 538214 433656 572591
rect 434626 538928 434682 538937
rect 434626 538863 434682 538872
rect 433628 538186 433840 538214
rect 433536 535350 433748 535378
rect 433444 535078 433564 535106
rect 433430 534984 433486 534993
rect 433430 534919 433486 534928
rect 433340 533792 433392 533798
rect 433340 533734 433392 533740
rect 429198 532672 429254 532681
rect 424508 532636 424560 532642
rect 429198 532607 429254 532616
rect 424508 532578 424560 532584
rect 415492 531820 415544 531826
rect 415492 531762 415544 531768
rect 433444 529514 433472 534919
rect 433536 529650 433564 535078
rect 433524 529644 433576 529650
rect 433524 529586 433576 529592
rect 433720 529582 433748 535350
rect 433812 533458 433840 538186
rect 434640 533730 434668 538863
rect 434628 533724 434680 533730
rect 434628 533666 434680 533672
rect 433800 533452 433852 533458
rect 433800 533394 433852 533400
rect 433708 529576 433760 529582
rect 433708 529518 433760 529524
rect 433432 529508 433484 529514
rect 433432 529450 433484 529456
rect 434732 529446 434760 700334
rect 434812 700324 434864 700330
rect 434812 700266 434864 700272
rect 434824 640257 434852 700266
rect 434904 653404 434956 653410
rect 434904 653346 434956 653352
rect 434810 640248 434866 640257
rect 434810 640183 434866 640192
rect 434810 596728 434866 596737
rect 434810 596663 434866 596672
rect 434720 529440 434772 529446
rect 434720 529382 434772 529388
rect 397458 529136 397514 529145
rect 397458 529071 397514 529080
rect 383660 491972 383712 491978
rect 383660 491914 383712 491920
rect 365168 490884 365220 490890
rect 365168 490826 365220 490832
rect 363696 490816 363748 490822
rect 363696 490758 363748 490764
rect 363708 58886 363736 490758
rect 363788 487892 363840 487898
rect 363788 487834 363840 487840
rect 363800 164801 363828 487834
rect 363880 486532 363932 486538
rect 363880 486474 363932 486480
rect 363892 164966 363920 486474
rect 364156 481228 364208 481234
rect 364156 481170 364208 481176
rect 363972 473204 364024 473210
rect 363972 473146 364024 473152
rect 363984 272610 364012 473146
rect 364064 467628 364116 467634
rect 364064 467570 364116 467576
rect 363972 272604 364024 272610
rect 363972 272546 364024 272552
rect 364076 270881 364104 467570
rect 364168 376650 364196 481170
rect 364892 481092 364944 481098
rect 364892 481034 364944 481040
rect 364248 478508 364300 478514
rect 364248 478450 364300 478456
rect 364260 380390 364288 478450
rect 364800 475720 364852 475726
rect 364800 475662 364852 475668
rect 364248 380384 364300 380390
rect 364248 380326 364300 380332
rect 364156 376644 364208 376650
rect 364156 376586 364208 376592
rect 364812 376378 364840 475662
rect 364904 380322 364932 481034
rect 364984 476808 365036 476814
rect 364984 476750 365036 476756
rect 364892 380316 364944 380322
rect 364892 380258 364944 380264
rect 364800 376372 364852 376378
rect 364800 376314 364852 376320
rect 364062 270872 364118 270881
rect 364062 270807 364118 270816
rect 363880 164960 363932 164966
rect 363880 164902 363932 164908
rect 363786 164792 363842 164801
rect 363786 164727 363842 164736
rect 363696 58880 363748 58886
rect 363696 58822 363748 58828
rect 364996 57730 365024 476750
rect 365076 472728 365128 472734
rect 365076 472670 365128 472676
rect 364984 57724 365036 57730
rect 364984 57666 365036 57672
rect 365088 57254 365116 472670
rect 365180 166190 365208 490826
rect 374644 490612 374696 490618
rect 374644 490554 374696 490560
rect 373540 489320 373592 489326
rect 373540 489262 373592 489268
rect 367928 487960 367980 487966
rect 367928 487902 367980 487908
rect 366732 486600 366784 486606
rect 366732 486542 366784 486548
rect 366548 483812 366600 483818
rect 366548 483754 366600 483760
rect 366456 483744 366508 483750
rect 366456 483686 366508 483692
rect 365628 481432 365680 481438
rect 365628 481374 365680 481380
rect 365444 480956 365496 480962
rect 365444 480898 365496 480904
rect 365260 470008 365312 470014
rect 365260 469950 365312 469956
rect 365272 166326 365300 469950
rect 365352 467424 365404 467430
rect 365352 467366 365404 467372
rect 365364 178022 365392 467366
rect 365456 271522 365484 480898
rect 365536 473136 365588 473142
rect 365536 473078 365588 473084
rect 365548 273057 365576 473078
rect 365640 375018 365668 481374
rect 366272 475584 366324 475590
rect 366272 475526 366324 475532
rect 366180 471776 366232 471782
rect 366180 471718 366232 471724
rect 366192 377398 366220 471718
rect 366284 380458 366312 475526
rect 366362 472696 366418 472705
rect 366362 472631 366418 472640
rect 366272 380452 366324 380458
rect 366272 380394 366324 380400
rect 366180 377392 366232 377398
rect 366180 377334 366232 377340
rect 365628 375012 365680 375018
rect 365628 374954 365680 374960
rect 365534 273048 365590 273057
rect 365534 272983 365590 272992
rect 365444 271516 365496 271522
rect 365444 271458 365496 271464
rect 365352 178016 365404 178022
rect 365352 177958 365404 177964
rect 365260 166320 365312 166326
rect 365260 166262 365312 166268
rect 365168 166184 365220 166190
rect 365168 166126 365220 166132
rect 365076 57248 365128 57254
rect 365076 57190 365128 57196
rect 363604 3528 363656 3534
rect 363604 3470 363656 3476
rect 366376 3466 366404 472631
rect 366468 57662 366496 483686
rect 366560 165170 366588 483754
rect 366640 469872 366692 469878
rect 366640 469814 366692 469820
rect 366652 167006 366680 469814
rect 366744 271794 366772 486542
rect 367008 481160 367060 481166
rect 367008 481102 367060 481108
rect 366824 468580 366876 468586
rect 366824 468522 366876 468528
rect 366836 273018 366864 468522
rect 366916 466132 366968 466138
rect 366916 466074 366968 466080
rect 366824 273012 366876 273018
rect 366824 272954 366876 272960
rect 366732 271788 366784 271794
rect 366732 271730 366784 271736
rect 366928 271318 366956 466074
rect 367020 376582 367048 481102
rect 367652 481024 367704 481030
rect 367652 480966 367704 480972
rect 367560 469124 367612 469130
rect 367560 469066 367612 469072
rect 367468 464432 367520 464438
rect 367468 464374 367520 464380
rect 367008 376576 367060 376582
rect 367008 376518 367060 376524
rect 367480 375222 367508 464374
rect 367572 377874 367600 469066
rect 367560 377868 367612 377874
rect 367560 377810 367612 377816
rect 367664 377670 367692 480966
rect 367744 479596 367796 479602
rect 367744 479538 367796 479544
rect 367652 377664 367704 377670
rect 367652 377606 367704 377612
rect 367468 375216 367520 375222
rect 367468 375158 367520 375164
rect 367008 374740 367060 374746
rect 367008 374682 367060 374688
rect 367020 271658 367048 374682
rect 367008 271652 367060 271658
rect 367008 271594 367060 271600
rect 366916 271312 366968 271318
rect 366916 271254 366968 271260
rect 366640 167000 366692 167006
rect 366640 166942 366692 166948
rect 366548 165164 366600 165170
rect 366548 165106 366600 165112
rect 366456 57656 366508 57662
rect 366456 57598 366508 57604
rect 367756 57458 367784 479538
rect 367836 467356 367888 467362
rect 367836 467298 367888 467304
rect 367848 166666 367876 467298
rect 367940 271250 367968 487902
rect 370504 487824 370556 487830
rect 370504 487766 370556 487772
rect 368020 485172 368072 485178
rect 368020 485114 368072 485120
rect 368032 271862 368060 485114
rect 369124 485104 369176 485110
rect 369124 485046 369176 485052
rect 368204 484356 368256 484362
rect 368204 484298 368256 484304
rect 368112 466064 368164 466070
rect 368112 466006 368164 466012
rect 368124 273358 368152 466006
rect 368216 375086 368244 484298
rect 368388 481364 368440 481370
rect 368388 481306 368440 481312
rect 368400 378962 368428 481306
rect 369032 474224 369084 474230
rect 369032 474166 369084 474172
rect 368848 468784 368900 468790
rect 368848 468726 368900 468732
rect 368860 380526 368888 468726
rect 368940 466404 368992 466410
rect 368940 466346 368992 466352
rect 368848 380520 368900 380526
rect 368848 380462 368900 380468
rect 368388 378956 368440 378962
rect 368388 378898 368440 378904
rect 368296 378548 368348 378554
rect 368296 378490 368348 378496
rect 368204 375080 368256 375086
rect 368204 375022 368256 375028
rect 368112 273352 368164 273358
rect 368112 273294 368164 273300
rect 368020 271856 368072 271862
rect 368020 271798 368072 271804
rect 367928 271244 367980 271250
rect 367928 271186 367980 271192
rect 368308 270366 368336 378490
rect 368952 378078 368980 466346
rect 369044 378418 369072 474166
rect 369032 378412 369084 378418
rect 369032 378354 369084 378360
rect 368940 378072 368992 378078
rect 368940 378014 368992 378020
rect 368388 376780 368440 376786
rect 368388 376722 368440 376728
rect 368296 270360 368348 270366
rect 368296 270302 368348 270308
rect 367836 166660 367888 166666
rect 367836 166602 367888 166608
rect 368308 147558 368336 270302
rect 368400 251938 368428 376722
rect 369032 273556 369084 273562
rect 369032 273498 369084 273504
rect 368388 251932 368440 251938
rect 368388 251874 368440 251880
rect 368296 147552 368348 147558
rect 368296 147494 368348 147500
rect 369044 145625 369072 273498
rect 369136 164898 369164 485046
rect 369400 483880 369452 483886
rect 369400 483822 369452 483828
rect 369216 478236 369268 478242
rect 369216 478178 369268 478184
rect 369228 165510 369256 478178
rect 369308 467288 369360 467294
rect 369308 467230 369360 467236
rect 369320 166598 369348 467230
rect 369412 271590 369440 483822
rect 370412 471640 370464 471646
rect 370412 471582 370464 471588
rect 369768 471572 369820 471578
rect 369768 471514 369820 471520
rect 369492 466268 369544 466274
rect 369492 466210 369544 466216
rect 369504 272882 369532 466210
rect 369584 380588 369636 380594
rect 369584 380530 369636 380536
rect 369596 379642 369624 380530
rect 369780 379710 369808 471514
rect 370320 468852 370372 468858
rect 370320 468794 370372 468800
rect 370228 464500 370280 464506
rect 370228 464442 370280 464448
rect 369768 379704 369820 379710
rect 369768 379646 369820 379652
rect 369584 379636 369636 379642
rect 369584 379578 369636 379584
rect 369676 379568 369728 379574
rect 369676 379510 369728 379516
rect 369584 378684 369636 378690
rect 369584 378626 369636 378632
rect 369596 378350 369624 378626
rect 369584 378344 369636 378350
rect 369584 378286 369636 378292
rect 369596 376961 369624 378286
rect 369582 376952 369638 376961
rect 369582 376887 369638 376896
rect 369584 376848 369636 376854
rect 369584 376790 369636 376796
rect 369492 272876 369544 272882
rect 369492 272818 369544 272824
rect 369400 271584 369452 271590
rect 369400 271526 369452 271532
rect 369596 270473 369624 376790
rect 369582 270464 369638 270473
rect 369582 270399 369638 270408
rect 369688 251870 369716 379510
rect 369768 379500 369820 379506
rect 369768 379442 369820 379448
rect 369780 377058 369808 379442
rect 369858 379128 369914 379137
rect 369858 379063 369914 379072
rect 369872 378729 369900 379063
rect 369858 378720 369914 378729
rect 369858 378655 369914 378664
rect 369768 377052 369820 377058
rect 369768 376994 369820 377000
rect 369766 376952 369822 376961
rect 369766 376887 369822 376896
rect 369780 270502 369808 376887
rect 370240 375154 370268 464442
rect 370332 377738 370360 468794
rect 370424 378622 370452 471582
rect 370412 378616 370464 378622
rect 370412 378558 370464 378564
rect 370320 377732 370372 377738
rect 370320 377674 370372 377680
rect 370228 375148 370280 375154
rect 370228 375090 370280 375096
rect 370412 271924 370464 271930
rect 370412 271866 370464 271872
rect 370424 271658 370452 271866
rect 370412 271652 370464 271658
rect 370412 271594 370464 271600
rect 369768 270496 369820 270502
rect 369768 270438 369820 270444
rect 369676 251864 369728 251870
rect 369676 251806 369728 251812
rect 369308 166592 369360 166598
rect 369308 166534 369360 166540
rect 370424 166122 370452 271594
rect 370412 166116 370464 166122
rect 370412 166058 370464 166064
rect 369216 165504 369268 165510
rect 369216 165446 369268 165452
rect 369124 164892 369176 164898
rect 369124 164834 369176 164840
rect 369030 145616 369086 145625
rect 369030 145551 369086 145560
rect 370516 70378 370544 487766
rect 370964 484016 371016 484022
rect 370964 483958 371016 483964
rect 370596 482384 370648 482390
rect 370596 482326 370648 482332
rect 370608 165374 370636 482326
rect 370872 476944 370924 476950
rect 370872 476886 370924 476892
rect 370688 472864 370740 472870
rect 370688 472806 370740 472812
rect 370596 165368 370648 165374
rect 370596 165310 370648 165316
rect 370700 164150 370728 472806
rect 370780 467152 370832 467158
rect 370780 467094 370832 467100
rect 370792 166734 370820 467094
rect 370884 271454 370912 476886
rect 370976 375970 371004 483958
rect 371884 476876 371936 476882
rect 371884 476818 371936 476824
rect 371792 471368 371844 471374
rect 371792 471310 371844 471316
rect 371240 467764 371292 467770
rect 371240 467706 371292 467712
rect 371148 379704 371200 379710
rect 371148 379646 371200 379652
rect 371054 379128 371110 379137
rect 371054 379063 371110 379072
rect 370964 375964 371016 375970
rect 370964 375906 371016 375912
rect 370964 374672 371016 374678
rect 370964 374614 371016 374620
rect 370872 271448 370924 271454
rect 370872 271390 370924 271396
rect 370976 269074 371004 374614
rect 371068 270026 371096 379063
rect 371160 270094 371188 379646
rect 371252 379574 371280 467706
rect 371240 379568 371292 379574
rect 371240 379510 371292 379516
rect 371606 379536 371662 379545
rect 371606 379471 371662 379480
rect 371148 270088 371200 270094
rect 371148 270030 371200 270036
rect 371056 270020 371108 270026
rect 371056 269962 371108 269968
rect 371620 269929 371648 379471
rect 371804 376242 371832 471310
rect 371792 376236 371844 376242
rect 371792 376178 371844 376184
rect 371790 273320 371846 273329
rect 371790 273255 371846 273264
rect 371700 270496 371752 270502
rect 371700 270438 371752 270444
rect 371712 270162 371740 270438
rect 371700 270156 371752 270162
rect 371700 270098 371752 270104
rect 371606 269920 371662 269929
rect 371606 269855 371662 269864
rect 370964 269068 371016 269074
rect 370964 269010 371016 269016
rect 371148 251932 371200 251938
rect 371148 251874 371200 251880
rect 371056 251864 371108 251870
rect 371056 251806 371108 251812
rect 370780 166728 370832 166734
rect 370780 166670 370832 166676
rect 370688 164144 370740 164150
rect 370688 164086 370740 164092
rect 371068 163441 371096 251806
rect 371160 163538 371188 251874
rect 371148 163532 371200 163538
rect 371148 163474 371200 163480
rect 371054 163432 371110 163441
rect 371054 163367 371110 163376
rect 371712 145518 371740 270098
rect 371804 146305 371832 273255
rect 371896 165238 371924 476818
rect 372068 474156 372120 474162
rect 372068 474098 372120 474104
rect 371976 467220 372028 467226
rect 371976 467162 372028 467168
rect 371988 166530 372016 467162
rect 372080 271386 372108 474098
rect 373080 471912 373132 471918
rect 373080 471854 373132 471860
rect 372436 471844 372488 471850
rect 372436 471786 372488 471792
rect 372252 468716 372304 468722
rect 372252 468658 372304 468664
rect 372160 466200 372212 466206
rect 372160 466142 372212 466148
rect 372172 272814 372200 466142
rect 372264 380594 372292 468658
rect 372252 380588 372304 380594
rect 372252 380530 372304 380536
rect 372342 378856 372398 378865
rect 372342 378791 372398 378800
rect 372252 377392 372304 377398
rect 372252 377334 372304 377340
rect 372160 272808 372212 272814
rect 372160 272750 372212 272756
rect 372068 271380 372120 271386
rect 372068 271322 372120 271328
rect 372158 270464 372214 270473
rect 372158 270399 372214 270408
rect 372068 270020 372120 270026
rect 372068 269962 372120 269968
rect 371976 166524 372028 166530
rect 371976 166466 372028 166472
rect 371884 165232 371936 165238
rect 371884 165174 371936 165180
rect 372080 148442 372108 269962
rect 372172 269793 372200 270399
rect 372158 269784 372214 269793
rect 372158 269719 372214 269728
rect 372172 163198 372200 269719
rect 372264 268530 372292 377334
rect 372356 269754 372384 378791
rect 372448 375290 372476 471786
rect 372988 466336 373040 466342
rect 372988 466278 373040 466284
rect 373000 377806 373028 466278
rect 372988 377800 373040 377806
rect 373092 377777 373120 471854
rect 373172 471300 373224 471306
rect 373172 471242 373224 471248
rect 372988 377742 373040 377748
rect 373078 377768 373134 377777
rect 373078 377703 373134 377712
rect 373184 377602 373212 471242
rect 373356 469940 373408 469946
rect 373356 469882 373408 469888
rect 373262 465760 373318 465769
rect 373262 465695 373318 465704
rect 373172 377596 373224 377602
rect 373172 377538 373224 377544
rect 372436 375284 372488 375290
rect 372436 375226 372488 375232
rect 373172 358148 373224 358154
rect 373172 358090 373224 358096
rect 372436 358080 372488 358086
rect 372436 358022 372488 358028
rect 372344 269748 372396 269754
rect 372344 269690 372396 269696
rect 372252 268524 372304 268530
rect 372252 268466 372304 268472
rect 372448 252006 372476 358022
rect 372528 273624 372580 273630
rect 372528 273566 372580 273572
rect 372436 252000 372488 252006
rect 372436 251942 372488 251948
rect 372160 163192 372212 163198
rect 372160 163134 372212 163140
rect 372068 148436 372120 148442
rect 372068 148378 372120 148384
rect 371790 146296 371846 146305
rect 371790 146231 371846 146240
rect 372540 145897 372568 273566
rect 373184 273426 373212 358090
rect 373172 273420 373224 273426
rect 373172 273362 373224 273368
rect 373184 148374 373212 273362
rect 373172 148368 373224 148374
rect 373172 148310 373224 148316
rect 372526 145888 372582 145897
rect 372526 145823 372582 145832
rect 371700 145512 371752 145518
rect 371700 145454 371752 145460
rect 370504 70372 370556 70378
rect 370504 70314 370556 70320
rect 367744 57452 367796 57458
rect 367744 57394 367796 57400
rect 373276 57322 373304 465695
rect 373368 166394 373396 469882
rect 373448 465860 373500 465866
rect 373448 465802 373500 465808
rect 373356 166388 373408 166394
rect 373356 166330 373408 166336
rect 373460 165034 373488 465802
rect 373552 271182 373580 489262
rect 374460 484152 374512 484158
rect 374460 484094 374512 484100
rect 373632 479732 373684 479738
rect 373632 479674 373684 479680
rect 373540 271176 373592 271182
rect 373540 271118 373592 271124
rect 373644 271046 373672 479674
rect 373724 473000 373776 473006
rect 373724 472942 373776 472948
rect 373736 272746 373764 472942
rect 373816 378412 373868 378418
rect 373816 378354 373868 378360
rect 373724 272740 373776 272746
rect 373724 272682 373776 272688
rect 373632 271040 373684 271046
rect 373632 270982 373684 270988
rect 373828 269890 373856 378354
rect 373906 377904 373962 377913
rect 373906 377839 373962 377848
rect 373816 269884 373868 269890
rect 373816 269826 373868 269832
rect 373632 269204 373684 269210
rect 373632 269146 373684 269152
rect 373540 269068 373592 269074
rect 373540 269010 373592 269016
rect 373552 268394 373580 269010
rect 373540 268388 373592 268394
rect 373540 268330 373592 268336
rect 373448 165028 373500 165034
rect 373448 164970 373500 164976
rect 373552 162178 373580 268330
rect 373540 162172 373592 162178
rect 373540 162114 373592 162120
rect 373356 148436 373408 148442
rect 373356 148378 373408 148384
rect 373264 57316 373316 57322
rect 373264 57258 373316 57264
rect 373368 55826 373396 148378
rect 373448 145512 373500 145518
rect 373448 145454 373500 145460
rect 373460 59362 373488 145454
rect 373644 144906 373672 269146
rect 373724 269136 373776 269142
rect 373724 269078 373776 269084
rect 373632 144900 373684 144906
rect 373632 144842 373684 144848
rect 373736 144838 373764 269078
rect 373724 144832 373776 144838
rect 373724 144774 373776 144780
rect 373448 59356 373500 59362
rect 373448 59298 373500 59304
rect 373920 57866 373948 377839
rect 374472 376514 374500 484094
rect 374552 471436 374604 471442
rect 374552 471378 374604 471384
rect 374564 378826 374592 471378
rect 374552 378820 374604 378826
rect 374552 378762 374604 378768
rect 374460 376508 374512 376514
rect 374460 376450 374512 376456
rect 374460 374944 374512 374950
rect 374460 374886 374512 374892
rect 374472 273222 374500 374886
rect 374460 273216 374512 273222
rect 374460 273158 374512 273164
rect 374564 272490 374592 378762
rect 374380 272462 374592 272490
rect 374380 271289 374408 272462
rect 374460 272332 374512 272338
rect 374460 272274 374512 272280
rect 374366 271280 374422 271289
rect 374366 271215 374422 271224
rect 374380 163742 374408 271215
rect 374472 268802 374500 272274
rect 374552 269544 374604 269550
rect 374552 269486 374604 269492
rect 374460 268796 374512 268802
rect 374460 268738 374512 268744
rect 374368 163736 374420 163742
rect 374368 163678 374420 163684
rect 374276 163192 374328 163198
rect 374276 163134 374328 163140
rect 373908 57860 373960 57866
rect 373908 57802 373960 57808
rect 374288 56438 374316 163134
rect 374472 162722 374500 268738
rect 374564 163810 374592 269486
rect 374552 163804 374604 163810
rect 374552 163746 374604 163752
rect 374460 162716 374512 162722
rect 374460 162658 374512 162664
rect 374472 151814 374500 162658
rect 374380 151786 374500 151814
rect 374380 59022 374408 151786
rect 374552 148368 374604 148374
rect 374552 148310 374604 148316
rect 374460 146192 374512 146198
rect 374460 146134 374512 146140
rect 374368 59016 374420 59022
rect 374368 58958 374420 58964
rect 374276 56432 374328 56438
rect 374276 56374 374328 56380
rect 374472 55894 374500 146134
rect 374564 56506 374592 148310
rect 374656 59294 374684 490554
rect 376024 489184 376076 489190
rect 376024 489126 376076 489132
rect 374828 486464 374880 486470
rect 374828 486406 374880 486412
rect 374736 472660 374788 472666
rect 374736 472602 374788 472608
rect 374644 59288 374696 59294
rect 374644 59230 374696 59236
rect 374748 57390 374776 472602
rect 374840 165345 374868 486406
rect 375012 482452 375064 482458
rect 375012 482394 375064 482400
rect 374920 465724 374972 465730
rect 374920 465666 374972 465672
rect 374932 166258 374960 465666
rect 375024 270978 375052 482394
rect 375196 473068 375248 473074
rect 375196 473010 375248 473016
rect 375104 468512 375156 468518
rect 375104 468454 375156 468460
rect 375116 271114 375144 468454
rect 375208 379370 375236 473010
rect 375932 471708 375984 471714
rect 375932 471650 375984 471656
rect 375288 471504 375340 471510
rect 375288 471446 375340 471452
rect 375300 379846 375328 471446
rect 375840 467696 375892 467702
rect 375840 467638 375892 467644
rect 375288 379840 375340 379846
rect 375288 379782 375340 379788
rect 375196 379364 375248 379370
rect 375196 379306 375248 379312
rect 375194 376000 375250 376009
rect 375194 375935 375250 375944
rect 375208 272338 375236 375935
rect 375196 272332 375248 272338
rect 375196 272274 375248 272280
rect 375300 272218 375328 379782
rect 375852 375902 375880 467638
rect 375840 375896 375892 375902
rect 375840 375838 375892 375844
rect 375944 375358 375972 471650
rect 375932 375352 375984 375358
rect 375932 375294 375984 375300
rect 375932 358420 375984 358426
rect 375932 358362 375984 358368
rect 375208 272190 375328 272218
rect 375104 271108 375156 271114
rect 375104 271050 375156 271056
rect 375012 270972 375064 270978
rect 375012 270914 375064 270920
rect 375010 270464 375066 270473
rect 375010 270399 375066 270408
rect 374920 166252 374972 166258
rect 374920 166194 374972 166200
rect 374826 165336 374882 165345
rect 374826 165271 374882 165280
rect 375024 162790 375052 270399
rect 375104 269612 375156 269618
rect 375104 269554 375156 269560
rect 375116 162858 375144 269554
rect 375208 269142 375236 272190
rect 375944 270473 375972 358362
rect 375930 270464 375986 270473
rect 375930 270399 375986 270408
rect 375748 270088 375800 270094
rect 375748 270030 375800 270036
rect 375288 269748 375340 269754
rect 375288 269690 375340 269696
rect 375196 269136 375248 269142
rect 375196 269078 375248 269084
rect 375196 163600 375248 163606
rect 375196 163542 375248 163548
rect 375208 163198 375236 163542
rect 375196 163192 375248 163198
rect 375196 163134 375248 163140
rect 375104 162852 375156 162858
rect 375104 162794 375156 162800
rect 375012 162784 375064 162790
rect 375012 162726 375064 162732
rect 374920 148640 374972 148646
rect 374920 148582 374972 148588
rect 374828 147552 374880 147558
rect 374828 147494 374880 147500
rect 374736 57384 374788 57390
rect 374736 57326 374788 57332
rect 374552 56500 374604 56506
rect 374552 56442 374604 56448
rect 374460 55888 374512 55894
rect 374460 55830 374512 55836
rect 373356 55820 373408 55826
rect 373356 55762 373408 55768
rect 374840 54466 374868 147494
rect 374932 54534 374960 148582
rect 375024 56574 375052 162726
rect 375196 162172 375248 162178
rect 375196 162114 375248 162120
rect 375012 56568 375064 56574
rect 375012 56510 375064 56516
rect 375208 55078 375236 162114
rect 375300 148986 375328 269690
rect 375288 148980 375340 148986
rect 375288 148922 375340 148928
rect 375300 148646 375328 148922
rect 375288 148640 375340 148646
rect 375288 148582 375340 148588
rect 375288 148504 375340 148510
rect 375288 148446 375340 148452
rect 375300 147558 375328 148446
rect 375288 147552 375340 147558
rect 375288 147494 375340 147500
rect 375760 146198 375788 270030
rect 375840 269884 375892 269890
rect 375840 269826 375892 269832
rect 375852 267734 375880 269826
rect 375852 267706 375972 267734
rect 375840 163532 375892 163538
rect 375840 163474 375892 163480
rect 375748 146192 375800 146198
rect 375748 146134 375800 146140
rect 375760 145790 375788 146134
rect 375748 145784 375800 145790
rect 375748 145726 375800 145732
rect 375852 55214 375880 163474
rect 375944 146198 375972 267706
rect 375932 146192 375984 146198
rect 375932 146134 375984 146140
rect 375932 146056 375984 146062
rect 375932 145998 375984 146004
rect 375944 56030 375972 145998
rect 376036 68105 376064 489126
rect 376576 484084 376628 484090
rect 376576 484026 376628 484032
rect 376116 479664 376168 479670
rect 376116 479606 376168 479612
rect 376128 164694 376156 479606
rect 376300 475448 376352 475454
rect 376300 475390 376352 475396
rect 376208 474020 376260 474026
rect 376208 473962 376260 473968
rect 376220 165481 376248 473962
rect 376312 272678 376340 475390
rect 376392 472932 376444 472938
rect 376392 472874 376444 472880
rect 376300 272672 376352 272678
rect 376300 272614 376352 272620
rect 376404 271658 376432 472874
rect 376484 380656 376536 380662
rect 376484 380598 376536 380604
rect 376496 379642 376524 380598
rect 376484 379636 376536 379642
rect 376484 379578 376536 379584
rect 376484 378616 376536 378622
rect 376484 378558 376536 378564
rect 376392 271652 376444 271658
rect 376392 271594 376444 271600
rect 376496 270230 376524 378558
rect 376588 378010 376616 484026
rect 377312 483948 377364 483954
rect 377312 483890 377364 483896
rect 376760 470280 376812 470286
rect 376760 470222 376812 470228
rect 376772 410553 376800 470222
rect 377220 468648 377272 468654
rect 377220 468590 377272 468596
rect 377128 467560 377180 467566
rect 377128 467502 377180 467508
rect 377034 417888 377090 417897
rect 377034 417823 377090 417832
rect 377048 417450 377076 417823
rect 377036 417444 377088 417450
rect 377036 417386 377088 417392
rect 377034 412040 377090 412049
rect 377034 411975 377090 411984
rect 377048 411942 377076 411975
rect 377036 411936 377088 411942
rect 377036 411878 377088 411884
rect 376758 410544 376814 410553
rect 376758 410479 376814 410488
rect 376852 391944 376904 391950
rect 376852 391886 376904 391892
rect 376864 390969 376892 391886
rect 376850 390960 376906 390969
rect 376850 390895 376906 390904
rect 376944 390516 376996 390522
rect 376944 390458 376996 390464
rect 376956 389337 376984 390458
rect 376942 389328 376998 389337
rect 376942 389263 376998 389272
rect 376944 389156 376996 389162
rect 376944 389098 376996 389104
rect 376956 389065 376984 389098
rect 376942 389056 376998 389065
rect 376942 388991 376998 389000
rect 377140 380662 377168 467502
rect 377128 380656 377180 380662
rect 377128 380598 377180 380604
rect 376668 379636 376720 379642
rect 376668 379578 376720 379584
rect 376576 378004 376628 378010
rect 376576 377946 376628 377952
rect 376576 375012 376628 375018
rect 376576 374954 376628 374960
rect 376484 270224 376536 270230
rect 376484 270166 376536 270172
rect 376390 269920 376446 269929
rect 376390 269855 376446 269864
rect 376404 267734 376432 269855
rect 376496 269210 376524 270166
rect 376588 269618 376616 374954
rect 376680 269958 376708 379578
rect 377232 377534 377260 468590
rect 377324 380730 377352 483890
rect 378784 483676 378836 483682
rect 378784 483618 378836 483624
rect 378232 470348 378284 470354
rect 378232 470290 378284 470296
rect 377404 470144 377456 470150
rect 377404 470086 377456 470092
rect 377416 422294 377444 470086
rect 377772 468920 377824 468926
rect 377772 468862 377824 468868
rect 377416 422266 377720 422294
rect 377588 417444 377640 417450
rect 377588 417386 377640 417392
rect 377494 412040 377550 412049
rect 377494 411975 377550 411984
rect 377402 410952 377458 410961
rect 377402 410887 377458 410896
rect 377416 410582 377444 410887
rect 377404 410576 377456 410582
rect 377404 410518 377456 410524
rect 377402 409184 377458 409193
rect 377402 409119 377404 409128
rect 377456 409119 377458 409128
rect 377404 409090 377456 409096
rect 377312 380724 377364 380730
rect 377312 380666 377364 380672
rect 377220 377528 377272 377534
rect 377220 377470 377272 377476
rect 376760 375352 376812 375358
rect 376758 375320 376760 375329
rect 376812 375320 376814 375329
rect 376758 375255 376814 375264
rect 377220 375216 377272 375222
rect 377220 375158 377272 375164
rect 377036 375148 377088 375154
rect 377036 375090 377088 375096
rect 377128 375148 377180 375154
rect 377128 375090 377180 375096
rect 377048 374882 377076 375090
rect 377036 374876 377088 374882
rect 377036 374818 377088 374824
rect 376942 310856 376998 310865
rect 376942 310791 376998 310800
rect 376956 287054 376984 310791
rect 376864 287026 376984 287054
rect 376760 282872 376812 282878
rect 376760 282814 376812 282820
rect 376772 282169 376800 282814
rect 376758 282160 376814 282169
rect 376758 282095 376814 282104
rect 376864 277394 376892 287026
rect 376944 284300 376996 284306
rect 376944 284242 376996 284248
rect 376956 284073 376984 284242
rect 376942 284064 376998 284073
rect 376942 283999 376998 284008
rect 376942 282296 376998 282305
rect 376942 282231 376998 282240
rect 376956 281586 376984 282231
rect 376944 281580 376996 281586
rect 376944 281522 376996 281528
rect 376864 277366 376984 277394
rect 376668 269952 376720 269958
rect 376668 269894 376720 269900
rect 376576 269612 376628 269618
rect 376576 269554 376628 269560
rect 376484 269204 376536 269210
rect 376484 269146 376536 269152
rect 376760 269068 376812 269074
rect 376760 269010 376812 269016
rect 376576 268864 376628 268870
rect 376576 268806 376628 268812
rect 376404 267706 376524 267734
rect 376392 252000 376444 252006
rect 376392 251942 376444 251948
rect 376206 165472 376262 165481
rect 376206 165407 376262 165416
rect 376116 164688 376168 164694
rect 376116 164630 376168 164636
rect 376404 164082 376432 251942
rect 376392 164076 376444 164082
rect 376392 164018 376444 164024
rect 376300 146192 376352 146198
rect 376300 146134 376352 146140
rect 376312 145994 376340 146134
rect 376300 145988 376352 145994
rect 376300 145930 376352 145936
rect 376206 145752 376262 145761
rect 376206 145687 376262 145696
rect 376116 144832 376168 144838
rect 376116 144774 376168 144780
rect 376022 68096 376078 68105
rect 376022 68031 376078 68040
rect 375932 56024 375984 56030
rect 375932 55966 375984 55972
rect 375840 55208 375892 55214
rect 375840 55150 375892 55156
rect 375196 55072 375248 55078
rect 375196 55014 375248 55020
rect 376128 54670 376156 144774
rect 376220 56234 376248 145687
rect 376208 56228 376260 56234
rect 376208 56170 376260 56176
rect 376312 54738 376340 145930
rect 376404 56370 376432 164018
rect 376496 162450 376524 267706
rect 376484 162444 376536 162450
rect 376484 162386 376536 162392
rect 376392 56364 376444 56370
rect 376392 56306 376444 56312
rect 376496 55146 376524 162386
rect 376588 161474 376616 268806
rect 376772 162518 376800 269010
rect 376956 203969 376984 277366
rect 377048 272406 377076 374818
rect 377140 374814 377168 375090
rect 377128 374808 377180 374814
rect 377128 374750 377180 374756
rect 377036 272400 377088 272406
rect 377036 272342 377088 272348
rect 377036 270292 377088 270298
rect 377036 270234 377088 270240
rect 376942 203960 376998 203969
rect 376942 203895 376998 203904
rect 376850 198792 376906 198801
rect 376850 198727 376906 198736
rect 376760 162512 376812 162518
rect 376760 162454 376812 162460
rect 376668 161492 376720 161498
rect 376588 161446 376668 161474
rect 376668 161434 376720 161440
rect 376574 146296 376630 146305
rect 376574 146231 376630 146240
rect 376588 145761 376616 146231
rect 376574 145752 376630 145761
rect 376574 145687 376630 145696
rect 376576 145580 376628 145586
rect 376576 145522 376628 145528
rect 376588 144838 376616 145522
rect 376576 144832 376628 144838
rect 376576 144774 376628 144780
rect 376680 59498 376708 161434
rect 376864 92857 376892 198727
rect 376956 176746 376984 203895
rect 377048 190454 377076 270234
rect 377140 269074 377168 374750
rect 377232 269074 377260 375158
rect 377508 305017 377536 411975
rect 377600 310865 377628 417386
rect 377692 416514 377720 422266
rect 377784 416945 377812 468862
rect 378140 468444 378192 468450
rect 378140 468386 378192 468392
rect 377770 416936 377826 416945
rect 377770 416871 377826 416880
rect 378046 416936 378102 416945
rect 378046 416871 378102 416880
rect 377692 416486 377812 416514
rect 377784 414769 377812 416486
rect 377770 414760 377826 414769
rect 377770 414695 377826 414704
rect 377678 413808 377734 413817
rect 377678 413743 377734 413752
rect 377692 413302 377720 413743
rect 377680 413296 377732 413302
rect 377680 413238 377732 413244
rect 377586 310856 377642 310865
rect 377586 310791 377642 310800
rect 377692 306785 377720 413238
rect 377784 307873 377812 414695
rect 377864 410576 377916 410582
rect 377864 410518 377916 410524
rect 377770 307864 377826 307873
rect 377770 307799 377826 307808
rect 377678 306776 377734 306785
rect 377678 306711 377734 306720
rect 377692 306374 377720 306711
rect 377600 306346 377720 306374
rect 377494 305008 377550 305017
rect 377494 304943 377550 304952
rect 377310 302152 377366 302161
rect 377310 302087 377366 302096
rect 377128 269068 377180 269074
rect 377128 269010 377180 269016
rect 377220 269068 377272 269074
rect 377220 269010 377272 269016
rect 377324 195265 377352 302087
rect 377508 198121 377536 304943
rect 377600 199889 377628 306346
rect 377678 303648 377734 303657
rect 377678 303583 377734 303592
rect 377586 199880 377642 199889
rect 377586 199815 377642 199824
rect 377600 198801 377628 199815
rect 377586 198792 377642 198801
rect 377586 198727 377642 198736
rect 377494 198112 377550 198121
rect 377494 198047 377550 198056
rect 377310 195256 377366 195265
rect 377310 195191 377366 195200
rect 377048 190426 377168 190454
rect 377036 178016 377088 178022
rect 377036 177958 377088 177964
rect 377048 177041 377076 177958
rect 377034 177032 377090 177041
rect 377034 176967 377090 176976
rect 376956 176718 377076 176746
rect 376944 176656 376996 176662
rect 376944 176598 376996 176604
rect 376956 175409 376984 176598
rect 376942 175400 376998 175409
rect 376942 175335 376998 175344
rect 377048 175250 377076 176718
rect 376956 175222 377076 175250
rect 376956 96937 376984 175222
rect 377140 161474 377168 190426
rect 377220 175228 377272 175234
rect 377220 175170 377272 175176
rect 377232 175137 377260 175170
rect 377218 175128 377274 175137
rect 377218 175063 377274 175072
rect 377312 164212 377364 164218
rect 377312 164154 377364 164160
rect 377324 163441 377352 164154
rect 377310 163432 377366 163441
rect 377310 163367 377366 163376
rect 377324 163033 377352 163367
rect 377310 163024 377366 163033
rect 377310 162959 377366 162968
rect 377048 161446 377168 161474
rect 377048 145314 377076 161446
rect 377312 145920 377364 145926
rect 377312 145862 377364 145868
rect 377036 145308 377088 145314
rect 377036 145250 377088 145256
rect 377048 142154 377076 145250
rect 377048 142126 377260 142154
rect 376942 96928 376998 96937
rect 376942 96863 376998 96872
rect 376850 92848 376906 92857
rect 376850 92783 376906 92792
rect 376944 70372 376996 70378
rect 376944 70314 376996 70320
rect 376956 70009 376984 70314
rect 376942 70000 376998 70009
rect 376942 69935 376998 69944
rect 376942 68368 376998 68377
rect 376942 68303 376944 68312
rect 376996 68303 376998 68312
rect 376944 68274 376996 68280
rect 376668 59492 376720 59498
rect 376668 59434 376720 59440
rect 376484 55140 376536 55146
rect 376484 55082 376536 55088
rect 377232 54874 377260 142126
rect 377220 54868 377272 54874
rect 377220 54810 377272 54816
rect 377324 54806 377352 145862
rect 377508 91089 377536 198047
rect 377692 197033 377720 303583
rect 377784 200841 377812 307799
rect 377876 303929 377904 410518
rect 377954 409184 378010 409193
rect 377954 409119 378010 409128
rect 377862 303920 377918 303929
rect 377862 303855 377918 303864
rect 377876 303657 377904 303855
rect 377862 303648 377918 303657
rect 377862 303583 377918 303592
rect 377968 302161 377996 409119
rect 378060 310049 378088 416871
rect 378152 398138 378180 468386
rect 378140 398132 378192 398138
rect 378140 398074 378192 398080
rect 378140 383988 378192 383994
rect 378140 383930 378192 383936
rect 378152 376786 378180 383930
rect 378244 379545 378272 470290
rect 378324 398132 378376 398138
rect 378324 398074 378376 398080
rect 378336 383994 378364 398074
rect 378324 383988 378376 383994
rect 378324 383930 378376 383936
rect 378230 379536 378286 379545
rect 378230 379471 378286 379480
rect 378244 379438 378272 379471
rect 378232 379432 378284 379438
rect 378232 379374 378284 379380
rect 378140 376780 378192 376786
rect 378140 376722 378192 376728
rect 378600 376780 378652 376786
rect 378600 376722 378652 376728
rect 378612 376106 378640 376722
rect 378600 376100 378652 376106
rect 378600 376042 378652 376048
rect 378140 375284 378192 375290
rect 378140 375226 378192 375232
rect 378152 374814 378180 375226
rect 378692 375080 378744 375086
rect 378692 375022 378744 375028
rect 378140 374808 378192 374814
rect 378140 374750 378192 374756
rect 378046 310040 378102 310049
rect 378046 309975 378102 309984
rect 377954 302152 378010 302161
rect 377954 302087 378010 302096
rect 377956 268252 378008 268258
rect 377956 268194 378008 268200
rect 377862 203008 377918 203017
rect 377862 202943 377918 202952
rect 377770 200832 377826 200841
rect 377770 200767 377826 200776
rect 377678 197024 377734 197033
rect 377678 196959 377734 196968
rect 377586 195256 377642 195265
rect 377586 195191 377642 195200
rect 377494 91080 377550 91089
rect 377494 91015 377550 91024
rect 377600 88233 377628 195191
rect 377692 90001 377720 196959
rect 377784 93809 377812 200767
rect 377876 95985 377904 202943
rect 377968 146062 377996 268194
rect 378060 203017 378088 309975
rect 378152 273562 378180 374750
rect 378140 273556 378192 273562
rect 378140 273498 378192 273504
rect 378600 273556 378652 273562
rect 378600 273498 378652 273504
rect 378612 273086 378640 273498
rect 378600 273080 378652 273086
rect 378600 273022 378652 273028
rect 378600 270428 378652 270434
rect 378600 270370 378652 270376
rect 378046 203008 378102 203017
rect 378046 202943 378102 202952
rect 378046 162616 378102 162625
rect 378102 162574 378180 162602
rect 378046 162551 378102 162560
rect 378152 162518 378180 162574
rect 378048 162512 378100 162518
rect 378048 162454 378100 162460
rect 378140 162512 378192 162518
rect 378140 162454 378192 162460
rect 378060 161566 378088 162454
rect 378048 161560 378100 161566
rect 378048 161502 378100 161508
rect 377956 146056 378008 146062
rect 377956 145998 378008 146004
rect 377968 145858 377996 145998
rect 377956 145852 378008 145858
rect 377956 145794 378008 145800
rect 377862 95976 377918 95985
rect 377862 95911 377918 95920
rect 377770 93800 377826 93809
rect 377770 93735 377826 93744
rect 377678 89992 377734 90001
rect 377678 89927 377734 89936
rect 377586 88224 377642 88233
rect 377586 88159 377642 88168
rect 378060 59566 378088 161502
rect 378612 161474 378640 270370
rect 378704 269006 378732 375022
rect 378692 269000 378744 269006
rect 378692 268942 378744 268948
rect 378704 268870 378732 268942
rect 378692 268864 378744 268870
rect 378692 268806 378744 268812
rect 378796 164762 378824 483618
rect 378876 482316 378928 482322
rect 378876 482258 378928 482264
rect 378888 164830 378916 482258
rect 434824 478174 434852 596663
rect 434916 544921 434944 653346
rect 494072 649330 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 542372 654838 542400 702406
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 542360 654832 542412 654838
rect 542360 654774 542412 654780
rect 494060 649324 494112 649330
rect 494060 649266 494112 649272
rect 457444 647284 457496 647290
rect 457444 647226 457496 647232
rect 436192 646468 436244 646474
rect 436192 646410 436244 646416
rect 436100 646400 436152 646406
rect 436100 646342 436152 646348
rect 436112 621761 436140 646342
rect 436204 626521 436232 646410
rect 436284 646332 436336 646338
rect 436284 646274 436336 646280
rect 436296 636041 436324 646274
rect 456984 645040 457036 645046
rect 456984 644982 457036 644988
rect 456996 639713 457024 644982
rect 456982 639704 457038 639713
rect 456982 639639 457038 639648
rect 436282 636032 436338 636041
rect 436282 635967 436338 635976
rect 436190 626512 436246 626521
rect 436190 626447 436246 626456
rect 436098 621752 436154 621761
rect 436098 621687 436154 621696
rect 436742 615904 436798 615913
rect 436742 615839 436798 615848
rect 436190 592104 436246 592113
rect 436190 592039 436246 592048
rect 436098 553480 436154 553489
rect 436098 553415 436154 553424
rect 434902 544912 434958 544921
rect 434902 544847 434958 544856
rect 436112 534002 436140 553415
rect 436204 542994 436232 592039
rect 436282 581768 436338 581777
rect 436282 581703 436338 581712
rect 436296 543114 436324 581703
rect 436374 577280 436430 577289
rect 436374 577215 436430 577224
rect 436284 543108 436336 543114
rect 436284 543050 436336 543056
rect 436204 542966 436324 542994
rect 436296 534070 436324 542966
rect 436284 534064 436336 534070
rect 436284 534006 436336 534012
rect 436100 533996 436152 534002
rect 436100 533938 436152 533944
rect 436388 533866 436416 577215
rect 436466 567624 436522 567633
rect 436466 567559 436522 567568
rect 436376 533860 436428 533866
rect 436376 533802 436428 533808
rect 436480 530806 436508 567559
rect 436558 563136 436614 563145
rect 436558 563071 436614 563080
rect 436572 535430 436600 563071
rect 436650 558104 436706 558113
rect 436650 558039 436706 558048
rect 436664 542994 436692 558039
rect 436756 543130 436784 615839
rect 457456 602313 457484 647226
rect 457536 646196 457588 646202
rect 457536 646138 457588 646144
rect 457548 621353 457576 646138
rect 494796 646128 494848 646134
rect 494796 646070 494848 646076
rect 457720 645108 457772 645114
rect 457720 645050 457772 645056
rect 457628 644904 457680 644910
rect 457628 644846 457680 644852
rect 457640 627473 457668 644846
rect 457732 633593 457760 645050
rect 471612 644972 471664 644978
rect 471612 644914 471664 644920
rect 465172 640348 465224 640354
rect 465172 640290 465224 640296
rect 465184 639963 465212 640290
rect 471624 639963 471652 644914
rect 483204 644836 483256 644842
rect 483204 644778 483256 644784
rect 477130 639976 477186 639985
rect 483216 639963 483244 644778
rect 488722 639976 488778 639985
rect 477186 639934 477434 639962
rect 477130 639911 477186 639920
rect 494808 639963 494836 646070
rect 580356 645176 580408 645182
rect 580356 645118 580408 645124
rect 512000 644768 512052 644774
rect 512000 644710 512052 644716
rect 501236 644564 501288 644570
rect 501236 644506 501288 644512
rect 501248 639963 501276 644506
rect 506754 639976 506810 639985
rect 488778 639934 489026 639962
rect 488722 639911 488778 639920
rect 506810 639934 507058 639962
rect 506754 639911 506810 639920
rect 457718 633584 457774 633593
rect 457718 633519 457774 633528
rect 457626 627464 457682 627473
rect 457626 627399 457682 627408
rect 512012 624073 512040 644710
rect 512092 644700 512144 644706
rect 512092 644642 512144 644648
rect 512104 630873 512132 644642
rect 512184 644632 512236 644638
rect 512184 644574 512236 644580
rect 512196 636993 512224 644574
rect 580264 640348 580316 640354
rect 580264 640290 580316 640296
rect 512182 636984 512238 636993
rect 512182 636919 512238 636928
rect 512090 630864 512146 630873
rect 512090 630799 512146 630808
rect 511998 624064 512054 624073
rect 511998 623999 512054 624008
rect 457534 621344 457590 621353
rect 457534 621279 457590 621288
rect 512090 617944 512146 617953
rect 512090 617879 512146 617888
rect 457626 614544 457682 614553
rect 457626 614479 457682 614488
rect 457534 608424 457590 608433
rect 457534 608359 457590 608368
rect 457442 602304 457498 602313
rect 457442 602239 457498 602248
rect 457442 596184 457498 596193
rect 457442 596119 457498 596128
rect 436834 548448 436890 548457
rect 436834 548383 436890 548392
rect 436848 543250 436876 548383
rect 436836 543244 436888 543250
rect 436836 543186 436888 543192
rect 436756 543102 436968 543130
rect 436836 543040 436888 543046
rect 436664 542966 436784 542994
rect 436836 542982 436888 542988
rect 436652 542904 436704 542910
rect 436652 542846 436704 542852
rect 436560 535424 436612 535430
rect 436560 535366 436612 535372
rect 436664 533526 436692 542846
rect 436756 533662 436784 542966
rect 436848 533934 436876 542982
rect 436836 533928 436888 533934
rect 436836 533870 436888 533876
rect 436744 533656 436796 533662
rect 436744 533598 436796 533604
rect 436940 533594 436968 543102
rect 436928 533588 436980 533594
rect 436928 533530 436980 533536
rect 436652 533520 436704 533526
rect 436652 533462 436704 533468
rect 457456 530942 457484 596119
rect 457444 530936 457496 530942
rect 457444 530878 457496 530884
rect 436468 530800 436520 530806
rect 436468 530742 436520 530748
rect 457548 480865 457576 608359
rect 457640 530874 457668 614479
rect 511998 605704 512054 605713
rect 511998 605639 512054 605648
rect 459572 590022 460046 590050
rect 465092 590022 465842 590050
rect 470612 590022 471638 590050
rect 476132 590022 477434 590050
rect 483032 590022 483230 590050
rect 488552 590022 489670 590050
rect 459572 531078 459600 590022
rect 459560 531072 459612 531078
rect 459560 531014 459612 531020
rect 457628 530868 457680 530874
rect 457628 530810 457680 530816
rect 465092 529718 465120 590022
rect 470612 529786 470640 590022
rect 476132 531010 476160 590022
rect 476120 531004 476172 531010
rect 476120 530946 476172 530952
rect 470600 529780 470652 529786
rect 470600 529722 470652 529728
rect 465080 529712 465132 529718
rect 465080 529654 465132 529660
rect 483032 493377 483060 590022
rect 488552 531146 488580 590022
rect 495452 531282 495480 590036
rect 500972 590022 501262 590050
rect 506492 590022 507058 590050
rect 495440 531276 495492 531282
rect 495440 531218 495492 531224
rect 488540 531140 488592 531146
rect 488540 531082 488592 531088
rect 500972 529854 501000 590022
rect 500960 529848 501012 529854
rect 500960 529790 501012 529796
rect 506492 527882 506520 590022
rect 506480 527876 506532 527882
rect 506480 527818 506532 527824
rect 483018 493368 483074 493377
rect 483018 493303 483074 493312
rect 512012 482225 512040 605639
rect 512104 526425 512132 617879
rect 512182 611824 512238 611833
rect 512182 611759 512238 611768
rect 512196 531214 512224 611759
rect 512274 599584 512330 599593
rect 512274 599519 512330 599528
rect 512184 531208 512236 531214
rect 512184 531150 512236 531156
rect 512288 529922 512316 599519
rect 513286 592784 513342 592793
rect 513286 592719 513342 592728
rect 513300 592074 513328 592719
rect 513288 592068 513340 592074
rect 513288 592010 513340 592016
rect 578884 592068 578936 592074
rect 578884 592010 578936 592016
rect 520924 529984 520976 529990
rect 520924 529926 520976 529932
rect 512276 529916 512328 529922
rect 512276 529858 512328 529864
rect 512090 526416 512146 526425
rect 512090 526351 512146 526360
rect 518164 499588 518216 499594
rect 518164 499530 518216 499536
rect 511998 482216 512054 482225
rect 511998 482151 512054 482160
rect 457534 480856 457590 480865
rect 457534 480791 457590 480800
rect 434812 478168 434864 478174
rect 434812 478110 434864 478116
rect 379244 470212 379296 470218
rect 379244 470154 379296 470160
rect 379060 465928 379112 465934
rect 379060 465870 379112 465876
rect 378968 465792 379020 465798
rect 378968 465734 379020 465740
rect 378980 165306 379008 465734
rect 379072 271697 379100 465870
rect 379256 375290 379284 470154
rect 379980 470076 380032 470082
rect 379980 470018 380032 470024
rect 379992 378962 380020 470018
rect 498476 466676 498528 466682
rect 498476 466618 498528 466624
rect 499488 466676 499540 466682
rect 499488 466618 499540 466624
rect 498488 466585 498516 466618
rect 498474 466576 498530 466585
rect 499500 466546 499528 466618
rect 499764 466608 499816 466614
rect 499762 466576 499764 466585
rect 517888 466608 517940 466614
rect 499816 466576 499818 466585
rect 498474 466511 498530 466520
rect 499488 466540 499540 466546
rect 499762 466511 499818 466520
rect 510894 466576 510950 466585
rect 517888 466550 517940 466556
rect 510894 466511 510896 466520
rect 499488 466482 499540 466488
rect 510948 466511 510950 466520
rect 517520 466540 517572 466546
rect 510896 466482 510948 466488
rect 517520 466482 517572 466488
rect 421104 380928 421156 380934
rect 413558 380896 413614 380905
rect 413558 380831 413614 380840
rect 421102 380896 421104 380905
rect 421156 380896 421158 380905
rect 421102 380831 421158 380840
rect 425978 380896 426034 380905
rect 425978 380831 426034 380840
rect 433614 380896 433670 380905
rect 433614 380831 433670 380840
rect 436006 380896 436062 380905
rect 436006 380831 436062 380840
rect 380992 380792 381044 380798
rect 380992 380734 381044 380740
rect 380898 380216 380954 380225
rect 380898 380151 380954 380160
rect 379612 378956 379664 378962
rect 379612 378898 379664 378904
rect 379980 378956 380032 378962
rect 379980 378898 380032 378904
rect 379520 378888 379572 378894
rect 379520 378830 379572 378836
rect 379532 378418 379560 378830
rect 379624 378486 379652 378898
rect 379612 378480 379664 378486
rect 379612 378422 379664 378428
rect 379520 378412 379572 378418
rect 379520 378354 379572 378360
rect 379336 375896 379388 375902
rect 379336 375838 379388 375844
rect 379244 375284 379296 375290
rect 379244 375226 379296 375232
rect 379256 365090 379284 375226
rect 379244 365084 379296 365090
rect 379244 365026 379296 365032
rect 379348 362386 379376 375838
rect 379428 365084 379480 365090
rect 379428 365026 379480 365032
rect 379164 362358 379376 362386
rect 379058 271688 379114 271697
rect 379058 271623 379114 271632
rect 379060 269068 379112 269074
rect 379060 269010 379112 269016
rect 379072 268462 379100 269010
rect 379164 268802 379192 362358
rect 379440 362250 379468 365026
rect 379256 362222 379468 362250
rect 379256 273630 379284 362222
rect 379428 358760 379480 358766
rect 379428 358702 379480 358708
rect 379336 357536 379388 357542
rect 379336 357478 379388 357484
rect 379244 273624 379296 273630
rect 379244 273566 379296 273572
rect 379256 273154 379284 273566
rect 379244 273148 379296 273154
rect 379244 273090 379296 273096
rect 379348 270502 379376 357478
rect 379440 273562 379468 358702
rect 379428 273556 379480 273562
rect 379428 273498 379480 273504
rect 379426 273320 379482 273329
rect 379426 273255 379482 273264
rect 379336 270496 379388 270502
rect 379336 270438 379388 270444
rect 379244 269068 379296 269074
rect 379244 269010 379296 269016
rect 379256 268870 379284 269010
rect 379244 268864 379296 268870
rect 379244 268806 379296 268812
rect 379152 268796 379204 268802
rect 379152 268738 379204 268744
rect 379060 268456 379112 268462
rect 379060 268398 379112 268404
rect 378968 165300 379020 165306
rect 378968 165242 379020 165248
rect 378876 164824 378928 164830
rect 378876 164766 378928 164772
rect 378784 164756 378836 164762
rect 378784 164698 378836 164704
rect 378612 161446 379008 161474
rect 378876 146192 378928 146198
rect 378876 146134 378928 146140
rect 378414 145888 378470 145897
rect 378414 145823 378470 145832
rect 378048 59560 378100 59566
rect 378048 59502 378100 59508
rect 378428 54942 378456 145823
rect 378888 145722 378916 146134
rect 378980 146062 379008 161446
rect 378968 146056 379020 146062
rect 378968 145998 379020 146004
rect 378876 145716 378928 145722
rect 378876 145658 378928 145664
rect 378784 145648 378836 145654
rect 378784 145590 378836 145596
rect 378600 145444 378652 145450
rect 378600 145386 378652 145392
rect 378612 59702 378640 145386
rect 378692 145376 378744 145382
rect 378692 145318 378744 145324
rect 378704 59770 378732 145318
rect 378796 144906 378824 145590
rect 378784 144900 378836 144906
rect 378784 144842 378836 144848
rect 378692 59764 378744 59770
rect 378692 59706 378744 59712
rect 378600 59696 378652 59702
rect 378600 59638 378652 59644
rect 378416 54936 378468 54942
rect 378416 54878 378468 54884
rect 377312 54800 377364 54806
rect 377312 54742 377364 54748
rect 376300 54732 376352 54738
rect 376300 54674 376352 54680
rect 376116 54664 376168 54670
rect 376116 54606 376168 54612
rect 378796 54602 378824 144842
rect 378888 59634 378916 145658
rect 378980 60722 379008 145998
rect 379072 145926 379100 268398
rect 379164 268258 379192 268738
rect 379244 268524 379296 268530
rect 379244 268466 379296 268472
rect 379152 268252 379204 268258
rect 379152 268194 379204 268200
rect 379152 252068 379204 252074
rect 379152 252010 379204 252016
rect 379164 163878 379192 252010
rect 379152 163872 379204 163878
rect 379152 163814 379204 163820
rect 379060 145920 379112 145926
rect 379060 145862 379112 145868
rect 379058 145616 379114 145625
rect 379058 145551 379114 145560
rect 378968 60716 379020 60722
rect 378968 60658 379020 60664
rect 378966 60616 379022 60625
rect 378966 60551 379022 60560
rect 378876 59628 378928 59634
rect 378876 59570 378928 59576
rect 378980 57798 379008 60551
rect 378968 57792 379020 57798
rect 378968 57734 379020 57740
rect 379072 55010 379100 145551
rect 379164 59226 379192 163814
rect 379256 146198 379284 268466
rect 379336 147688 379388 147694
rect 379336 147630 379388 147636
rect 379244 146192 379296 146198
rect 379244 146134 379296 146140
rect 379244 60716 379296 60722
rect 379244 60658 379296 60664
rect 379152 59220 379204 59226
rect 379152 59162 379204 59168
rect 379256 55962 379284 60658
rect 379348 56098 379376 147630
rect 379440 57594 379468 273255
rect 379532 271028 379560 378354
rect 379624 272066 379652 378422
rect 379888 377460 379940 377466
rect 379888 377402 379940 377408
rect 379796 273556 379848 273562
rect 379796 273498 379848 273504
rect 379704 272400 379756 272406
rect 379704 272342 379756 272348
rect 379612 272060 379664 272066
rect 379612 272002 379664 272008
rect 379716 271998 379744 272342
rect 379704 271992 379756 271998
rect 379704 271934 379756 271940
rect 379532 271000 379652 271028
rect 379520 270496 379572 270502
rect 379520 270438 379572 270444
rect 379532 269822 379560 270438
rect 379624 270434 379652 271000
rect 379612 270428 379664 270434
rect 379612 270370 379664 270376
rect 379520 269816 379572 269822
rect 379520 269758 379572 269764
rect 379532 149054 379560 269758
rect 379624 269618 379652 270370
rect 379612 269612 379664 269618
rect 379612 269554 379664 269560
rect 379716 163946 379744 271934
rect 379808 164014 379836 273498
rect 379900 268870 379928 377402
rect 379992 270502 380020 378898
rect 380912 358766 380940 380151
rect 381004 379778 381032 380734
rect 413572 380730 413600 380831
rect 413560 380724 413612 380730
rect 413560 380666 413612 380672
rect 425992 380662 426020 380831
rect 425980 380656 426032 380662
rect 404174 380624 404230 380633
rect 404174 380559 404230 380568
rect 405462 380624 405518 380633
rect 405462 380559 405518 380568
rect 413466 380624 413522 380633
rect 425980 380598 426032 380604
rect 433628 380594 433656 380831
rect 413466 380559 413522 380568
rect 433616 380588 433668 380594
rect 380992 379772 381044 379778
rect 380992 379714 381044 379720
rect 380900 358760 380952 358766
rect 380900 358702 380952 358708
rect 381004 357542 381032 379714
rect 404188 379710 404216 380559
rect 405476 379846 405504 380559
rect 405464 379840 405516 379846
rect 405464 379782 405516 379788
rect 413480 379778 413508 380559
rect 433616 380530 433668 380536
rect 436020 380526 436048 380831
rect 438490 380760 438546 380769
rect 438490 380695 438546 380704
rect 440882 380760 440938 380769
rect 440882 380695 440938 380704
rect 443458 380760 443514 380769
rect 443458 380695 443514 380704
rect 448242 380760 448298 380769
rect 448242 380695 448298 380704
rect 436008 380520 436060 380526
rect 436008 380462 436060 380468
rect 438504 380458 438532 380695
rect 438492 380452 438544 380458
rect 438492 380394 438544 380400
rect 440896 380390 440924 380695
rect 440884 380384 440936 380390
rect 440884 380326 440936 380332
rect 443472 380254 443500 380695
rect 445942 380624 445998 380633
rect 445942 380559 445998 380568
rect 443460 380248 443512 380254
rect 443460 380190 443512 380196
rect 445956 380186 445984 380559
rect 448256 380322 448284 380695
rect 503350 380624 503406 380633
rect 503350 380559 503406 380568
rect 448244 380316 448296 380322
rect 448244 380258 448296 380264
rect 445944 380180 445996 380186
rect 445944 380122 445996 380128
rect 413468 379772 413520 379778
rect 413468 379714 413520 379720
rect 404176 379704 404228 379710
rect 404176 379646 404228 379652
rect 420644 379636 420696 379642
rect 420644 379578 420696 379584
rect 420656 379409 420684 379578
rect 431132 379568 431184 379574
rect 431132 379510 431184 379516
rect 431144 379409 431172 379510
rect 437940 379500 437992 379506
rect 437940 379442 437992 379448
rect 434260 379432 434312 379438
rect 396078 379400 396134 379409
rect 396078 379335 396134 379344
rect 396354 379400 396410 379409
rect 396354 379335 396410 379344
rect 398194 379400 398250 379409
rect 398194 379335 398250 379344
rect 399482 379400 399538 379409
rect 399482 379335 399538 379344
rect 405830 379400 405886 379409
rect 405830 379335 405886 379344
rect 407578 379400 407634 379409
rect 407578 379335 407634 379344
rect 408314 379400 408370 379409
rect 408314 379335 408316 379344
rect 396092 378962 396120 379335
rect 396080 378956 396132 378962
rect 396080 378898 396132 378904
rect 381082 378856 381138 378865
rect 396368 378826 396396 379335
rect 381082 378791 381138 378800
rect 396356 378820 396408 378826
rect 381096 358086 381124 378791
rect 396356 378762 396408 378768
rect 381174 378720 381230 378729
rect 398208 378690 398236 379335
rect 381174 378655 381230 378664
rect 398196 378684 398248 378690
rect 381188 358154 381216 378655
rect 398196 378626 398248 378632
rect 399496 378554 399524 379335
rect 402978 379264 403034 379273
rect 402978 379199 403034 379208
rect 399484 378548 399536 378554
rect 399484 378490 399536 378496
rect 402992 377398 403020 379199
rect 405844 378622 405872 379335
rect 405832 378616 405884 378622
rect 405832 378558 405884 378564
rect 407592 378350 407620 379335
rect 408368 379335 408370 379344
rect 410338 379400 410394 379409
rect 410338 379335 410394 379344
rect 411258 379400 411314 379409
rect 411258 379335 411314 379344
rect 412362 379400 412418 379409
rect 412362 379335 412418 379344
rect 420642 379400 420698 379409
rect 420642 379335 420698 379344
rect 428186 379400 428242 379409
rect 428186 379335 428242 379344
rect 431130 379400 431186 379409
rect 431130 379335 431186 379344
rect 434258 379400 434260 379409
rect 437952 379409 437980 379442
rect 434312 379400 434314 379409
rect 434258 379335 434314 379344
rect 437938 379400 437994 379409
rect 437938 379335 437994 379344
rect 451002 379400 451058 379409
rect 451002 379335 451058 379344
rect 453026 379400 453082 379409
rect 453026 379335 453082 379344
rect 455602 379400 455658 379409
rect 455602 379335 455658 379344
rect 460938 379400 460994 379409
rect 460938 379335 460994 379344
rect 463514 379400 463570 379409
rect 463514 379335 463570 379344
rect 473450 379400 473506 379409
rect 473450 379335 473506 379344
rect 480626 379400 480682 379409
rect 480626 379335 480682 379344
rect 485962 379400 486018 379409
rect 485962 379335 486018 379344
rect 408316 379306 408368 379312
rect 408682 378584 408738 378593
rect 408682 378519 408738 378528
rect 407580 378344 407632 378350
rect 407580 378286 407632 378292
rect 402980 377392 403032 377398
rect 402980 377334 403032 377340
rect 408696 375902 408724 378519
rect 409970 378176 410026 378185
rect 409970 378111 410026 378120
rect 408684 375896 408736 375902
rect 408684 375838 408736 375844
rect 381266 375320 381322 375329
rect 381266 375255 381322 375264
rect 381280 374649 381308 375255
rect 409984 375222 410012 378111
rect 410352 377534 410380 379335
rect 411272 378418 411300 379335
rect 412376 378486 412404 379335
rect 414570 379264 414626 379273
rect 414570 379199 414626 379208
rect 415858 379264 415914 379273
rect 415858 379199 415914 379208
rect 416042 379264 416098 379273
rect 416042 379199 416098 379208
rect 422850 379264 422906 379273
rect 422850 379199 422906 379208
rect 412364 378480 412416 378486
rect 412364 378422 412416 378428
rect 411260 378412 411312 378418
rect 411260 378354 411312 378360
rect 410340 377528 410392 377534
rect 410340 377470 410392 377476
rect 414584 377466 414612 379199
rect 414572 377460 414624 377466
rect 414572 377402 414624 377408
rect 409972 375216 410024 375222
rect 409972 375158 410024 375164
rect 415872 375154 415900 379199
rect 416056 375970 416084 379199
rect 419354 379128 419410 379137
rect 419354 379063 419410 379072
rect 418434 378584 418490 378593
rect 418434 378519 418490 378528
rect 416962 378176 417018 378185
rect 416962 378111 417018 378120
rect 418158 378176 418214 378185
rect 418158 378111 418214 378120
rect 416044 375964 416096 375970
rect 416044 375906 416096 375912
rect 415860 375148 415912 375154
rect 415860 375090 415912 375096
rect 416976 374950 417004 378111
rect 418172 375018 418200 378111
rect 418448 376174 418476 378519
rect 418436 376168 418488 376174
rect 418436 376110 418488 376116
rect 419368 375086 419396 379063
rect 421746 378584 421802 378593
rect 421746 378519 421802 378528
rect 421760 376009 421788 378519
rect 422574 378312 422630 378321
rect 422574 378247 422630 378256
rect 421746 376000 421802 376009
rect 421746 375935 421802 375944
rect 422588 375358 422616 378247
rect 422864 376310 422892 379199
rect 423954 378176 424010 378185
rect 423954 378111 424010 378120
rect 425150 378176 425206 378185
rect 425150 378111 425206 378120
rect 426438 378176 426494 378185
rect 426438 378111 426494 378120
rect 422852 376304 422904 376310
rect 422852 376246 422904 376252
rect 422576 375352 422628 375358
rect 422576 375294 422628 375300
rect 423968 375290 423996 378111
rect 423956 375284 424008 375290
rect 423956 375226 424008 375232
rect 419356 375080 419408 375086
rect 419356 375022 419408 375028
rect 418160 375012 418212 375018
rect 418160 374954 418212 374960
rect 416964 374944 417016 374950
rect 416964 374886 417016 374892
rect 425164 374882 425192 378111
rect 425152 374876 425204 374882
rect 425152 374818 425204 374824
rect 426452 374814 426480 378111
rect 428200 377602 428228 379335
rect 430670 378584 430726 378593
rect 430670 378519 430726 378528
rect 436190 378584 436246 378593
rect 436190 378519 436246 378528
rect 428278 378176 428334 378185
rect 428278 378111 428334 378120
rect 428188 377596 428240 377602
rect 428188 377538 428240 377544
rect 426440 374808 426492 374814
rect 426440 374750 426492 374756
rect 428292 374746 428320 378111
rect 430684 376242 430712 378519
rect 432234 378176 432290 378185
rect 432234 378111 432290 378120
rect 435178 378176 435234 378185
rect 435178 378111 435234 378120
rect 430672 376236 430724 376242
rect 430672 376178 430724 376184
rect 428280 374740 428332 374746
rect 428280 374682 428332 374688
rect 432248 374678 432276 378111
rect 432236 374672 432288 374678
rect 381266 374640 381322 374649
rect 435192 374649 435220 378111
rect 436204 376106 436232 378519
rect 438122 378176 438178 378185
rect 438122 378111 438178 378120
rect 438136 377913 438164 378111
rect 438122 377904 438178 377913
rect 438122 377839 438178 377848
rect 436192 376100 436244 376106
rect 436192 376042 436244 376048
rect 432236 374614 432288 374620
rect 435178 374640 435234 374649
rect 381266 374575 381322 374584
rect 435178 374575 435234 374584
rect 381280 358426 381308 374575
rect 438136 359582 438164 377839
rect 451016 377670 451044 379335
rect 453040 377738 453068 379335
rect 455616 377806 455644 379335
rect 460952 377942 460980 379335
rect 460940 377936 460992 377942
rect 460940 377878 460992 377884
rect 463528 377874 463556 379335
rect 465078 379128 465134 379137
rect 465078 379063 465134 379072
rect 463516 377868 463568 377874
rect 463516 377810 463568 377816
rect 455604 377800 455656 377806
rect 455604 377742 455656 377748
rect 453028 377732 453080 377738
rect 453028 377674 453080 377680
rect 451004 377664 451056 377670
rect 451004 377606 451056 377612
rect 465092 376378 465120 379063
rect 470874 378992 470930 379001
rect 470874 378927 470930 378936
rect 467930 378856 467986 378865
rect 467930 378791 467986 378800
rect 467944 376446 467972 378791
rect 470888 376718 470916 378927
rect 473464 378146 473492 379335
rect 474738 378856 474794 378865
rect 474738 378791 474794 378800
rect 477498 378856 477554 378865
rect 477498 378791 477554 378800
rect 473452 378140 473504 378146
rect 473452 378082 473504 378088
rect 470876 376712 470928 376718
rect 470876 376654 470928 376660
rect 474752 376650 474780 378791
rect 474740 376644 474792 376650
rect 474740 376586 474792 376592
rect 477512 376582 477540 378791
rect 480640 378078 480668 379335
rect 483386 378856 483442 378865
rect 483386 378791 483442 378800
rect 480628 378072 480680 378078
rect 480628 378014 480680 378020
rect 477500 376576 477552 376582
rect 477500 376518 477552 376524
rect 483400 376514 483428 378791
rect 485976 378010 486004 379335
rect 503364 378214 503392 380559
rect 503626 379400 503682 379409
rect 503626 379335 503682 379344
rect 503640 378758 503668 379335
rect 503628 378752 503680 378758
rect 503628 378694 503680 378700
rect 503640 378282 503668 378694
rect 517532 378418 517560 466482
rect 517796 466472 517848 466478
rect 517796 466414 517848 466420
rect 511908 378412 511960 378418
rect 511908 378354 511960 378360
rect 517520 378412 517572 378418
rect 517520 378354 517572 378360
rect 503628 378276 503680 378282
rect 503628 378218 503680 378224
rect 503352 378208 503404 378214
rect 503352 378150 503404 378156
rect 485964 378004 486016 378010
rect 485964 377946 486016 377952
rect 483388 376508 483440 376514
rect 483388 376450 483440 376456
rect 467932 376440 467984 376446
rect 467932 376382 467984 376388
rect 465080 376372 465132 376378
rect 465080 376314 465132 376320
rect 500776 359712 500828 359718
rect 500776 359654 500828 359660
rect 498844 359644 498896 359650
rect 498844 359586 498896 359592
rect 438124 359576 438176 359582
rect 438124 359518 438176 359524
rect 498856 358873 498884 359586
rect 500788 358873 500816 359654
rect 498842 358864 498898 358873
rect 498842 358799 498898 358808
rect 500774 358864 500830 358873
rect 500774 358799 500830 358808
rect 510894 358864 510950 358873
rect 511920 358834 511948 378354
rect 517612 378276 517664 378282
rect 517612 378218 517664 378224
rect 516600 359576 516652 359582
rect 516600 359518 516652 359524
rect 510894 358799 510896 358808
rect 510948 358799 510950 358808
rect 511908 358828 511960 358834
rect 510896 358770 510948 358776
rect 511908 358770 511960 358776
rect 381268 358420 381320 358426
rect 381268 358362 381320 358368
rect 381176 358148 381228 358154
rect 381176 358090 381228 358096
rect 381084 358080 381136 358086
rect 381084 358022 381136 358028
rect 380992 357536 381044 357542
rect 380992 357478 381044 357484
rect 440882 273728 440938 273737
rect 440882 273663 440938 273672
rect 416042 273592 416098 273601
rect 416042 273527 416098 273536
rect 427634 273592 427690 273601
rect 427634 273527 427636 273536
rect 416056 273494 416084 273527
rect 427688 273527 427690 273536
rect 433338 273592 433394 273601
rect 433338 273527 433394 273536
rect 427636 273498 427688 273504
rect 416044 273488 416096 273494
rect 416044 273430 416096 273436
rect 433352 273426 433380 273527
rect 433340 273420 433392 273426
rect 433340 273362 433392 273368
rect 440896 273358 440924 273663
rect 440884 273352 440936 273358
rect 430946 273320 431002 273329
rect 440884 273294 440936 273300
rect 430946 273255 430948 273264
rect 431000 273255 431002 273264
rect 430948 273226 431000 273232
rect 396724 273216 396776 273222
rect 396724 273158 396776 273164
rect 380072 272060 380124 272066
rect 380072 272002 380124 272008
rect 379980 270496 380032 270502
rect 379980 270438 380032 270444
rect 379992 269550 380020 270438
rect 380084 270434 380112 272002
rect 396736 271153 396764 273158
rect 423772 273148 423824 273154
rect 423772 273090 423824 273096
rect 423404 273012 423456 273018
rect 423404 272954 423456 272960
rect 423416 272921 423444 272954
rect 423784 272921 423812 273090
rect 426440 273080 426492 273086
rect 426440 273022 426492 273028
rect 426452 272921 426480 273022
rect 428188 272944 428240 272950
rect 423402 272912 423458 272921
rect 423402 272847 423458 272856
rect 423770 272912 423826 272921
rect 423770 272847 423826 272856
rect 426438 272912 426494 272921
rect 426438 272847 426494 272856
rect 428186 272912 428188 272921
rect 428240 272912 428242 272921
rect 428186 272847 428242 272856
rect 468482 272912 468538 272921
rect 468482 272847 468484 272856
rect 468536 272847 468538 272856
rect 470874 272912 470930 272921
rect 470874 272847 470930 272856
rect 468484 272818 468536 272824
rect 470888 272814 470916 272847
rect 470876 272808 470928 272814
rect 470876 272750 470928 272756
rect 478418 272776 478474 272785
rect 478418 272711 478420 272720
rect 478472 272711 478474 272720
rect 480810 272776 480866 272785
rect 480810 272711 480866 272720
rect 478420 272682 478472 272688
rect 480824 272678 480852 272711
rect 480812 272672 480864 272678
rect 473450 272640 473506 272649
rect 473450 272575 473506 272584
rect 475842 272640 475898 272649
rect 480812 272614 480864 272620
rect 475842 272575 475844 272584
rect 473464 272542 473492 272575
rect 475896 272575 475898 272584
rect 475844 272546 475896 272552
rect 473452 272536 473504 272542
rect 473452 272478 473504 272484
rect 401690 272232 401746 272241
rect 401690 272167 401746 272176
rect 455786 272232 455842 272241
rect 455786 272167 455842 272176
rect 396722 271144 396778 271153
rect 396722 271079 396778 271088
rect 396078 270600 396134 270609
rect 396078 270535 396134 270544
rect 396092 270502 396120 270535
rect 396080 270496 396132 270502
rect 396080 270438 396132 270444
rect 380072 270428 380124 270434
rect 380072 270370 380124 270376
rect 380084 270298 380112 270370
rect 380072 270292 380124 270298
rect 380072 270234 380124 270240
rect 380256 270224 380308 270230
rect 380256 270166 380308 270172
rect 379980 269544 380032 269550
rect 379980 269486 380032 269492
rect 380268 269142 380296 270166
rect 389180 269952 389232 269958
rect 389180 269894 389232 269900
rect 380256 269136 380308 269142
rect 380256 269078 380308 269084
rect 379888 268864 379940 268870
rect 379888 268806 379940 268812
rect 379900 267734 379928 268806
rect 379900 267706 380020 267734
rect 379796 164008 379848 164014
rect 379796 163950 379848 163956
rect 379704 163940 379756 163946
rect 379704 163882 379756 163888
rect 379612 162852 379664 162858
rect 379612 162794 379664 162800
rect 379624 162246 379652 162794
rect 379612 162240 379664 162246
rect 379612 162182 379664 162188
rect 379520 149048 379572 149054
rect 379520 148990 379572 148996
rect 379532 147694 379560 148990
rect 379520 147688 379572 147694
rect 379520 147630 379572 147636
rect 379624 59158 379652 162182
rect 379612 59152 379664 59158
rect 379612 59094 379664 59100
rect 379716 59090 379744 163882
rect 379704 59084 379756 59090
rect 379704 59026 379756 59032
rect 379428 57588 379480 57594
rect 379428 57530 379480 57536
rect 379808 56302 379836 163950
rect 379888 162784 379940 162790
rect 379888 162726 379940 162732
rect 379900 162450 379928 162726
rect 379888 162444 379940 162450
rect 379888 162386 379940 162392
rect 379992 146130 380020 267706
rect 389192 251841 389220 269894
rect 391940 269680 391992 269686
rect 391940 269622 391992 269628
rect 391952 268734 391980 269622
rect 391940 268728 391992 268734
rect 391940 268670 391992 268676
rect 396736 252074 396764 271079
rect 397458 270600 397514 270609
rect 397458 270535 397514 270544
rect 398838 270600 398894 270609
rect 398838 270535 398894 270544
rect 400218 270600 400274 270609
rect 400218 270535 400274 270544
rect 397472 270162 397500 270535
rect 398852 270366 398880 270535
rect 398840 270360 398892 270366
rect 398840 270302 398892 270308
rect 397460 270156 397512 270162
rect 397460 270098 397512 270104
rect 400232 270026 400260 270535
rect 400220 270020 400272 270026
rect 400220 269962 400272 269968
rect 401704 269754 401732 272167
rect 425060 271992 425112 271998
rect 425060 271934 425112 271940
rect 425072 271833 425100 271934
rect 428004 271924 428056 271930
rect 428004 271866 428056 271872
rect 440148 271924 440200 271930
rect 440148 271866 440200 271872
rect 428016 271833 428044 271866
rect 440160 271833 440188 271866
rect 403530 271824 403586 271833
rect 403530 271759 403586 271768
rect 425058 271824 425114 271833
rect 425058 271759 425114 271768
rect 428002 271824 428058 271833
rect 428002 271759 428058 271768
rect 440146 271824 440202 271833
rect 440146 271759 440202 271768
rect 447138 271824 447194 271833
rect 447138 271759 447194 271768
rect 449898 271824 449954 271833
rect 449898 271759 449954 271768
rect 452658 271824 452714 271833
rect 455800 271794 455828 272167
rect 516612 271930 516640 359518
rect 517520 358828 517572 358834
rect 517520 358770 517572 358776
rect 516600 271924 516652 271930
rect 516600 271866 516652 271872
rect 458180 271856 458232 271862
rect 458178 271824 458180 271833
rect 458232 271824 458234 271833
rect 452658 271759 452714 271768
rect 455788 271788 455840 271794
rect 402978 270600 403034 270609
rect 402978 270535 403034 270544
rect 401692 269748 401744 269754
rect 401692 269690 401744 269696
rect 402992 268530 403020 270535
rect 403544 270094 403572 271759
rect 442998 271552 443054 271561
rect 442998 271487 443000 271496
rect 443052 271487 443054 271496
rect 443000 271458 443052 271464
rect 447152 271454 447180 271759
rect 449912 271726 449940 271759
rect 449900 271720 449952 271726
rect 449900 271662 449952 271668
rect 452672 271590 452700 271759
rect 458178 271759 458234 271768
rect 460938 271824 460994 271833
rect 460938 271759 460994 271768
rect 455788 271730 455840 271736
rect 460952 271658 460980 271759
rect 460940 271652 460992 271658
rect 460940 271594 460992 271600
rect 452660 271584 452712 271590
rect 452660 271526 452712 271532
rect 503626 271552 503682 271561
rect 503626 271487 503682 271496
rect 447140 271448 447192 271454
rect 418342 271416 418398 271425
rect 418342 271351 418398 271360
rect 434718 271416 434774 271425
rect 434718 271351 434774 271360
rect 445758 271416 445814 271425
rect 447140 271390 447192 271396
rect 503534 271416 503590 271425
rect 445758 271351 445760 271360
rect 418356 271046 418384 271351
rect 434732 271318 434760 271351
rect 445812 271351 445814 271360
rect 503534 271351 503590 271360
rect 445760 271322 445812 271328
rect 434720 271312 434772 271318
rect 433338 271280 433394 271289
rect 434720 271254 434772 271260
rect 437478 271280 437534 271289
rect 433338 271215 433394 271224
rect 437478 271215 437534 271224
rect 420918 271144 420974 271153
rect 433352 271114 433380 271215
rect 437492 271182 437520 271215
rect 503548 271182 503576 271351
rect 503640 271318 503668 271487
rect 503628 271312 503680 271318
rect 503628 271254 503680 271260
rect 437480 271176 437532 271182
rect 437480 271118 437532 271124
rect 503536 271176 503588 271182
rect 503536 271118 503588 271124
rect 420918 271079 420920 271088
rect 420972 271079 420974 271088
rect 433340 271108 433392 271114
rect 420920 271050 420972 271056
rect 433340 271050 433392 271056
rect 418344 271040 418396 271046
rect 409878 271008 409934 271017
rect 418344 270982 418396 270988
rect 429198 271008 429254 271017
rect 409878 270943 409880 270952
rect 409932 270943 409934 270952
rect 429198 270943 429254 270952
rect 437478 271008 437534 271017
rect 437478 270943 437534 270952
rect 409880 270914 409932 270920
rect 429212 270910 429240 270943
rect 425704 270904 425756 270910
rect 425704 270846 425756 270852
rect 429200 270904 429252 270910
rect 429200 270846 429252 270852
rect 411350 270736 411406 270745
rect 411350 270671 411406 270680
rect 404358 270600 404414 270609
rect 404358 270535 404414 270544
rect 405738 270600 405794 270609
rect 405738 270535 405794 270544
rect 407118 270600 407174 270609
rect 407118 270535 407174 270544
rect 408498 270600 408554 270609
rect 408498 270535 408554 270544
rect 409878 270600 409934 270609
rect 409878 270535 409934 270544
rect 411258 270600 411314 270609
rect 411258 270535 411314 270544
rect 404372 270230 404400 270535
rect 405752 270298 405780 270535
rect 405740 270292 405792 270298
rect 405740 270234 405792 270240
rect 404360 270224 404412 270230
rect 404360 270166 404412 270172
rect 403532 270088 403584 270094
rect 403532 270030 403584 270036
rect 407132 269890 407160 270535
rect 407120 269884 407172 269890
rect 407120 269826 407172 269832
rect 408512 268802 408540 270535
rect 408500 268796 408552 268802
rect 408500 268738 408552 268744
rect 402980 268524 403032 268530
rect 402980 268466 403032 268472
rect 409892 268462 409920 270535
rect 411272 270434 411300 270535
rect 411260 270428 411312 270434
rect 411260 270370 411312 270376
rect 411364 269618 411392 270671
rect 422944 270632 422996 270638
rect 413006 270600 413062 270609
rect 413006 270535 413062 270544
rect 414018 270600 414074 270609
rect 414018 270535 414074 270544
rect 415398 270600 415454 270609
rect 415398 270535 415454 270544
rect 418158 270600 418214 270609
rect 418158 270535 418214 270544
rect 418526 270600 418582 270609
rect 418526 270535 418582 270544
rect 419538 270600 419594 270609
rect 419538 270535 419594 270544
rect 420918 270600 420974 270609
rect 422944 270574 422996 270580
rect 420918 270535 420974 270544
rect 421564 270564 421616 270570
rect 413020 269822 413048 270535
rect 413008 269816 413060 269822
rect 413008 269758 413060 269764
rect 411352 269612 411404 269618
rect 411352 269554 411404 269560
rect 414032 268870 414060 270535
rect 415412 268938 415440 270535
rect 415400 268932 415452 268938
rect 415400 268874 415452 268880
rect 414020 268864 414072 268870
rect 414020 268806 414072 268812
rect 418172 268734 418200 270535
rect 418540 269006 418568 270535
rect 419552 269958 419580 270535
rect 419540 269952 419592 269958
rect 419540 269894 419592 269900
rect 420932 269074 420960 270535
rect 421564 270506 421616 270512
rect 420920 269068 420972 269074
rect 420920 269010 420972 269016
rect 418528 269000 418580 269006
rect 418528 268942 418580 268948
rect 418160 268728 418212 268734
rect 418160 268670 418212 268676
rect 409880 268456 409932 268462
rect 409880 268398 409932 268404
rect 396724 252068 396776 252074
rect 396724 252010 396776 252016
rect 421576 251938 421604 270506
rect 421564 251932 421616 251938
rect 421564 251874 421616 251880
rect 422956 251870 422984 270574
rect 425716 252006 425744 270846
rect 431958 270736 432014 270745
rect 431958 270671 432014 270680
rect 431972 268394 432000 270671
rect 437492 270638 437520 270943
rect 437480 270632 437532 270638
rect 436098 270600 436154 270609
rect 437480 270574 437532 270580
rect 436098 270535 436100 270544
rect 436152 270535 436154 270544
rect 436100 270506 436152 270512
rect 431960 268388 432012 268394
rect 431960 268330 432012 268336
rect 500868 253360 500920 253366
rect 500866 253328 500868 253337
rect 500920 253328 500922 253337
rect 499212 253292 499264 253298
rect 500866 253263 500922 253272
rect 499212 253234 499264 253240
rect 499224 252793 499252 253234
rect 499210 252784 499266 252793
rect 499210 252719 499266 252728
rect 510894 252648 510950 252657
rect 510894 252583 510896 252592
rect 510948 252583 510950 252592
rect 510896 252554 510948 252560
rect 425704 252000 425756 252006
rect 425704 251942 425756 251948
rect 422944 251864 422996 251870
rect 389178 251832 389234 251841
rect 422944 251806 422996 251812
rect 389178 251767 389234 251776
rect 423404 167000 423456 167006
rect 423404 166942 423456 166948
rect 416044 166932 416096 166938
rect 416044 166874 416096 166880
rect 416056 166841 416084 166874
rect 418436 166864 418488 166870
rect 416042 166832 416098 166841
rect 416042 166767 416098 166776
rect 418434 166832 418436 166841
rect 423416 166841 423444 166942
rect 418488 166832 418490 166841
rect 418434 166767 418490 166776
rect 423402 166832 423458 166841
rect 423402 166767 423458 166776
rect 425978 166832 426034 166841
rect 425978 166767 425980 166776
rect 426032 166767 426034 166776
rect 470966 166832 471022 166841
rect 470966 166767 471022 166776
rect 473450 166832 473506 166841
rect 473450 166767 473506 166776
rect 475842 166832 475898 166841
rect 475842 166767 475898 166776
rect 478418 166832 478474 166841
rect 478418 166767 478474 166776
rect 480902 166832 480958 166841
rect 480902 166767 480958 166776
rect 425980 166738 426032 166744
rect 413558 166560 413614 166569
rect 413558 166495 413614 166504
rect 408130 166288 408186 166297
rect 408130 166223 408186 166232
rect 408144 166190 408172 166223
rect 408132 166184 408184 166190
rect 408132 166126 408184 166132
rect 380900 166116 380952 166122
rect 380900 166058 380952 166064
rect 380912 146305 380940 166058
rect 397458 165608 397514 165617
rect 397458 165543 397514 165552
rect 401598 165608 401654 165617
rect 401598 165543 401654 165552
rect 404358 165608 404414 165617
rect 404358 165543 404414 165552
rect 410430 165608 410486 165617
rect 410430 165543 410486 165552
rect 396170 164384 396226 164393
rect 396170 164319 396226 164328
rect 396078 164248 396134 164257
rect 396078 164183 396134 164192
rect 396092 163810 396120 164183
rect 396080 163804 396132 163810
rect 396080 163746 396132 163752
rect 395344 161560 395396 161566
rect 395344 161502 395396 161508
rect 380898 146296 380954 146305
rect 380898 146231 380954 146240
rect 395356 146169 395384 161502
rect 395342 146160 395398 146169
rect 379980 146124 380032 146130
rect 395342 146095 395398 146104
rect 379980 146066 380032 146072
rect 379796 56296 379848 56302
rect 379796 56238 379848 56244
rect 379992 56166 380020 146066
rect 396092 145382 396120 163746
rect 396184 163742 396212 164319
rect 396172 163736 396224 163742
rect 396172 163678 396224 163684
rect 396184 145450 396212 163678
rect 396724 161492 396776 161498
rect 396724 161434 396776 161440
rect 396736 146198 396764 161434
rect 396724 146192 396776 146198
rect 396724 146134 396776 146140
rect 397472 145518 397500 165543
rect 398838 164248 398894 164257
rect 398838 164183 398894 164192
rect 400218 164248 400274 164257
rect 400218 164183 400274 164192
rect 398852 148510 398880 164183
rect 398840 148504 398892 148510
rect 398840 148446 398892 148452
rect 400232 148442 400260 164183
rect 401612 148986 401640 165543
rect 402978 164384 403034 164393
rect 402978 164319 403034 164328
rect 401600 148980 401652 148986
rect 401600 148922 401652 148928
rect 400220 148436 400272 148442
rect 400220 148378 400272 148384
rect 402992 145790 403020 164319
rect 403070 164248 403126 164257
rect 403070 164183 403126 164192
rect 402980 145784 403032 145790
rect 402980 145726 403032 145732
rect 403084 145722 403112 164183
rect 403072 145716 403124 145722
rect 403072 145658 403124 145664
rect 404372 145586 404400 165543
rect 410444 164694 410472 165543
rect 413572 164762 413600 166495
rect 470980 166462 471008 166767
rect 473464 166734 473492 166767
rect 473452 166728 473504 166734
rect 473452 166670 473504 166676
rect 475856 166666 475884 166767
rect 475844 166660 475896 166666
rect 475844 166602 475896 166608
rect 478432 166598 478460 166767
rect 478420 166592 478472 166598
rect 478420 166534 478472 166540
rect 480916 166530 480944 166767
rect 483386 166696 483442 166705
rect 483386 166631 483442 166640
rect 485962 166696 486018 166705
rect 485962 166631 486018 166640
rect 480904 166524 480956 166530
rect 480904 166466 480956 166472
rect 470968 166456 471020 166462
rect 470968 166398 471020 166404
rect 483400 166326 483428 166631
rect 485976 166394 486004 166631
rect 503258 166560 503314 166569
rect 503258 166495 503314 166504
rect 485964 166388 486016 166394
rect 485964 166330 486016 166336
rect 483388 166320 483440 166326
rect 428186 166288 428242 166297
rect 483388 166262 483440 166268
rect 428186 166223 428188 166232
rect 428240 166223 428242 166232
rect 428188 166194 428240 166200
rect 415398 165608 415454 165617
rect 415398 165543 415454 165552
rect 416870 165608 416926 165617
rect 416870 165543 416926 165552
rect 418158 165608 418214 165617
rect 418158 165543 418214 165552
rect 423770 165608 423826 165617
rect 423770 165543 423826 165552
rect 426438 165608 426494 165617
rect 426438 165543 426494 165552
rect 434626 165608 434682 165617
rect 434810 165608 434866 165617
rect 434682 165566 434760 165594
rect 434626 165543 434682 165552
rect 413560 164756 413612 164762
rect 413560 164698 413612 164704
rect 410432 164688 410484 164694
rect 410432 164630 410484 164636
rect 411350 164384 411406 164393
rect 411350 164319 411406 164328
rect 405738 164248 405794 164257
rect 405738 164183 405794 164192
rect 407118 164248 407174 164257
rect 407118 164183 407174 164192
rect 408498 164248 408554 164257
rect 408498 164183 408554 164192
rect 409970 164248 410026 164257
rect 409970 164183 410026 164192
rect 411258 164248 411314 164257
rect 411258 164183 411314 164192
rect 405752 145654 405780 164183
rect 407132 145994 407160 164183
rect 407120 145988 407172 145994
rect 407120 145930 407172 145936
rect 408512 145858 408540 164183
rect 409984 145926 410012 164183
rect 411272 146062 411300 164183
rect 411260 146056 411312 146062
rect 411260 145998 411312 146004
rect 409972 145920 410024 145926
rect 409972 145862 410024 145868
rect 408500 145852 408552 145858
rect 408500 145794 408552 145800
rect 405740 145648 405792 145654
rect 405740 145590 405792 145596
rect 404360 145580 404412 145586
rect 404360 145522 404412 145528
rect 397460 145512 397512 145518
rect 397460 145454 397512 145460
rect 396172 145444 396224 145450
rect 396172 145386 396224 145392
rect 396080 145376 396132 145382
rect 396080 145318 396132 145324
rect 411364 145314 411392 164319
rect 412730 164248 412786 164257
rect 412730 164183 412786 164192
rect 414018 164248 414074 164257
rect 414018 164183 414074 164192
rect 412744 149054 412772 164183
rect 412732 149048 412784 149054
rect 412732 148990 412784 148996
rect 414032 146130 414060 164183
rect 415412 146169 415440 165543
rect 416884 163878 416912 165543
rect 416872 163872 416924 163878
rect 416872 163814 416924 163820
rect 418172 146198 418200 165543
rect 422944 165096 422996 165102
rect 422944 165038 422996 165044
rect 420918 164928 420974 164937
rect 420918 164863 420974 164872
rect 420932 164830 420960 164863
rect 422956 164830 422984 165038
rect 420920 164824 420972 164830
rect 420920 164766 420972 164772
rect 422944 164824 422996 164830
rect 422944 164766 422996 164772
rect 418250 164248 418306 164257
rect 418250 164183 418306 164192
rect 419538 164248 419594 164257
rect 419538 164183 419594 164192
rect 420918 164248 420974 164257
rect 420918 164183 420974 164192
rect 423586 164248 423642 164257
rect 423642 164206 423720 164234
rect 423586 164183 423642 164192
rect 418264 162246 418292 164183
rect 419552 162654 419580 164183
rect 420932 162722 420960 164183
rect 420920 162716 420972 162722
rect 420920 162658 420972 162664
rect 419540 162648 419592 162654
rect 419540 162590 419592 162596
rect 418252 162240 418304 162246
rect 418252 162182 418304 162188
rect 418160 146192 418212 146198
rect 415398 146160 415454 146169
rect 414020 146124 414072 146130
rect 418160 146134 418212 146140
rect 415398 146095 415454 146104
rect 414020 146066 414072 146072
rect 423692 145761 423720 164206
rect 423784 145897 423812 165543
rect 425058 164248 425114 164257
rect 425058 164183 425114 164192
rect 425072 163946 425100 164183
rect 426452 164014 426480 165543
rect 433338 164928 433394 164937
rect 433338 164863 433394 164872
rect 433352 164830 433380 164863
rect 433340 164824 433392 164830
rect 433340 164766 433392 164772
rect 433338 164656 433394 164665
rect 433338 164591 433394 164600
rect 433352 164558 433380 164591
rect 428832 164552 428884 164558
rect 428832 164494 428884 164500
rect 433340 164552 433392 164558
rect 433340 164494 433392 164500
rect 427726 164248 427782 164257
rect 427782 164206 427860 164234
rect 427726 164183 427782 164192
rect 426440 164008 426492 164014
rect 426440 163950 426492 163956
rect 425060 163940 425112 163946
rect 425060 163882 425112 163888
rect 423770 145888 423826 145897
rect 423770 145823 423826 145832
rect 423678 145752 423734 145761
rect 423678 145687 423734 145696
rect 427832 145625 427860 164206
rect 428844 162790 428872 164494
rect 429290 164384 429346 164393
rect 429290 164319 429346 164328
rect 430670 164384 430726 164393
rect 430670 164319 430726 164328
rect 429106 164248 429162 164257
rect 429162 164206 429240 164234
rect 429106 164183 429162 164192
rect 428832 162784 428884 162790
rect 428832 162726 428884 162732
rect 429212 146305 429240 164206
rect 429304 164082 429332 164319
rect 430578 164248 430634 164257
rect 430578 164183 430634 164192
rect 430592 164150 430620 164183
rect 430580 164144 430632 164150
rect 430580 164086 430632 164092
rect 429292 164076 429344 164082
rect 429292 164018 429344 164024
rect 430684 163606 430712 164319
rect 431958 164248 432014 164257
rect 431958 164183 432014 164192
rect 430672 163600 430724 163606
rect 430672 163542 430724 163548
rect 431972 162178 432000 164183
rect 431960 162172 432012 162178
rect 431960 162114 432012 162120
rect 434732 148374 434760 165566
rect 434810 165543 434866 165552
rect 437846 165608 437902 165617
rect 437846 165543 437902 165552
rect 440238 165608 440294 165617
rect 440238 165543 440294 165552
rect 442998 165608 443054 165617
rect 442998 165543 443054 165552
rect 447322 165608 447378 165617
rect 447322 165543 447378 165552
rect 449898 165608 449954 165617
rect 449898 165543 449954 165552
rect 452658 165608 452714 165617
rect 452658 165543 452660 165552
rect 434824 164966 434852 165543
rect 437754 165064 437810 165073
rect 437754 164999 437810 165008
rect 434812 164960 434864 164966
rect 434812 164902 434864 164908
rect 437768 164898 437796 164999
rect 437756 164892 437808 164898
rect 437756 164834 437808 164840
rect 434810 164248 434866 164257
rect 434810 164183 434866 164192
rect 436098 164248 436154 164257
rect 437860 164218 437888 165543
rect 440252 165170 440280 165543
rect 443012 165442 443040 165543
rect 443000 165436 443052 165442
rect 443000 165378 443052 165384
rect 447336 165238 447364 165543
rect 449912 165374 449940 165543
rect 452712 165543 452714 165552
rect 455418 165608 455474 165617
rect 455418 165543 455474 165552
rect 458362 165608 458418 165617
rect 458362 165543 458418 165552
rect 452660 165514 452712 165520
rect 455432 165510 455460 165543
rect 455420 165504 455472 165510
rect 455420 165446 455472 165452
rect 449900 165368 449952 165374
rect 449900 165310 449952 165316
rect 458376 165306 458404 165543
rect 458364 165300 458416 165306
rect 458364 165242 458416 165248
rect 447324 165232 447376 165238
rect 447324 165174 447376 165180
rect 440240 165164 440292 165170
rect 440240 165106 440292 165112
rect 445758 165064 445814 165073
rect 503272 165034 503300 166495
rect 503628 165164 503680 165170
rect 503628 165106 503680 165112
rect 445758 164999 445760 165008
rect 445812 164999 445814 165008
rect 503260 165028 503312 165034
rect 445760 164970 445812 164976
rect 503260 164970 503312 164976
rect 440240 164960 440292 164966
rect 440240 164902 440292 164908
rect 440146 164248 440202 164257
rect 436098 164183 436154 164192
rect 437848 164212 437900 164218
rect 434824 162858 434852 164183
rect 436112 163538 436140 164183
rect 440252 164234 440280 164902
rect 503640 164665 503668 165106
rect 516612 165034 516640 271866
rect 517532 252618 517560 358770
rect 517624 271182 517652 378218
rect 517704 378208 517756 378214
rect 517704 378150 517756 378156
rect 517716 271318 517744 378150
rect 517808 364334 517836 466414
rect 517900 383654 517928 466550
rect 517900 383626 518112 383654
rect 517808 364306 518020 364334
rect 517992 359650 518020 364306
rect 518084 359718 518112 383626
rect 518072 359712 518124 359718
rect 518072 359654 518124 359660
rect 517980 359644 518032 359650
rect 517980 359586 518032 359592
rect 517704 271312 517756 271318
rect 517704 271254 517756 271260
rect 517612 271176 517664 271182
rect 517612 271118 517664 271124
rect 517624 270842 517652 271118
rect 517612 270836 517664 270842
rect 517612 270778 517664 270784
rect 517716 267734 517744 271254
rect 517888 270836 517940 270842
rect 517888 270778 517940 270784
rect 517716 267706 517836 267734
rect 517704 253360 517756 253366
rect 517704 253302 517756 253308
rect 517612 253292 517664 253298
rect 517612 253234 517664 253240
rect 517520 252612 517572 252618
rect 517520 252554 517572 252560
rect 516600 165028 516652 165034
rect 516600 164970 516652 164976
rect 517532 164966 517560 252554
rect 510528 164960 510580 164966
rect 510528 164902 510580 164908
rect 517520 164960 517572 164966
rect 517520 164902 517572 164908
rect 503626 164656 503682 164665
rect 503626 164591 503682 164600
rect 440202 164206 440280 164234
rect 440146 164183 440202 164192
rect 437848 164154 437900 164160
rect 436100 163532 436152 163538
rect 436100 163474 436152 163480
rect 434812 162852 434864 162858
rect 434812 162794 434864 162800
rect 434720 148368 434772 148374
rect 434720 148310 434772 148316
rect 429198 146296 429254 146305
rect 429198 146231 429254 146240
rect 427818 145616 427874 145625
rect 427818 145551 427874 145560
rect 411352 145308 411404 145314
rect 411352 145250 411404 145256
rect 440252 144129 440280 164206
rect 498660 146192 498712 146198
rect 498660 146134 498712 146140
rect 498672 144945 498700 146134
rect 499856 146124 499908 146130
rect 499856 146066 499908 146072
rect 499868 144945 499896 146066
rect 503640 145722 503668 164591
rect 510540 146282 510568 164902
rect 510540 146266 510660 146282
rect 510540 146260 510672 146266
rect 510540 146254 510620 146260
rect 510620 146202 510672 146208
rect 510632 146169 510660 146202
rect 517624 146198 517652 253234
rect 517716 253230 517744 253302
rect 517704 253224 517756 253230
rect 517704 253166 517756 253172
rect 517612 146192 517664 146198
rect 510618 146160 510674 146169
rect 517612 146134 517664 146140
rect 517716 146130 517744 253166
rect 517808 165170 517836 267706
rect 517796 165164 517848 165170
rect 517796 165106 517848 165112
rect 517900 165102 517928 270778
rect 517992 253298 518020 359586
rect 517980 253292 518032 253298
rect 517980 253234 518032 253240
rect 518084 253230 518112 359654
rect 518176 353258 518204 499530
rect 518900 465112 518952 465118
rect 518900 465054 518952 465060
rect 518912 459649 518940 465054
rect 518898 459640 518954 459649
rect 518898 459575 518954 459584
rect 519450 459640 519506 459649
rect 519450 459575 519506 459584
rect 519358 400344 519414 400353
rect 519358 400279 519414 400288
rect 518990 398168 519046 398177
rect 518990 398103 519046 398112
rect 519004 365022 519032 398103
rect 519174 396808 519230 396817
rect 519174 396743 519230 396752
rect 519082 395312 519138 395321
rect 519082 395247 519138 395256
rect 519096 376038 519124 395247
rect 519084 376032 519136 376038
rect 519084 375974 519136 375980
rect 518992 365016 519044 365022
rect 518992 364958 519044 364964
rect 519004 354674 519032 364958
rect 518912 354646 519032 354674
rect 518164 353252 518216 353258
rect 518164 353194 518216 353200
rect 518912 291689 518940 354646
rect 518898 291680 518954 291689
rect 518954 291638 519032 291666
rect 518898 291615 518954 291624
rect 518072 253224 518124 253230
rect 518072 253166 518124 253172
rect 518898 186416 518954 186425
rect 518898 186351 518954 186360
rect 517888 165096 517940 165102
rect 517888 165038 517940 165044
rect 510618 146095 510674 146104
rect 517520 146124 517572 146130
rect 517520 146066 517572 146072
rect 517704 146124 517756 146130
rect 517704 146066 517756 146072
rect 503628 145716 503680 145722
rect 503628 145658 503680 145664
rect 517532 145654 517560 146066
rect 517796 145716 517848 145722
rect 517796 145658 517848 145664
rect 517520 145648 517572 145654
rect 517520 145590 517572 145596
rect 498658 144936 498714 144945
rect 498658 144871 498714 144880
rect 499854 144936 499910 144945
rect 499854 144871 499910 144880
rect 440238 144120 440294 144129
rect 440238 144055 440294 144064
rect 396078 59800 396134 59809
rect 396078 59735 396080 59744
rect 396132 59735 396134 59744
rect 397090 59800 397146 59809
rect 397090 59735 397146 59744
rect 403070 59800 403126 59809
rect 403070 59735 403126 59744
rect 413558 59800 413614 59809
rect 413558 59735 413614 59744
rect 415858 59800 415914 59809
rect 415858 59735 415914 59744
rect 419446 59800 419502 59809
rect 419446 59735 419502 59744
rect 396080 59706 396132 59712
rect 397104 59702 397132 59735
rect 397092 59696 397144 59702
rect 397092 59638 397144 59644
rect 403084 59634 403112 59735
rect 403072 59628 403124 59634
rect 403072 59570 403124 59576
rect 413572 59430 413600 59735
rect 415872 59566 415900 59735
rect 415860 59560 415912 59566
rect 415860 59502 415912 59508
rect 419460 59498 419488 59735
rect 423494 59664 423550 59673
rect 423494 59599 423550 59608
rect 503258 59664 503314 59673
rect 503258 59599 503314 59608
rect 419448 59492 419500 59498
rect 419448 59434 419500 59440
rect 413560 59424 413612 59430
rect 398194 59392 398250 59401
rect 398194 59327 398196 59336
rect 398248 59327 398250 59336
rect 410706 59392 410762 59401
rect 413560 59366 413612 59372
rect 416962 59392 417018 59401
rect 410706 59327 410762 59336
rect 416962 59327 417018 59336
rect 418158 59392 418214 59401
rect 418158 59327 418214 59336
rect 421010 59392 421066 59401
rect 421010 59327 421066 59336
rect 421746 59392 421802 59401
rect 421746 59327 421802 59336
rect 398196 59298 398248 59304
rect 410720 59294 410748 59327
rect 410708 59288 410760 59294
rect 410708 59230 410760 59236
rect 416976 59226 417004 59327
rect 416964 59220 417016 59226
rect 416964 59162 417016 59168
rect 418172 59158 418200 59327
rect 418160 59152 418212 59158
rect 418160 59094 418212 59100
rect 421024 58750 421052 59327
rect 421760 59022 421788 59327
rect 421748 59016 421800 59022
rect 421748 58958 421800 58964
rect 423508 58954 423536 59599
rect 425242 59392 425298 59401
rect 425242 59327 425298 59336
rect 425978 59392 426034 59401
rect 425978 59327 426034 59336
rect 428186 59392 428242 59401
rect 428186 59327 428242 59336
rect 468482 59392 468538 59401
rect 468482 59327 468538 59336
rect 425256 59090 425284 59327
rect 425244 59084 425296 59090
rect 425244 59026 425296 59032
rect 423496 58948 423548 58954
rect 423496 58890 423548 58896
rect 425992 58818 426020 59327
rect 425980 58812 426032 58818
rect 425980 58754 426032 58760
rect 421012 58744 421064 58750
rect 421012 58686 421064 58692
rect 428200 58682 428228 59327
rect 468496 58886 468524 59327
rect 468484 58880 468536 58886
rect 468484 58822 468536 58828
rect 428188 58676 428240 58682
rect 428188 58618 428240 58624
rect 430948 57996 431000 58002
rect 430948 57938 431000 57944
rect 430960 57905 430988 57938
rect 475844 57928 475896 57934
rect 398838 57896 398894 57905
rect 398838 57831 398894 57840
rect 400402 57896 400458 57905
rect 400402 57831 400458 57840
rect 401598 57896 401654 57905
rect 401598 57831 401654 57840
rect 404082 57896 404138 57905
rect 404082 57831 404138 57840
rect 404358 57896 404414 57905
rect 404358 57831 404414 57840
rect 405830 57896 405886 57905
rect 405830 57831 405886 57840
rect 407118 57896 407174 57905
rect 407118 57831 407174 57840
rect 408314 57896 408370 57905
rect 408314 57831 408370 57840
rect 408682 57896 408738 57905
rect 408682 57831 408738 57840
rect 409878 57896 409934 57905
rect 409878 57831 409934 57840
rect 411350 57896 411406 57905
rect 411350 57831 411406 57840
rect 413466 57896 413522 57905
rect 413466 57831 413522 57840
rect 414570 57896 414626 57905
rect 414570 57831 414626 57840
rect 418434 57896 418490 57905
rect 418434 57831 418490 57840
rect 422850 57896 422906 57905
rect 422850 57831 422906 57840
rect 423678 57896 423734 57905
rect 423678 57831 423734 57840
rect 426530 57896 426586 57905
rect 426530 57831 426586 57840
rect 427634 57896 427690 57905
rect 427634 57831 427690 57840
rect 427818 57896 427874 57905
rect 427818 57831 427874 57840
rect 429658 57896 429714 57905
rect 429658 57831 429714 57840
rect 430946 57896 431002 57905
rect 430946 57831 431002 57840
rect 431958 57896 432014 57905
rect 431958 57831 432014 57840
rect 433338 57896 433394 57905
rect 433338 57831 433394 57840
rect 433522 57896 433578 57905
rect 433522 57831 433578 57840
rect 435086 57896 435142 57905
rect 435086 57831 435142 57840
rect 435914 57896 435970 57905
rect 435914 57831 435970 57840
rect 438490 57896 438546 57905
rect 438490 57831 438546 57840
rect 460938 57896 460994 57905
rect 460938 57831 460994 57840
rect 465906 57896 465962 57905
rect 465906 57831 465962 57840
rect 470874 57896 470930 57905
rect 470874 57831 470930 57840
rect 475842 57896 475844 57905
rect 475896 57896 475898 57905
rect 475842 57831 475898 57840
rect 480626 57896 480682 57905
rect 480626 57831 480628 57840
rect 379980 56160 380032 56166
rect 379980 56102 380032 56108
rect 379336 56092 379388 56098
rect 379336 56034 379388 56040
rect 379244 55956 379296 55962
rect 379244 55898 379296 55904
rect 379060 55004 379112 55010
rect 379060 54946 379112 54952
rect 378784 54596 378836 54602
rect 378784 54538 378836 54544
rect 374920 54528 374972 54534
rect 374920 54470 374972 54476
rect 398852 54466 398880 57831
rect 400416 55826 400444 57831
rect 400404 55820 400456 55826
rect 400404 55762 400456 55768
rect 401612 54534 401640 57831
rect 404096 55894 404124 57831
rect 404084 55888 404136 55894
rect 404084 55830 404136 55836
rect 404372 54670 404400 57831
rect 404360 54664 404412 54670
rect 404360 54606 404412 54612
rect 405844 54602 405872 57831
rect 407132 54738 407160 57831
rect 408328 57254 408356 57831
rect 408316 57248 408368 57254
rect 408316 57190 408368 57196
rect 408696 56030 408724 57831
rect 408684 56024 408736 56030
rect 408684 55966 408736 55972
rect 409892 54806 409920 57831
rect 411258 56944 411314 56953
rect 411258 56879 411314 56888
rect 411272 55962 411300 56879
rect 411260 55956 411312 55962
rect 411260 55898 411312 55904
rect 411364 54874 411392 57831
rect 413480 56098 413508 57831
rect 414584 56166 414612 57831
rect 418448 57322 418476 57831
rect 418436 57316 418488 57322
rect 418436 57258 418488 57264
rect 422864 56234 422892 57831
rect 422852 56228 422904 56234
rect 422852 56170 422904 56176
rect 414572 56160 414624 56166
rect 414572 56102 414624 56108
rect 413468 56092 413520 56098
rect 413468 56034 413520 56040
rect 423692 54942 423720 57831
rect 426544 55010 426572 57831
rect 427648 56302 427676 57831
rect 427636 56296 427688 56302
rect 427636 56238 427688 56244
rect 427832 55049 427860 57831
rect 429672 56370 429700 57831
rect 430578 57080 430634 57089
rect 430578 57015 430634 57024
rect 430592 56438 430620 57015
rect 430580 56432 430632 56438
rect 430580 56374 430632 56380
rect 429660 56364 429712 56370
rect 429660 56306 429712 56312
rect 431972 55078 432000 57831
rect 433352 56506 433380 57831
rect 433536 57526 433564 57831
rect 433524 57520 433576 57526
rect 433430 57488 433486 57497
rect 433524 57462 433576 57468
rect 433706 57488 433762 57497
rect 433430 57423 433486 57432
rect 433706 57423 433762 57432
rect 433444 57089 433472 57423
rect 433430 57080 433486 57089
rect 433430 57015 433486 57024
rect 433340 56500 433392 56506
rect 433340 56442 433392 56448
rect 433720 55146 433748 57423
rect 435100 56574 435128 57831
rect 435928 57390 435956 57831
rect 436098 57488 436154 57497
rect 438504 57458 438532 57831
rect 460952 57662 460980 57831
rect 465920 57730 465948 57831
rect 465908 57724 465960 57730
rect 465908 57666 465960 57672
rect 460940 57656 460992 57662
rect 460940 57598 460992 57604
rect 470888 57594 470916 57831
rect 480680 57831 480682 57840
rect 483386 57896 483442 57905
rect 503272 57866 503300 59599
rect 517808 57934 517836 145658
rect 503352 57928 503404 57934
rect 503350 57896 503352 57905
rect 517796 57928 517848 57934
rect 503404 57896 503406 57905
rect 483386 57831 483442 57840
rect 503260 57860 503312 57866
rect 480628 57802 480680 57808
rect 483400 57798 483428 57831
rect 517796 57870 517848 57876
rect 517900 57866 517928 165038
rect 518440 146192 518492 146198
rect 518440 146134 518492 146140
rect 518452 145586 518480 146134
rect 518440 145580 518492 145586
rect 518440 145522 518492 145528
rect 518912 93854 518940 186351
rect 519004 184793 519032 291638
rect 519096 288833 519124 375974
rect 519188 370530 519216 396743
rect 519266 394088 519322 394097
rect 519266 394023 519322 394032
rect 519280 373318 519308 394023
rect 519268 373312 519320 373318
rect 519268 373254 519320 373260
rect 519280 372638 519308 373254
rect 519268 372632 519320 372638
rect 519268 372574 519320 372580
rect 519176 370524 519228 370530
rect 519176 370466 519228 370472
rect 519372 369238 519400 400279
rect 519360 369232 519412 369238
rect 519360 369174 519412 369180
rect 519266 352880 519322 352889
rect 519266 352815 519322 352824
rect 519082 288824 519138 288833
rect 519082 288759 519138 288768
rect 518990 184784 519046 184793
rect 518990 184719 519046 184728
rect 519096 181937 519124 288759
rect 519174 287600 519230 287609
rect 519174 287535 519230 287544
rect 519188 287094 519216 287535
rect 519176 287088 519228 287094
rect 519176 287030 519228 287036
rect 519082 181928 519138 181937
rect 519082 181863 519138 181872
rect 518912 93826 519032 93854
rect 519004 79937 519032 93826
rect 518990 79928 519046 79937
rect 518990 79863 519046 79872
rect 519096 75449 519124 181863
rect 519188 180713 519216 287030
rect 519280 246265 519308 352815
rect 519372 293865 519400 369174
rect 519464 352889 519492 459575
rect 520936 405686 520964 529926
rect 578896 511329 578924 592010
rect 580276 577697 580304 640290
rect 580368 630873 580396 645118
rect 580354 630864 580410 630873
rect 580354 630799 580410 630808
rect 580262 577688 580318 577697
rect 580262 577623 580318 577632
rect 578882 511320 578938 511329
rect 578882 511255 578938 511264
rect 580264 494760 580316 494766
rect 580264 494702 580316 494708
rect 580276 458153 580304 494702
rect 580262 458144 580318 458153
rect 580262 458079 580318 458088
rect 520924 405680 520976 405686
rect 520924 405622 520976 405628
rect 580172 405680 580224 405686
rect 580172 405622 580224 405628
rect 580184 404977 580212 405622
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580264 378276 580316 378282
rect 580264 378218 580316 378224
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 519636 372632 519688 372638
rect 519636 372574 519688 372580
rect 519544 370524 519596 370530
rect 519544 370466 519596 370472
rect 519450 352880 519506 352889
rect 519450 352815 519506 352824
rect 519358 293856 519414 293865
rect 519358 293791 519414 293800
rect 519266 246256 519322 246265
rect 519266 246191 519322 246200
rect 519174 180704 519230 180713
rect 519174 180639 519230 180648
rect 519082 75440 519138 75449
rect 519082 75375 519138 75384
rect 519188 74225 519216 180639
rect 519280 139369 519308 246191
rect 519372 186425 519400 293791
rect 519556 290329 519584 370466
rect 519542 290320 519598 290329
rect 519542 290255 519598 290264
rect 519556 277394 519584 290255
rect 519648 287094 519676 372574
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 580276 325281 580304 378218
rect 580262 325272 580318 325281
rect 580262 325207 580318 325216
rect 520186 288824 520242 288833
rect 520186 288759 520242 288768
rect 520200 288454 520228 288759
rect 520188 288448 520240 288454
rect 520188 288390 520240 288396
rect 580264 288448 580316 288454
rect 580264 288390 580316 288396
rect 519636 287088 519688 287094
rect 519636 287030 519688 287036
rect 519464 277366 519584 277394
rect 519358 186416 519414 186425
rect 519358 186351 519414 186360
rect 519360 183592 519412 183598
rect 519360 183534 519412 183540
rect 519266 139360 519322 139369
rect 519266 139295 519322 139304
rect 519372 78305 519400 183534
rect 519464 183433 519492 277366
rect 580276 232393 580304 288390
rect 580356 287088 580408 287094
rect 580356 287030 580408 287036
rect 580368 272241 580396 287030
rect 580354 272232 580410 272241
rect 580354 272167 580410 272176
rect 580262 232384 580318 232393
rect 580262 232319 580318 232328
rect 580354 192536 580410 192545
rect 580354 192471 580410 192480
rect 520186 184784 520242 184793
rect 520186 184719 520242 184728
rect 520200 183598 520228 184719
rect 520188 183592 520240 183598
rect 520188 183534 520240 183540
rect 580264 183592 580316 183598
rect 580264 183534 580316 183540
rect 520096 183524 520148 183530
rect 520096 183466 520148 183472
rect 520108 183433 520136 183466
rect 519450 183424 519506 183433
rect 519450 183359 519506 183368
rect 520094 183424 520150 183433
rect 520094 183359 520150 183368
rect 519358 78296 519414 78305
rect 519358 78231 519414 78240
rect 519464 76809 519492 183359
rect 580276 152697 580304 183534
rect 580368 183530 580396 192471
rect 580356 183524 580408 183530
rect 580356 183466 580408 183472
rect 580262 152688 580318 152697
rect 580262 152623 580318 152632
rect 580264 145648 580316 145654
rect 580264 145590 580316 145596
rect 520188 80028 520240 80034
rect 520188 79970 520240 79976
rect 520200 79937 520228 79970
rect 520186 79928 520242 79937
rect 520186 79863 520242 79872
rect 519450 76800 519506 76809
rect 519450 76735 519506 76744
rect 519174 74216 519230 74225
rect 519174 74151 519230 74160
rect 503350 57831 503406 57840
rect 517888 57860 517940 57866
rect 503260 57802 503312 57808
rect 517888 57802 517940 57808
rect 483388 57792 483440 57798
rect 483388 57734 483440 57740
rect 470876 57588 470928 57594
rect 470876 57530 470928 57536
rect 438858 57488 438914 57497
rect 436098 57423 436154 57432
rect 438492 57452 438544 57458
rect 435916 57384 435968 57390
rect 435916 57326 435968 57332
rect 435088 56568 435140 56574
rect 435088 56510 435140 56516
rect 436112 55214 436140 57423
rect 438858 57423 438914 57432
rect 438492 57394 438544 57400
rect 436100 55208 436152 55214
rect 438872 55185 438900 57423
rect 436100 55150 436152 55156
rect 438858 55176 438914 55185
rect 433708 55140 433760 55146
rect 438858 55111 438914 55120
rect 433708 55082 433760 55088
rect 431960 55072 432012 55078
rect 427818 55040 427874 55049
rect 426532 55004 426584 55010
rect 431960 55014 432012 55020
rect 427818 54975 427874 54984
rect 426532 54946 426584 54952
rect 423680 54936 423732 54942
rect 423680 54878 423732 54884
rect 411352 54868 411404 54874
rect 411352 54810 411404 54816
rect 409880 54800 409932 54806
rect 409880 54742 409932 54748
rect 407120 54732 407172 54738
rect 407120 54674 407172 54680
rect 405832 54596 405884 54602
rect 405832 54538 405884 54544
rect 401600 54528 401652 54534
rect 401600 54470 401652 54476
rect 374828 54460 374880 54466
rect 374828 54402 374880 54408
rect 398840 54460 398892 54466
rect 398840 54402 398892 54408
rect 580276 33153 580304 145590
rect 580356 145580 580408 145586
rect 580356 145522 580408 145528
rect 580368 73001 580396 145522
rect 580446 112840 580502 112849
rect 580446 112775 580502 112784
rect 580460 80034 580488 112775
rect 580448 80028 580500 80034
rect 580448 79970 580500 79976
rect 580354 72992 580410 73001
rect 580354 72927 580410 72936
rect 580262 33144 580318 33153
rect 580262 33079 580318 33088
rect 366364 3460 366416 3466
rect 366364 3402 366416 3408
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3422 632032 3478 632088
rect 3146 579944 3202 580000
rect 2962 410488 3018 410544
rect 3330 358400 3386 358456
rect 3514 514800 3570 514856
rect 3422 97552 3478 97608
rect 3606 462576 3662 462632
rect 3514 58520 3570 58576
rect 57702 640600 57758 640656
rect 57610 631760 57666 631816
rect 57518 613400 57574 613456
rect 57426 607280 57482 607336
rect 57334 601160 57390 601216
rect 57242 591640 57298 591696
rect 57150 585520 57206 585576
rect 57058 582800 57114 582856
rect 57794 634480 57850 634536
rect 59082 637880 59138 637936
rect 58898 628360 58954 628416
rect 58530 625640 58586 625696
rect 57886 616120 57942 616176
rect 58438 597760 58494 597816
rect 58806 610000 58862 610056
rect 58622 603880 58678 603936
rect 58714 588920 58770 588976
rect 58990 622240 59046 622296
rect 59174 619520 59230 619576
rect 59174 595040 59230 595096
rect 120814 618296 120870 618352
rect 120722 581576 120778 581632
rect 121090 603200 121146 603256
rect 121550 633800 121606 633856
rect 121826 631080 121882 631136
rect 121734 627680 121790 627736
rect 121918 621560 121974 621616
rect 122010 606600 122066 606656
rect 122102 600480 122158 600536
rect 122194 597080 122250 597136
rect 122286 588240 122342 588296
rect 122930 639920 122986 639976
rect 123114 637200 123170 637256
rect 123022 612720 123078 612776
rect 123206 624960 123262 625016
rect 123114 584840 123170 584896
rect 123390 615440 123446 615496
rect 123298 594360 123354 594416
rect 124034 609320 124090 609376
rect 123482 590960 123538 591016
rect 146298 640600 146354 640656
rect 146298 631760 146354 631816
rect 146298 628360 146354 628416
rect 147218 625640 147274 625696
rect 146206 616120 146262 616176
rect 146298 610020 146354 610056
rect 146298 610000 146300 610020
rect 146300 610000 146352 610020
rect 146352 610000 146354 610020
rect 147126 607280 147182 607336
rect 146298 597760 146354 597816
rect 146942 595040 146998 595096
rect 146298 591640 146354 591696
rect 147034 588920 147090 588976
rect 147402 634480 147458 634536
rect 147310 619520 147366 619576
rect 147310 601160 147366 601216
rect 148230 603880 148286 603936
rect 148598 637880 148654 637936
rect 148506 613400 148562 613456
rect 148690 622240 148746 622296
rect 149058 585520 149114 585576
rect 148966 582800 149022 582856
rect 210790 584296 210846 584352
rect 210882 581576 210938 581632
rect 211250 639376 211306 639432
rect 212630 636656 212686 636712
rect 211342 630672 211398 630728
rect 212538 627136 212594 627192
rect 211526 624416 211582 624472
rect 211434 621016 211490 621072
rect 211710 606192 211766 606248
rect 211618 600616 211674 600672
rect 211802 596672 211858 596728
rect 211894 587968 211950 588024
rect 212722 633392 212778 633448
rect 212814 618296 212870 618352
rect 212998 614896 213054 614952
rect 212906 612856 212962 612912
rect 213826 608776 213882 608832
rect 213090 603336 213146 603392
rect 213274 593816 213330 593872
rect 213182 590688 213238 590744
rect 237378 640736 237434 640792
rect 237378 634344 237434 634400
rect 237378 631624 237434 631680
rect 237378 625504 237434 625560
rect 237378 622104 237434 622160
rect 238022 616120 238078 616176
rect 237378 613264 237434 613320
rect 237378 610020 237434 610056
rect 237378 610000 237380 610020
rect 237380 610000 237432 610020
rect 237432 610000 237434 610020
rect 237378 607280 237434 607336
rect 237378 603744 237434 603800
rect 237378 601024 237434 601080
rect 237378 597624 237434 597680
rect 237378 594904 237434 594960
rect 237378 591504 237434 591560
rect 237378 588784 237434 588840
rect 237378 585384 237434 585440
rect 237378 582664 237434 582720
rect 238206 637744 238262 637800
rect 238298 628224 238354 628280
rect 238850 619520 238906 619576
rect 238666 554920 238722 554976
rect 300858 639376 300914 639432
rect 300674 581576 300730 581632
rect 241518 555056 241574 555112
rect 249430 553832 249486 553888
rect 255134 555464 255190 555520
rect 286690 555192 286746 555248
rect 285954 554784 286010 554840
rect 293130 553696 293186 553752
rect 293774 553560 293830 553616
rect 294510 553424 294566 553480
rect 300950 636656 301006 636712
rect 302238 633392 302294 633448
rect 301042 630672 301098 630728
rect 301134 624416 301190 624472
rect 301226 612856 301282 612912
rect 301318 606192 301374 606248
rect 301410 600616 301466 600672
rect 301502 593816 301558 593872
rect 301594 587968 301650 588024
rect 302330 627136 302386 627192
rect 302422 621016 302478 621072
rect 302606 618296 302662 618352
rect 302514 614896 302570 614952
rect 303158 609456 303214 609512
rect 302698 603336 302754 603392
rect 302974 596672 303030 596728
rect 302882 590688 302938 590744
rect 298098 555328 298154 555384
rect 300214 554920 300270 554976
rect 300582 555056 300638 555112
rect 300582 534520 300638 534576
rect 301962 553832 302018 553888
rect 302238 545400 302294 545456
rect 301962 532616 302018 532672
rect 302422 530440 302478 530496
rect 57702 522960 57758 523016
rect 57886 522960 57942 523016
rect 41326 485560 41382 485616
rect 43994 485016 44050 485072
rect 46110 379344 46166 379400
rect 46662 488008 46718 488064
rect 46478 487872 46534 487928
rect 46570 485152 46626 485208
rect 47490 379072 47546 379128
rect 47674 379208 47730 379264
rect 47490 271768 47546 271824
rect 48134 485288 48190 485344
rect 47858 271632 47914 271688
rect 49146 488144 49202 488200
rect 49054 271768 49110 271824
rect 49054 271224 49110 271280
rect 50894 490456 50950 490512
rect 49238 164600 49294 164656
rect 50342 272992 50398 273048
rect 50526 272856 50582 272912
rect 50710 465160 50766 465216
rect 50618 165416 50674 165472
rect 51630 272720 51686 272776
rect 52182 379480 52238 379536
rect 52458 271532 52460 271552
rect 52460 271532 52512 271552
rect 52512 271532 52514 271552
rect 52458 271496 52514 271532
rect 52734 271496 52790 271552
rect 53010 271088 53066 271144
rect 52366 145560 52422 145616
rect 53286 165280 53342 165336
rect 303066 584296 303122 584352
rect 302882 554784 302938 554840
rect 302790 515480 302846 515536
rect 302882 500520 302938 500576
rect 305642 555328 305698 555384
rect 53746 388456 53802 388512
rect 54758 485424 54814 485480
rect 54482 377984 54538 378040
rect 54574 272856 54630 272912
rect 53838 250960 53894 251016
rect 54574 270544 54630 270600
rect 54390 250960 54446 251016
rect 54574 145560 54630 145616
rect 56322 490048 56378 490104
rect 56230 471280 56286 471336
rect 55494 380976 55550 381032
rect 54850 145832 54906 145888
rect 56690 311072 56746 311128
rect 56690 204176 56746 204232
rect 56690 202952 56746 203008
rect 56322 165144 56378 165200
rect 56506 145696 56562 145752
rect 57242 417560 57298 417616
rect 57242 389000 57298 389056
rect 56966 301552 57022 301608
rect 57150 310392 57206 310448
rect 56782 175072 56838 175128
rect 57794 417832 57850 417888
rect 57794 414160 57850 414216
rect 57794 413208 57850 413264
rect 57794 411440 57850 411496
rect 57794 410352 57850 410408
rect 57794 408584 57850 408640
rect 57702 391584 57758 391640
rect 57426 389272 57482 389328
rect 57334 306720 57390 306776
rect 57150 204176 57206 204232
rect 57058 203904 57114 203960
rect 56966 195200 57022 195256
rect 56690 96464 56746 96520
rect 57150 198736 57206 198792
rect 57058 97416 57114 97472
rect 58346 390632 58402 390688
rect 57886 311072 57942 311128
rect 57702 310392 57758 310448
rect 57610 307808 57666 307864
rect 57518 304952 57574 305008
rect 57426 303864 57482 303920
rect 57334 199824 57390 199880
rect 57334 198736 57390 198792
rect 57518 282240 57574 282296
rect 58806 284144 58862 284200
rect 58714 281968 58770 282024
rect 58714 270544 58770 270600
rect 57886 203904 57942 203960
rect 57610 200776 57666 200832
rect 57518 197376 57574 197432
rect 57426 196288 57482 196344
rect 57242 175344 57298 175400
rect 57150 93336 57206 93392
rect 57518 163240 57574 163296
rect 57702 197376 57758 197432
rect 57610 93744 57666 93800
rect 57794 195200 57850 195256
rect 57702 91024 57758 91080
rect 57426 90480 57482 90536
rect 57886 175344 57942 175400
rect 57794 88168 57850 88224
rect 57518 70080 57574 70136
rect 58530 251096 58586 251152
rect 58898 177520 58954 177576
rect 58530 145968 58586 146024
rect 57886 68856 57942 68912
rect 2778 19352 2834 19408
rect 59358 357312 59414 357368
rect 59634 272584 59690 272640
rect 59910 471416 59966 471472
rect 59450 164192 59506 164248
rect 59450 140800 59506 140856
rect 66350 490592 66406 490648
rect 65890 471688 65946 471744
rect 68926 490592 68982 490648
rect 68650 490320 68706 490376
rect 68098 467064 68154 467120
rect 69846 469784 69902 469840
rect 70674 468832 70730 468888
rect 70306 468696 70362 468752
rect 71594 491136 71650 491192
rect 71778 491136 71834 491192
rect 72054 490864 72110 490920
rect 72238 491000 72294 491056
rect 73802 490728 73858 490784
rect 74630 490456 74686 490512
rect 73342 490184 73398 490240
rect 75090 466384 75146 466440
rect 76010 466248 76066 466304
rect 77758 491136 77814 491192
rect 77298 491000 77354 491056
rect 76838 466112 76894 466168
rect 76470 465976 76526 466032
rect 78678 490592 78734 490648
rect 78218 465840 78274 465896
rect 79966 468560 80022 468616
rect 80794 485560 80850 485616
rect 82634 471144 82690 471200
rect 80426 468424 80482 468480
rect 79046 465704 79102 465760
rect 91006 471552 91062 471608
rect 90546 471280 90602 471336
rect 69386 465568 69442 465624
rect 92754 471416 92810 471472
rect 116490 485288 116546 485344
rect 117410 485424 117466 485480
rect 120446 488144 120502 488200
rect 120078 488008 120134 488064
rect 121366 488280 121422 488336
rect 120906 487872 120962 487928
rect 118698 485152 118754 485208
rect 118238 485016 118294 485072
rect 107750 465704 107806 465760
rect 122194 474000 122250 474056
rect 126610 487736 126666 487792
rect 125322 482296 125378 482352
rect 124034 482160 124090 482216
rect 128450 482432 128506 482488
rect 145102 490456 145158 490512
rect 145562 479440 145618 479496
rect 146482 490592 146538 490648
rect 146942 482160 146998 482216
rect 146022 474272 146078 474328
rect 147770 490728 147826 490784
rect 149150 489096 149206 489152
rect 151266 483656 151322 483712
rect 150438 480936 150494 480992
rect 148690 476720 148746 476776
rect 152646 485016 152702 485072
rect 153934 475360 153990 475416
rect 151726 474136 151782 474192
rect 155682 482432 155738 482488
rect 156142 482296 156198 482352
rect 158810 483792 158866 483848
rect 158350 478080 158406 478136
rect 157062 476856 157118 476912
rect 160558 471280 160614 471336
rect 154854 468560 154910 468616
rect 147310 468424 147366 468480
rect 162766 471416 162822 471472
rect 163594 471144 163650 471200
rect 161846 468832 161902 468888
rect 165802 474408 165858 474464
rect 167182 465976 167238 466032
rect 169850 468696 169906 468752
rect 172886 472504 172942 472560
rect 173346 471824 173402 471880
rect 172426 471688 172482 471744
rect 171138 467064 171194 467120
rect 178038 466556 178040 466576
rect 178040 466556 178092 466576
rect 178092 466556 178094 466576
rect 178038 466520 178094 466556
rect 179418 466540 179474 466576
rect 179418 466520 179420 466540
rect 179420 466520 179472 466540
rect 179472 466520 179474 466540
rect 179970 490864 180026 490920
rect 180062 466112 180118 466168
rect 168930 465840 168986 465896
rect 181258 468968 181314 469024
rect 182546 471552 182602 471608
rect 92294 464344 92350 464400
rect 184754 491000 184810 491056
rect 185674 491136 185730 491192
rect 186962 490320 187018 490376
rect 190918 466520 190974 466576
rect 183466 464344 183522 464400
rect 110970 380316 111026 380352
rect 110970 380296 110972 380316
rect 110972 380296 111024 380316
rect 111024 380296 111026 380316
rect 113546 380332 113548 380352
rect 113548 380332 113600 380352
rect 113600 380332 113602 380352
rect 113546 380296 113602 380332
rect 115938 380296 115994 380352
rect 118330 380296 118386 380352
rect 120998 380296 121054 380352
rect 123482 380296 123538 380352
rect 128358 380296 128414 380352
rect 135902 380296 135958 380352
rect 143630 380296 143686 380352
rect 148598 380316 148654 380352
rect 148598 380296 148600 380316
rect 148600 380296 148652 380316
rect 148652 380296 148654 380316
rect 99378 380160 99434 380216
rect 155958 380296 156014 380352
rect 158534 380296 158590 380352
rect 160926 380296 160982 380352
rect 163502 380332 163504 380352
rect 163504 380332 163556 380352
rect 163556 380332 163558 380352
rect 163502 380296 163558 380332
rect 166078 380296 166134 380352
rect 77206 379344 77262 379400
rect 80426 379344 80482 379400
rect 85486 379364 85542 379400
rect 85486 379344 85488 379364
rect 85488 379344 85540 379364
rect 85540 379344 85542 379364
rect 76838 379208 76894 379264
rect 76838 378800 76894 378856
rect 86590 379380 86592 379400
rect 86592 379380 86644 379400
rect 86644 379380 86646 379400
rect 86590 379344 86646 379380
rect 88338 379344 88394 379400
rect 88798 379344 88854 379400
rect 90730 379344 90786 379400
rect 91374 379344 91430 379400
rect 92386 379344 92442 379400
rect 93582 379344 93638 379400
rect 96066 379344 96122 379400
rect 98458 379344 98514 379400
rect 90822 379208 90878 379264
rect 93490 379208 93546 379264
rect 80426 378664 80482 378720
rect 77114 378528 77170 378584
rect 101034 379344 101090 379400
rect 103518 379344 103574 379400
rect 105358 379344 105414 379400
rect 108210 379344 108266 379400
rect 108854 379344 108910 379400
rect 109774 379344 109830 379400
rect 111246 379344 111302 379400
rect 112350 379344 112406 379400
rect 113454 379344 113510 379400
rect 114466 379344 114522 379400
rect 115846 379344 115902 379400
rect 117134 379344 117190 379400
rect 141054 379344 141110 379400
rect 146022 379344 146078 379400
rect 150990 379344 151046 379400
rect 153566 379344 153622 379400
rect 99470 379208 99526 379264
rect 97078 378528 97134 378584
rect 98550 378528 98606 378584
rect 102966 379208 103022 379264
rect 101862 378528 101918 378584
rect 100758 378256 100814 378312
rect 104254 379208 104310 379264
rect 107566 378528 107622 378584
rect 125966 378392 126022 378448
rect 131026 378392 131082 378448
rect 133510 378392 133566 378448
rect 138478 378392 138534 378448
rect 108854 377712 108910 377768
rect 182362 378392 182418 378448
rect 182270 378256 182326 378312
rect 182822 378256 182878 378312
rect 178590 358828 178646 358864
rect 178590 358808 178592 358828
rect 178592 358808 178644 358828
rect 178644 358808 178646 358828
rect 179694 358844 179696 358864
rect 179696 358844 179748 358864
rect 179748 358844 179750 358864
rect 179694 358808 179750 358844
rect 197358 490184 197414 490240
rect 190918 358808 190974 358864
rect 95974 273808 96030 273864
rect 77114 273128 77170 273184
rect 88338 273128 88394 273184
rect 90730 273128 90786 273184
rect 93674 273128 93730 273184
rect 60922 272448 60978 272504
rect 60738 252456 60794 252512
rect 95698 272720 95754 272776
rect 95882 272720 95938 272776
rect 83002 272332 83058 272368
rect 83002 272312 83004 272332
rect 83004 272312 83056 272332
rect 83056 272312 83058 272332
rect 95698 272312 95754 272368
rect 131026 273672 131082 273728
rect 145930 273692 145986 273728
rect 145930 273672 145932 273692
rect 145932 273672 145984 273692
rect 145984 273672 145986 273692
rect 133418 273556 133474 273592
rect 133418 273536 133420 273556
rect 133420 273536 133472 273556
rect 133472 273536 133474 273556
rect 135902 273536 135958 273592
rect 138478 273536 138534 273592
rect 140870 273536 140926 273592
rect 98090 273128 98146 273184
rect 98458 272856 98514 272912
rect 99378 272856 99434 272912
rect 85394 272196 85450 272232
rect 85394 272176 85396 272196
rect 85396 272176 85448 272196
rect 85448 272176 85450 272196
rect 113546 272176 113602 272232
rect 75918 271768 75974 271824
rect 84198 271768 84254 271824
rect 88338 271768 88394 271824
rect 94226 271768 94282 271824
rect 102138 271768 102194 271824
rect 107658 271768 107714 271824
rect 67546 271496 67602 271552
rect 77298 271360 77354 271416
rect 78678 270972 78734 271008
rect 78678 270952 78680 270972
rect 78680 270952 78732 270972
rect 78732 270952 78734 270972
rect 103518 271632 103574 271688
rect 110418 271632 110474 271688
rect 100758 271496 100814 271552
rect 91190 271360 91246 271416
rect 85578 270680 85634 270736
rect 89718 270680 89774 270736
rect 86958 270544 87014 270600
rect 91098 270544 91154 270600
rect 104898 271360 104954 271416
rect 125598 271788 125654 271824
rect 125598 271768 125600 271788
rect 125600 271768 125652 271788
rect 125652 271768 125654 271788
rect 143538 271804 143540 271824
rect 143540 271804 143592 271824
rect 143592 271804 143594 271824
rect 143538 271768 143594 271804
rect 154486 271804 154488 271824
rect 154488 271804 154540 271824
rect 154540 271804 154542 271824
rect 154486 271768 154542 271804
rect 157246 271788 157302 271824
rect 157246 271768 157248 271788
rect 157248 271768 157300 271788
rect 157300 271768 157302 271788
rect 158626 271768 158682 271824
rect 120078 271652 120134 271688
rect 120078 271632 120080 271652
rect 120080 271632 120132 271652
rect 120132 271632 120134 271652
rect 123114 271632 123170 271688
rect 161386 271632 161442 271688
rect 164146 271632 164202 271688
rect 115938 271496 115994 271552
rect 117318 271516 117374 271552
rect 198738 460128 198794 460184
rect 198646 396616 198702 396672
rect 198554 380976 198610 381032
rect 117318 271496 117320 271516
rect 117320 271496 117372 271516
rect 117372 271496 117374 271516
rect 183466 271360 183522 271416
rect 106278 271224 106334 271280
rect 104898 270952 104954 271008
rect 96618 270816 96674 270872
rect 92478 270680 92534 270736
rect 103702 270544 103758 270600
rect 128358 271088 128414 271144
rect 183466 271124 183468 271144
rect 183468 271124 183520 271144
rect 183520 271124 183522 271144
rect 183466 271088 183522 271124
rect 115938 270816 115994 270872
rect 106370 270544 106426 270600
rect 107658 270544 107714 270600
rect 110418 270544 110474 270600
rect 113178 270564 113234 270600
rect 113178 270544 113180 270564
rect 113180 270544 113232 270564
rect 113232 270544 113234 270564
rect 114466 270544 114522 270600
rect 115846 270544 115902 270600
rect 147678 270816 147734 270872
rect 180154 253308 180156 253328
rect 180156 253308 180208 253328
rect 180208 253308 180210 253328
rect 180154 253272 180210 253308
rect 179326 253172 179328 253192
rect 179328 253172 179380 253192
rect 179380 253172 179382 253192
rect 179326 253136 179382 253172
rect 191746 252612 191802 252648
rect 191746 252592 191748 252612
rect 191748 252592 191800 252612
rect 191800 252592 191802 252612
rect 138478 166776 138534 166832
rect 143538 166776 143594 166832
rect 145930 166776 145986 166832
rect 98458 166640 98514 166696
rect 101034 166640 101090 166696
rect 105818 166640 105874 166696
rect 108210 166640 108266 166696
rect 163318 166640 163374 166696
rect 165894 166640 165950 166696
rect 113270 166504 113326 166560
rect 150898 166524 150954 166560
rect 150898 166504 150900 166524
rect 150900 166504 150952 166524
rect 150952 166504 150954 166524
rect 96066 166252 96122 166288
rect 96066 166232 96068 166252
rect 96068 166232 96120 166252
rect 96120 166232 96122 166252
rect 153290 166504 153346 166560
rect 81438 165552 81494 165608
rect 84290 165552 84346 165608
rect 89902 165552 89958 165608
rect 91098 165552 91154 165608
rect 95238 165552 95294 165608
rect 99378 165552 99434 165608
rect 103518 165552 103574 165608
rect 109682 165552 109738 165608
rect 110878 165552 110934 165608
rect 111154 165552 111210 165608
rect 111890 165552 111946 165608
rect 113546 165552 113602 165608
rect 115938 165552 115994 165608
rect 116398 165552 116454 165608
rect 117870 165552 117926 165608
rect 118330 165552 118386 165608
rect 120906 165552 120962 165608
rect 123482 165552 123538 165608
rect 125874 165552 125930 165608
rect 128358 165552 128414 165608
rect 129738 165552 129794 165608
rect 132498 165572 132554 165608
rect 132498 165552 132500 165572
rect 132500 165552 132552 165572
rect 132552 165552 132554 165572
rect 76010 164328 76066 164384
rect 75918 164192 75974 164248
rect 77298 164192 77354 164248
rect 78678 164192 78734 164248
rect 80058 164192 80114 164248
rect 82818 164192 82874 164248
rect 84198 164192 84254 164248
rect 88338 164756 88394 164792
rect 88338 164736 88340 164756
rect 88340 164736 88392 164756
rect 88392 164736 88394 164756
rect 85578 164192 85634 164248
rect 86958 164192 87014 164248
rect 88430 164192 88486 164248
rect 89810 164192 89866 164248
rect 91190 164192 91246 164248
rect 92478 164192 92534 164248
rect 93858 164192 93914 164248
rect 91098 145968 91154 146024
rect 96618 164192 96674 164248
rect 96618 145832 96674 145888
rect 97998 164192 98054 164248
rect 97262 145696 97318 145752
rect 104898 164892 104954 164928
rect 104898 164872 104900 164892
rect 104900 164872 104952 164892
rect 104952 164872 104954 164892
rect 107566 164872 107622 164928
rect 106278 164736 106334 164792
rect 100758 164464 100814 164520
rect 100758 164192 100814 164248
rect 102138 164192 102194 164248
rect 103610 164192 103666 164248
rect 99378 145560 99434 145616
rect 107750 164484 107806 164520
rect 107750 164464 107752 164484
rect 107752 164464 107804 164484
rect 107804 164464 107806 164484
rect 114466 164872 114522 164928
rect 116030 164464 116086 164520
rect 183190 165552 183246 165608
rect 118882 165008 118938 165064
rect 183466 165028 183522 165064
rect 183466 165008 183468 165028
rect 183468 165008 183520 165028
rect 183520 165008 183522 165028
rect 191746 145424 191802 145480
rect 179050 144880 179106 144936
rect 179694 144880 179750 144936
rect 77114 59780 77116 59800
rect 77116 59780 77168 59800
rect 77168 59780 77170 59800
rect 77114 59744 77170 59780
rect 83094 59744 83150 59800
rect 84198 59764 84254 59800
rect 84198 59744 84200 59764
rect 84200 59744 84252 59764
rect 84252 59744 84254 59764
rect 99470 59744 99526 59800
rect 102782 59744 102838 59800
rect 107566 59744 107622 59800
rect 100758 59644 100760 59664
rect 100760 59644 100812 59664
rect 100812 59644 100814 59664
rect 100758 59608 100814 59644
rect 103886 59608 103942 59664
rect 85394 59356 85450 59392
rect 85394 59336 85396 59356
rect 85396 59336 85448 59356
rect 85448 59336 85450 59356
rect 95882 59336 95938 59392
rect 98090 59336 98146 59392
rect 114374 59608 114430 59664
rect 143538 59608 143594 59664
rect 105266 59336 105322 59392
rect 106370 59336 106426 59392
rect 138386 59064 138442 59120
rect 148506 59200 148562 59256
rect 150898 59200 150954 59256
rect 76010 57840 76066 57896
rect 78218 57840 78274 57896
rect 78678 57840 78734 57896
rect 80426 57840 80482 57896
rect 81438 57840 81494 57896
rect 86498 57840 86554 57896
rect 86958 57840 87014 57896
rect 88338 57840 88394 57896
rect 89994 57840 90050 57896
rect 90730 57840 90786 57896
rect 91190 57840 91246 57896
rect 92202 57840 92258 57896
rect 92478 57840 92534 57896
rect 93674 57840 93730 57896
rect 94410 57840 94466 57896
rect 98458 57840 98514 57896
rect 101770 57840 101826 57896
rect 108578 57840 108634 57896
rect 109498 57840 109554 57896
rect 111154 57840 111210 57896
rect 113546 57840 113602 57896
rect 116490 57840 116546 57896
rect 117962 57840 118018 57896
rect 120722 57840 120778 57896
rect 123482 57840 123538 57896
rect 130842 57840 130898 57896
rect 145562 57860 145618 57896
rect 145562 57840 145564 57860
rect 145564 57840 145616 57860
rect 145616 57840 145618 57860
rect 88430 57024 88486 57080
rect 98642 57432 98698 57488
rect 98642 57160 98698 57216
rect 114558 57568 114614 57624
rect 111798 57432 111854 57488
rect 113178 57432 113234 57488
rect 118698 57568 118754 57624
rect 116490 56072 116546 56128
rect 153290 57840 153346 57896
rect 183466 57860 183522 57896
rect 183466 57840 183468 57860
rect 183468 57840 183520 57860
rect 183520 57840 183522 57860
rect 198922 400288 198978 400344
rect 198922 395256 198978 395312
rect 199198 397296 199254 397352
rect 199566 398248 199622 398304
rect 199474 397296 199530 397352
rect 198830 353096 198886 353152
rect 198738 291624 198794 291680
rect 199198 292712 199254 292768
rect 198922 290944 198978 291000
rect 198830 246200 198886 246256
rect 198738 184864 198794 184920
rect 198738 183504 198794 183560
rect 199106 289720 199162 289776
rect 199106 288768 199162 288824
rect 199014 288360 199070 288416
rect 199014 287544 199070 287600
rect 198922 183504 198978 183560
rect 198922 182008 198978 182064
rect 198830 139168 198886 139224
rect 198738 76336 198794 76392
rect 199842 394576 199898 394632
rect 199382 291624 199438 291680
rect 199566 292712 199622 292768
rect 199474 290944 199530 291000
rect 199658 289720 199714 289776
rect 199750 288360 199806 288416
rect 200762 490900 200764 490920
rect 200764 490900 200816 490920
rect 200816 490900 200818 490920
rect 200762 490864 200818 490900
rect 200578 490320 200634 490376
rect 201406 380976 201462 381032
rect 199290 186360 199346 186416
rect 199198 184864 199254 184920
rect 199106 182008 199162 182064
rect 199014 180648 199070 180704
rect 198922 74840 198978 74896
rect 199290 79328 199346 79384
rect 199198 77696 199254 77752
rect 199106 73616 199162 73672
rect 201590 491036 201592 491056
rect 201592 491036 201644 491056
rect 201644 491036 201646 491056
rect 201590 491000 201646 491036
rect 202878 490592 202934 490648
rect 202234 471280 202290 471336
rect 202418 471416 202474 471472
rect 202510 270408 202566 270464
rect 204258 490900 204260 490920
rect 204260 490900 204312 490920
rect 204312 490900 204314 490920
rect 204258 490864 204314 490900
rect 204258 490492 204260 490512
rect 204260 490492 204312 490512
rect 204312 490492 204314 490512
rect 204258 490456 204314 490492
rect 204258 379072 204314 379128
rect 204258 378392 204314 378448
rect 205638 491036 205640 491056
rect 205640 491036 205692 491056
rect 205692 491036 205694 491056
rect 205638 491000 205694 491036
rect 205638 490320 205694 490376
rect 204718 380160 204774 380216
rect 204718 379888 204774 379944
rect 204718 378936 204774 378992
rect 204810 378528 204866 378584
rect 204718 378120 204774 378176
rect 203522 165416 203578 165472
rect 205178 464344 205234 464400
rect 205914 380160 205970 380216
rect 205730 379072 205786 379128
rect 205546 378256 205602 378312
rect 205362 377848 205418 377904
rect 205454 377712 205510 377768
rect 207018 380704 207074 380760
rect 207018 380296 207074 380352
rect 207018 379072 207074 379128
rect 206466 271496 206522 271552
rect 207294 374584 207350 374640
rect 208398 490320 208454 490376
rect 208306 379908 208362 379944
rect 208306 379888 208308 379908
rect 208308 379888 208360 379908
rect 208360 379888 208362 379908
rect 208122 378392 208178 378448
rect 207754 270952 207810 271008
rect 208122 270272 208178 270328
rect 209226 471144 209282 471200
rect 209870 378936 209926 378992
rect 209686 378528 209742 378584
rect 210330 378800 210386 378856
rect 211066 379480 211122 379536
rect 210974 378120 211030 378176
rect 183190 57740 183192 57760
rect 183192 57740 183244 57760
rect 183244 57740 183246 57760
rect 183190 57704 183246 57740
rect 155958 57568 156014 57624
rect 160098 57568 160154 57624
rect 165618 57568 165674 57624
rect 153290 56208 153346 56264
rect 212078 491000 212134 491056
rect 212538 490592 212594 490648
rect 211250 380704 211306 380760
rect 212630 380568 212686 380624
rect 212446 378120 212502 378176
rect 212446 377984 212502 378040
rect 211710 146104 211766 146160
rect 211802 145832 211858 145888
rect 213366 491136 213422 491192
rect 212998 380432 213054 380488
rect 212998 379752 213054 379808
rect 212998 379344 213054 379400
rect 212998 378936 213054 378992
rect 212906 270136 212962 270192
rect 213642 380704 213698 380760
rect 213826 379208 213882 379264
rect 213826 378936 213882 378992
rect 213550 271360 213606 271416
rect 213826 377984 213882 378040
rect 165618 55120 165674 55176
rect 212170 55120 212226 55176
rect 160098 54984 160154 55040
rect 155958 54848 156014 54904
rect 118698 54712 118754 54768
rect 214378 380024 214434 380080
rect 214102 271768 214158 271824
rect 214470 270136 214526 270192
rect 215114 376624 215170 376680
rect 215022 376488 215078 376544
rect 214194 146240 214250 146296
rect 214838 146240 214894 146296
rect 214838 146104 214894 146160
rect 214838 145560 214894 145616
rect 215298 380296 215354 380352
rect 215390 377848 215446 377904
rect 216218 271632 216274 271688
rect 216770 417832 216826 417888
rect 216862 416880 216918 416936
rect 216862 414704 216918 414760
rect 216678 413752 216734 413808
rect 216770 409148 216826 409184
rect 216770 409128 216772 409148
rect 216772 409128 216824 409148
rect 216824 409128 216826 409148
rect 217230 410896 217286 410952
rect 216678 389308 216680 389328
rect 216680 389308 216732 389328
rect 216732 389308 216734 389328
rect 216678 389272 216734 389308
rect 216586 377984 216642 378040
rect 216402 145696 216458 145752
rect 216678 374584 216734 374640
rect 216954 390904 217010 390960
rect 216954 389000 217010 389056
rect 216954 307672 217010 307728
rect 217046 304952 217102 305008
rect 217322 379652 217324 379672
rect 217324 379652 217376 379672
rect 217376 379652 217378 379672
rect 217322 379616 217378 379652
rect 217138 303864 217194 303920
rect 217046 302096 217102 302152
rect 216678 284008 216734 284064
rect 216678 282376 216734 282432
rect 216770 282104 216826 282160
rect 216862 202952 216918 203008
rect 216678 176976 216734 177032
rect 216678 175344 216734 175400
rect 216678 175072 216734 175128
rect 216678 162696 216734 162752
rect 217782 417832 217838 417888
rect 217690 411984 217746 412040
rect 217414 375672 217470 375728
rect 217506 310800 217562 310856
rect 217414 309984 217470 310040
rect 217322 302096 217378 302152
rect 217322 270020 217378 270056
rect 217322 270000 217324 270020
rect 217324 270000 217376 270020
rect 217376 270000 217378 270020
rect 217046 195200 217102 195256
rect 217874 416880 217930 416936
rect 217782 310800 217838 310856
rect 217966 379752 218022 379808
rect 217874 309984 217930 310040
rect 217598 307808 217654 307864
rect 217506 203904 217562 203960
rect 217414 202952 217470 203008
rect 217414 198736 217470 198792
rect 216862 95920 216918 95976
rect 216678 68348 216680 68368
rect 216680 68348 216732 68368
rect 216732 68348 216734 68368
rect 216678 68312 216734 68348
rect 216770 68040 216826 68096
rect 217690 307672 217746 307728
rect 217690 306720 217746 306776
rect 217598 200776 217654 200832
rect 217506 96872 217562 96928
rect 217414 92792 217470 92848
rect 217874 304952 217930 305008
rect 217782 303864 217838 303920
rect 217690 199824 217746 199880
rect 217690 198736 217746 198792
rect 217966 252492 217968 252512
rect 217968 252492 218020 252512
rect 218020 252492 218022 252512
rect 217966 252456 218022 252492
rect 217874 198056 217930 198112
rect 217782 196968 217838 197024
rect 217690 195200 217746 195256
rect 217598 93744 217654 93800
rect 217874 91024 217930 91080
rect 217782 89936 217838 89992
rect 217690 88168 217746 88224
rect 218610 162596 218612 162616
rect 218612 162596 218664 162616
rect 218664 162596 218666 162616
rect 218610 162560 218666 162596
rect 218426 146104 218482 146160
rect 218426 144880 218482 144936
rect 218978 468560 219034 468616
rect 218794 468424 218850 468480
rect 218886 163532 218942 163568
rect 218886 163512 218888 163532
rect 218888 163512 218940 163532
rect 218940 163512 218942 163532
rect 218886 162716 218942 162752
rect 218886 162696 218888 162716
rect 218888 162696 218940 162716
rect 218940 162696 218942 162716
rect 219070 465840 219126 465896
rect 219346 379480 219402 379536
rect 219254 377848 219310 377904
rect 219070 59472 219126 59528
rect 223946 480936 224002 480992
rect 224866 491136 224922 491192
rect 226154 490728 226210 490784
rect 225694 490592 225750 490648
rect 226614 490456 226670 490512
rect 228822 487736 228878 487792
rect 229282 486376 229338 486432
rect 229742 485016 229798 485072
rect 228362 483656 228418 483712
rect 230570 490728 230626 490784
rect 231490 490864 231546 490920
rect 232318 490456 232374 490512
rect 231030 475360 231086 475416
rect 230110 474000 230166 474056
rect 234066 490592 234122 490648
rect 234986 491136 235042 491192
rect 235446 482296 235502 482352
rect 236274 491000 236330 491056
rect 235906 479440 235962 479496
rect 234526 476720 234582 476776
rect 233698 472504 233754 472560
rect 224406 465704 224462 465760
rect 247314 489096 247370 489152
rect 253478 481072 253534 481128
rect 252558 475496 252614 475552
rect 255686 478080 255742 478136
rect 276386 468424 276442 468480
rect 295338 471416 295394 471472
rect 296166 471144 296222 471200
rect 297546 471280 297602 471336
rect 316682 647264 316738 647320
rect 321558 643592 321614 643648
rect 321558 638988 321614 639024
rect 321558 638968 321560 638988
rect 321560 638968 321612 638988
rect 321612 638968 321614 638988
rect 321558 634072 321614 634128
rect 321558 629448 321614 629504
rect 321558 625232 321614 625288
rect 321558 619928 321614 619984
rect 321558 615576 321614 615632
rect 321558 610272 321614 610328
rect 321558 600752 321614 600808
rect 321558 596400 321614 596456
rect 321558 591232 321614 591288
rect 321098 585792 321154 585848
rect 321006 582256 321062 582312
rect 321834 576816 321890 576872
rect 321558 571648 321614 571704
rect 321558 567296 321614 567352
rect 321558 562808 321614 562864
rect 324226 606736 324282 606792
rect 316958 553696 317014 553752
rect 321558 557776 321614 557832
rect 319626 553424 319682 553480
rect 319810 553560 319866 553616
rect 321558 553324 321560 553344
rect 321560 553324 321612 553344
rect 321612 553324 321614 553344
rect 321558 553288 321614 553324
rect 321650 548936 321706 548992
rect 321558 543668 321560 543688
rect 321560 543668 321612 543688
rect 321612 543668 321614 543688
rect 321558 543632 321614 543668
rect 321558 539280 321614 539336
rect 322386 555192 322442 555248
rect 322754 532480 322810 532536
rect 333058 646176 333114 646232
rect 351090 646040 351146 646096
rect 423862 647264 423918 647320
rect 410338 645904 410394 645960
rect 433338 630808 433394 630864
rect 433338 611360 433394 611416
rect 323950 555464 324006 555520
rect 323858 532344 323914 532400
rect 342718 532344 342774 532400
rect 360750 532480 360806 532536
rect 338486 466556 338488 466576
rect 338488 466556 338540 466576
rect 338540 466556 338542 466576
rect 338486 466520 338542 466556
rect 339774 466540 339830 466576
rect 339774 466520 339776 466540
rect 339776 466520 339828 466540
rect 339828 466520 339830 466540
rect 350998 466520 351054 466576
rect 298374 465840 298430 465896
rect 235998 380704 236054 380760
rect 237102 380704 237158 380760
rect 243082 380704 243138 380760
rect 248234 380704 248290 380760
rect 254490 380704 254546 380760
rect 255870 380704 255926 380760
rect 313462 380704 313518 380760
rect 220726 380296 220782 380352
rect 244278 380432 244334 380488
rect 220082 379344 220138 379400
rect 219990 379072 220046 379128
rect 220726 379344 220782 379400
rect 239586 379344 239642 379400
rect 220726 378528 220782 378584
rect 220910 378664 220966 378720
rect 238206 379208 238262 379264
rect 258078 380568 258134 380624
rect 261758 380568 261814 380624
rect 270958 380568 271014 380624
rect 244922 379344 244978 379400
rect 246210 379344 246266 379400
rect 248602 379344 248658 379400
rect 250074 379344 250130 379400
rect 251178 379344 251234 379400
rect 252282 379344 252338 379400
rect 253386 379344 253442 379400
rect 263874 379344 263930 379400
rect 264978 379344 265034 379400
rect 268290 379344 268346 379400
rect 269762 379380 269764 379400
rect 269764 379380 269816 379400
rect 269816 379380 269818 379400
rect 269762 379344 269818 379380
rect 250626 378800 250682 378856
rect 253202 378800 253258 378856
rect 258354 378528 258410 378584
rect 260562 378528 260618 378584
rect 260930 378528 260986 378584
rect 253202 378392 253258 378448
rect 253386 378392 253442 378448
rect 255962 378392 256018 378448
rect 262770 378528 262826 378584
rect 263598 378528 263654 378584
rect 265898 378528 265954 378584
rect 266358 378548 266414 378584
rect 266358 378528 266360 378548
rect 266360 378528 266412 378548
rect 266412 378528 266414 378548
rect 267554 378528 267610 378584
rect 268014 378528 268070 378584
rect 315854 380568 315910 380624
rect 271050 379364 271106 379400
rect 271050 379344 271052 379364
rect 271052 379344 271104 379364
rect 271104 379344 271106 379364
rect 272154 379344 272210 379400
rect 273258 379344 273314 379400
rect 275742 379344 275798 379400
rect 285954 379344 286010 379400
rect 287702 379344 287758 379400
rect 290186 379344 290242 379400
rect 293314 379344 293370 379400
rect 295890 379344 295946 379400
rect 298098 379344 298154 379400
rect 305826 379380 305828 379400
rect 305828 379380 305880 379400
rect 305880 379380 305882 379400
rect 305826 379344 305882 379380
rect 307850 379344 307906 379400
rect 310978 379344 311034 379400
rect 317786 379344 317842 379400
rect 320914 379344 320970 379400
rect 325882 379344 325938 379400
rect 273442 378936 273498 378992
rect 274638 378392 274694 378448
rect 276110 379208 276166 379264
rect 277030 379208 277086 379264
rect 278410 379208 278466 379264
rect 280802 379208 280858 379264
rect 283102 379208 283158 379264
rect 276018 378256 276074 378312
rect 277306 378936 277362 378992
rect 280066 378120 280122 378176
rect 300858 379208 300914 379264
rect 302514 378936 302570 378992
rect 343454 379072 343510 379128
rect 343546 378936 343602 378992
rect 338486 358828 338542 358864
rect 338486 358808 338488 358828
rect 338488 358808 338540 358828
rect 338540 358808 338542 358828
rect 339774 358844 339776 358864
rect 339776 358844 339828 358864
rect 339828 358844 339830 358864
rect 339774 358808 339830 358844
rect 351734 358808 351790 358864
rect 250718 273536 250774 273592
rect 272246 273536 272302 273592
rect 280894 273536 280950 273592
rect 273258 273400 273314 273456
rect 283378 272720 283434 272776
rect 288162 272720 288218 272776
rect 290922 272740 290978 272776
rect 290922 272720 290924 272740
rect 290924 272720 290976 272740
rect 290976 272720 290978 272740
rect 295890 272756 295892 272776
rect 295892 272756 295944 272776
rect 295944 272756 295946 272776
rect 295890 272720 295946 272756
rect 298466 272604 298522 272640
rect 298466 272584 298468 272604
rect 298468 272584 298520 272604
rect 298520 272584 298522 272604
rect 300858 272584 300914 272640
rect 235998 272176 236054 272232
rect 255318 271768 255374 271824
rect 263598 271768 263654 271824
rect 264978 271768 265034 271824
rect 268014 271768 268070 271824
rect 270498 271768 270554 271824
rect 273258 271768 273314 271824
rect 275926 271768 275982 271824
rect 276110 271768 276166 271824
rect 277214 271768 277270 271824
rect 278686 271768 278742 271824
rect 302238 271788 302294 271824
rect 302238 271768 302240 271788
rect 302240 271768 302292 271788
rect 302292 271768 302294 271788
rect 258262 271224 258318 271280
rect 260838 271244 260894 271280
rect 260838 271224 260840 271244
rect 260840 271224 260892 271244
rect 260892 271224 260894 271244
rect 307758 271804 307760 271824
rect 307760 271804 307812 271824
rect 307812 271804 307814 271824
rect 307758 271768 307814 271804
rect 343546 271632 343602 271688
rect 343454 271496 343510 271552
rect 280066 271244 280122 271280
rect 280066 271224 280068 271244
rect 280068 271224 280120 271244
rect 280120 271224 280122 271244
rect 239126 271088 239182 271144
rect 247038 271088 247094 271144
rect 252558 271088 252614 271144
rect 260838 271088 260894 271144
rect 266358 271088 266414 271144
rect 268106 271108 268162 271144
rect 268106 271088 268108 271108
rect 268108 271088 268160 271108
rect 268160 271088 268162 271108
rect 235998 270544 236054 270600
rect 237378 270544 237434 270600
rect 219622 167048 219678 167104
rect 219346 58520 219402 58576
rect 252558 270816 252614 270872
rect 244278 270680 244334 270736
rect 251270 270680 251326 270736
rect 242898 270544 242954 270600
rect 244370 270544 244426 270600
rect 245658 270544 245714 270600
rect 247038 270544 247094 270600
rect 248510 270544 248566 270600
rect 249798 270544 249854 270600
rect 251178 270544 251234 270600
rect 259550 270680 259606 270736
rect 253938 270544 253994 270600
rect 255318 270544 255374 270600
rect 256698 270544 256754 270600
rect 258078 270544 258134 270600
rect 259458 270544 259514 270600
rect 229098 268368 229154 268424
rect 230386 268404 230388 268424
rect 230388 268404 230440 268424
rect 230440 268404 230442 268424
rect 230386 268368 230442 268404
rect 270498 271088 270554 271144
rect 262218 270544 262274 270600
rect 263598 270544 263654 270600
rect 264978 270816 265034 270872
rect 265622 270680 265678 270736
rect 269118 270544 269174 270600
rect 273258 270564 273314 270600
rect 273258 270544 273260 270564
rect 273260 270544 273312 270564
rect 273312 270544 273314 270564
rect 340786 253408 340842 253464
rect 339406 253000 339462 253056
rect 351826 253172 351828 253192
rect 351828 253172 351880 253192
rect 351880 253172 351882 253192
rect 351826 253136 351882 253172
rect 231858 251776 231914 251832
rect 298466 166776 298522 166832
rect 303526 166776 303582 166832
rect 288254 166660 288310 166696
rect 288254 166640 288256 166660
rect 288256 166640 288308 166660
rect 288308 166640 288310 166660
rect 295890 166640 295946 166696
rect 253570 166504 253626 166560
rect 265898 166504 265954 166560
rect 270866 166504 270922 166560
rect 308494 166640 308550 166696
rect 315854 166640 315910 166696
rect 236090 165552 236146 165608
rect 238758 165552 238814 165608
rect 242898 165552 242954 165608
rect 247130 165552 247186 165608
rect 258170 165552 258226 165608
rect 260838 165552 260894 165608
rect 273442 165552 273498 165608
rect 276018 165552 276074 165608
rect 278410 165552 278466 165608
rect 280802 165552 280858 165608
rect 285954 165552 286010 165608
rect 293314 165552 293370 165608
rect 300858 165552 300914 165608
rect 310978 165572 311034 165608
rect 310978 165552 310980 165572
rect 310980 165552 311032 165572
rect 311032 165552 311034 165572
rect 235998 164192 236054 164248
rect 237378 164192 237434 164248
rect 240138 164192 240194 164248
rect 241518 164192 241574 164248
rect 237378 145832 237434 145888
rect 247038 164872 247094 164928
rect 244370 164328 244426 164384
rect 244278 164192 244334 164248
rect 245658 164192 245714 164248
rect 249798 164872 249854 164928
rect 255318 164872 255374 164928
rect 258078 164892 258134 164928
rect 258078 164872 258080 164892
rect 258080 164872 258132 164892
rect 258132 164872 258134 164892
rect 251270 164328 251326 164384
rect 256698 164328 256754 164384
rect 248418 164192 248474 164248
rect 249890 164192 249946 164248
rect 251178 164192 251234 164248
rect 252558 164192 252614 164248
rect 253938 164192 253994 164248
rect 255410 164192 255466 164248
rect 259550 164328 259606 164384
rect 259458 164192 259514 164248
rect 263598 165144 263654 165200
rect 266266 165144 266322 165200
rect 262218 164192 262274 164248
rect 263782 164192 263838 164248
rect 271878 165144 271934 165200
rect 267738 165008 267794 165064
rect 266542 164328 266598 164384
rect 266450 164192 266506 164248
rect 267738 164212 267794 164248
rect 267738 164192 267740 164212
rect 267740 164192 267792 164212
rect 267792 164192 267794 164212
rect 269118 164192 269174 164248
rect 270498 164192 270554 164248
rect 269118 146240 269174 146296
rect 266542 146104 266598 146160
rect 270498 145696 270554 145752
rect 275282 165144 275338 165200
rect 280066 165144 280122 165200
rect 325882 165552 325938 165608
rect 343270 165572 343326 165608
rect 343270 165552 343272 165572
rect 343272 165552 343324 165572
rect 343324 165552 343326 165572
rect 273810 164328 273866 164384
rect 274546 164192 274602 164248
rect 276662 164192 276718 164248
rect 277398 164192 277454 164248
rect 276018 148960 276074 149016
rect 276662 148960 276718 149016
rect 276018 148280 276074 148336
rect 343546 164892 343602 164928
rect 343546 164872 343548 164892
rect 343548 164872 343600 164892
rect 343600 164872 343602 164892
rect 325882 164056 325938 164112
rect 271878 145560 271934 145616
rect 357162 148960 357218 149016
rect 338486 144880 338542 144936
rect 340234 144880 340290 144936
rect 351642 144880 351698 144936
rect 255870 59744 255926 59800
rect 260654 59744 260710 59800
rect 261758 59744 261814 59800
rect 262862 59744 262918 59800
rect 263874 59744 263930 59800
rect 256974 59608 257030 59664
rect 308494 59608 308550 59664
rect 259458 59336 259514 59392
rect 295890 59200 295946 59256
rect 298466 59200 298522 59256
rect 303434 59200 303490 59256
rect 222934 58520 222990 58576
rect 222934 58248 222990 58304
rect 236090 57840 236146 57896
rect 238114 57840 238170 57896
rect 238758 57840 238814 57896
rect 240506 57840 240562 57896
rect 241518 57840 241574 57896
rect 242898 57840 242954 57896
rect 244370 57840 244426 57896
rect 245290 57840 245346 57896
rect 245658 57840 245714 57896
rect 247682 57840 247738 57896
rect 248142 57840 248198 57896
rect 248418 57840 248474 57896
rect 249798 57840 249854 57896
rect 251178 57840 251234 57896
rect 251362 57840 251418 57896
rect 253386 57840 253442 57896
rect 253938 57840 253994 57896
rect 271234 57840 271290 57896
rect 271878 57840 271934 57896
rect 273258 57840 273314 57896
rect 275650 57840 275706 57896
rect 278042 57840 278098 57896
rect 279054 57840 279110 57896
rect 287610 57840 287666 57896
rect 293314 57840 293370 57896
rect 300858 57840 300914 57896
rect 305826 57840 305882 57896
rect 310978 57840 311034 57896
rect 313370 57840 313426 57896
rect 315026 57840 315082 57896
rect 318246 57840 318302 57896
rect 325882 57860 325938 57896
rect 325882 57840 325884 57860
rect 325884 57840 325936 57860
rect 325936 57840 325938 57860
rect 235998 56888 236054 56944
rect 263598 57704 263654 57760
rect 265438 57704 265494 57760
rect 266450 57704 266506 57760
rect 268198 57704 268254 57760
rect 268658 57704 268714 57760
rect 269118 57704 269174 57760
rect 266358 57296 266414 57352
rect 265438 56072 265494 56128
rect 273350 57704 273406 57760
rect 276018 57704 276074 57760
rect 273350 55120 273406 55176
rect 343178 57876 343180 57896
rect 343180 57876 343232 57896
rect 343232 57876 343234 57896
rect 343178 57840 343234 57876
rect 343454 57860 343510 57896
rect 343454 57840 343456 57860
rect 343456 57840 343508 57860
rect 343508 57840 343510 57860
rect 359370 460128 359426 460184
rect 359094 400288 359150 400344
rect 359002 398112 359058 398168
rect 358542 273128 358598 273184
rect 358910 290944 358966 291000
rect 359186 288768 359242 288824
rect 359002 245656 359058 245712
rect 358910 183504 358966 183560
rect 359738 396752 359794 396808
rect 359462 353096 359518 353152
rect 359370 292712 359426 292768
rect 359278 288360 359334 288416
rect 359922 395256 359978 395312
rect 359830 394032 359886 394088
rect 359554 292712 359610 292768
rect 359646 291760 359702 291816
rect 359554 288360 359610 288416
rect 359554 287544 359610 287600
rect 359462 245656 359518 245712
rect 359462 186360 359518 186416
rect 359278 184864 359334 184920
rect 359186 181872 359242 181928
rect 359094 179424 359150 179480
rect 359002 139304 359058 139360
rect 359370 183504 359426 183560
rect 359278 78240 359334 78296
rect 359646 184864 359702 184920
rect 359554 180648 359610 180704
rect 359554 179424 359610 179480
rect 359462 79872 359518 79928
rect 359370 76880 359426 76936
rect 359186 75384 359242 75440
rect 359094 74024 359150 74080
rect 361486 379480 361542 379536
rect 315026 56208 315082 56264
rect 276018 54984 276074 55040
rect 143538 3984 143594 4040
rect 136454 3848 136510 3904
rect 132958 3440 133014 3496
rect 129370 3304 129426 3360
rect 140042 3712 140098 3768
rect 150622 3576 150678 3632
rect 433430 601704 433486 601760
rect 433522 586744 433578 586800
rect 433614 572600 433670 572656
rect 434626 538872 434682 538928
rect 433430 534928 433486 534984
rect 429198 532616 429254 532672
rect 434810 640192 434866 640248
rect 434810 596672 434866 596728
rect 397458 529080 397514 529136
rect 364062 270816 364118 270872
rect 363786 164736 363842 164792
rect 366362 472640 366418 472696
rect 365534 272992 365590 273048
rect 369582 376896 369638 376952
rect 369582 270408 369638 270464
rect 369858 379072 369914 379128
rect 369858 378664 369914 378720
rect 369766 376896 369822 376952
rect 369030 145560 369086 145616
rect 371054 379072 371110 379128
rect 371606 379480 371662 379536
rect 371790 273264 371846 273320
rect 371606 269864 371662 269920
rect 371054 163376 371110 163432
rect 372342 378800 372398 378856
rect 372158 270408 372214 270464
rect 372158 269728 372214 269784
rect 373078 377712 373134 377768
rect 373262 465704 373318 465760
rect 371790 146240 371846 146296
rect 372526 145832 372582 145888
rect 373906 377848 373962 377904
rect 374366 271224 374422 271280
rect 375194 375944 375250 376000
rect 375010 270408 375066 270464
rect 374826 165280 374882 165336
rect 375930 270408 375986 270464
rect 377034 417832 377090 417888
rect 377034 411984 377090 412040
rect 376758 410488 376814 410544
rect 376850 390904 376906 390960
rect 376942 389272 376998 389328
rect 376942 389000 376998 389056
rect 376390 269864 376446 269920
rect 377494 411984 377550 412040
rect 377402 410896 377458 410952
rect 377402 409148 377458 409184
rect 377402 409128 377404 409148
rect 377404 409128 377456 409148
rect 377456 409128 377458 409148
rect 376758 375300 376760 375320
rect 376760 375300 376812 375320
rect 376812 375300 376814 375320
rect 376758 375264 376814 375300
rect 376942 310800 376998 310856
rect 376758 282104 376814 282160
rect 376942 284008 376998 284064
rect 376942 282240 376998 282296
rect 376206 165416 376262 165472
rect 376206 145696 376262 145752
rect 376022 68040 376078 68096
rect 376942 203904 376998 203960
rect 376850 198736 376906 198792
rect 376574 146240 376630 146296
rect 376574 145696 376630 145752
rect 377770 416880 377826 416936
rect 378046 416880 378102 416936
rect 377770 414704 377826 414760
rect 377678 413752 377734 413808
rect 377586 310800 377642 310856
rect 377770 307808 377826 307864
rect 377678 306720 377734 306776
rect 377494 304952 377550 305008
rect 377310 302096 377366 302152
rect 377678 303592 377734 303648
rect 377586 199824 377642 199880
rect 377586 198736 377642 198792
rect 377494 198056 377550 198112
rect 377310 195200 377366 195256
rect 377034 176976 377090 177032
rect 376942 175344 376998 175400
rect 377218 175072 377274 175128
rect 377310 163376 377366 163432
rect 377310 162968 377366 163024
rect 376942 96872 376998 96928
rect 376850 92792 376906 92848
rect 376942 69944 376998 70000
rect 376942 68332 376998 68368
rect 376942 68312 376944 68332
rect 376944 68312 376996 68332
rect 376996 68312 376998 68332
rect 377954 409128 378010 409184
rect 377862 303864 377918 303920
rect 377862 303592 377918 303648
rect 378230 379480 378286 379536
rect 378046 309984 378102 310040
rect 377954 302096 378010 302152
rect 377862 202952 377918 203008
rect 377770 200776 377826 200832
rect 377678 196968 377734 197024
rect 377586 195200 377642 195256
rect 377494 91024 377550 91080
rect 378046 202952 378102 203008
rect 378046 162560 378102 162616
rect 377862 95920 377918 95976
rect 377770 93744 377826 93800
rect 377678 89936 377734 89992
rect 377586 88168 377642 88224
rect 580170 683848 580226 683904
rect 456982 639648 457038 639704
rect 436282 635976 436338 636032
rect 436190 626456 436246 626512
rect 436098 621696 436154 621752
rect 436742 615848 436798 615904
rect 436190 592048 436246 592104
rect 436098 553424 436154 553480
rect 434902 544856 434958 544912
rect 436282 581712 436338 581768
rect 436374 577224 436430 577280
rect 436466 567568 436522 567624
rect 436558 563080 436614 563136
rect 436650 558048 436706 558104
rect 477130 639920 477186 639976
rect 488722 639920 488778 639976
rect 506754 639920 506810 639976
rect 457718 633528 457774 633584
rect 457626 627408 457682 627464
rect 512182 636928 512238 636984
rect 512090 630808 512146 630864
rect 511998 624008 512054 624064
rect 457534 621288 457590 621344
rect 512090 617888 512146 617944
rect 457626 614488 457682 614544
rect 457534 608368 457590 608424
rect 457442 602248 457498 602304
rect 457442 596128 457498 596184
rect 436834 548392 436890 548448
rect 511998 605648 512054 605704
rect 483018 493312 483074 493368
rect 512182 611768 512238 611824
rect 512274 599528 512330 599584
rect 513286 592728 513342 592784
rect 512090 526360 512146 526416
rect 511998 482160 512054 482216
rect 457534 480800 457590 480856
rect 498474 466520 498530 466576
rect 499762 466556 499764 466576
rect 499764 466556 499816 466576
rect 499816 466556 499818 466576
rect 499762 466520 499818 466556
rect 510894 466540 510950 466576
rect 510894 466520 510896 466540
rect 510896 466520 510948 466540
rect 510948 466520 510950 466540
rect 413558 380840 413614 380896
rect 421102 380876 421104 380896
rect 421104 380876 421156 380896
rect 421156 380876 421158 380896
rect 421102 380840 421158 380876
rect 425978 380840 426034 380896
rect 433614 380840 433670 380896
rect 436006 380840 436062 380896
rect 380898 380160 380954 380216
rect 379058 271632 379114 271688
rect 379426 273264 379482 273320
rect 378414 145832 378470 145888
rect 379058 145560 379114 145616
rect 378966 60560 379022 60616
rect 404174 380568 404230 380624
rect 405462 380568 405518 380624
rect 413466 380568 413522 380624
rect 438490 380704 438546 380760
rect 440882 380704 440938 380760
rect 443458 380704 443514 380760
rect 448242 380704 448298 380760
rect 445942 380568 445998 380624
rect 503350 380568 503406 380624
rect 396078 379344 396134 379400
rect 396354 379344 396410 379400
rect 398194 379344 398250 379400
rect 399482 379344 399538 379400
rect 405830 379344 405886 379400
rect 407578 379344 407634 379400
rect 408314 379364 408370 379400
rect 408314 379344 408316 379364
rect 408316 379344 408368 379364
rect 408368 379344 408370 379364
rect 381082 378800 381138 378856
rect 381174 378664 381230 378720
rect 402978 379208 403034 379264
rect 410338 379344 410394 379400
rect 411258 379344 411314 379400
rect 412362 379344 412418 379400
rect 420642 379344 420698 379400
rect 428186 379344 428242 379400
rect 431130 379344 431186 379400
rect 434258 379380 434260 379400
rect 434260 379380 434312 379400
rect 434312 379380 434314 379400
rect 434258 379344 434314 379380
rect 437938 379344 437994 379400
rect 451002 379344 451058 379400
rect 453026 379344 453082 379400
rect 455602 379344 455658 379400
rect 460938 379344 460994 379400
rect 463514 379344 463570 379400
rect 473450 379344 473506 379400
rect 480626 379344 480682 379400
rect 485962 379344 486018 379400
rect 408682 378528 408738 378584
rect 409970 378120 410026 378176
rect 381266 375264 381322 375320
rect 414570 379208 414626 379264
rect 415858 379208 415914 379264
rect 416042 379208 416098 379264
rect 422850 379208 422906 379264
rect 419354 379072 419410 379128
rect 418434 378528 418490 378584
rect 416962 378120 417018 378176
rect 418158 378120 418214 378176
rect 421746 378528 421802 378584
rect 422574 378256 422630 378312
rect 421746 375944 421802 376000
rect 423954 378120 424010 378176
rect 425150 378120 425206 378176
rect 426438 378120 426494 378176
rect 430670 378528 430726 378584
rect 436190 378528 436246 378584
rect 428278 378120 428334 378176
rect 432234 378120 432290 378176
rect 435178 378120 435234 378176
rect 381266 374584 381322 374640
rect 438122 378120 438178 378176
rect 438122 377848 438178 377904
rect 435178 374584 435234 374640
rect 465078 379072 465134 379128
rect 470874 378936 470930 378992
rect 467930 378800 467986 378856
rect 474738 378800 474794 378856
rect 477498 378800 477554 378856
rect 483386 378800 483442 378856
rect 503626 379344 503682 379400
rect 498842 358808 498898 358864
rect 500774 358808 500830 358864
rect 510894 358828 510950 358864
rect 510894 358808 510896 358828
rect 510896 358808 510948 358828
rect 510948 358808 510950 358828
rect 440882 273672 440938 273728
rect 416042 273536 416098 273592
rect 427634 273556 427690 273592
rect 427634 273536 427636 273556
rect 427636 273536 427688 273556
rect 427688 273536 427690 273556
rect 433338 273536 433394 273592
rect 430946 273284 431002 273320
rect 430946 273264 430948 273284
rect 430948 273264 431000 273284
rect 431000 273264 431002 273284
rect 423402 272856 423458 272912
rect 423770 272856 423826 272912
rect 426438 272856 426494 272912
rect 428186 272892 428188 272912
rect 428188 272892 428240 272912
rect 428240 272892 428242 272912
rect 428186 272856 428242 272892
rect 468482 272876 468538 272912
rect 468482 272856 468484 272876
rect 468484 272856 468536 272876
rect 468536 272856 468538 272876
rect 470874 272856 470930 272912
rect 478418 272740 478474 272776
rect 478418 272720 478420 272740
rect 478420 272720 478472 272740
rect 478472 272720 478474 272740
rect 480810 272720 480866 272776
rect 473450 272584 473506 272640
rect 475842 272604 475898 272640
rect 475842 272584 475844 272604
rect 475844 272584 475896 272604
rect 475896 272584 475898 272604
rect 401690 272176 401746 272232
rect 455786 272176 455842 272232
rect 396722 271088 396778 271144
rect 396078 270544 396134 270600
rect 397458 270544 397514 270600
rect 398838 270544 398894 270600
rect 400218 270544 400274 270600
rect 403530 271768 403586 271824
rect 425058 271768 425114 271824
rect 428002 271768 428058 271824
rect 440146 271768 440202 271824
rect 447138 271768 447194 271824
rect 449898 271768 449954 271824
rect 452658 271768 452714 271824
rect 458178 271804 458180 271824
rect 458180 271804 458232 271824
rect 458232 271804 458234 271824
rect 402978 270544 403034 270600
rect 442998 271516 443054 271552
rect 442998 271496 443000 271516
rect 443000 271496 443052 271516
rect 443052 271496 443054 271516
rect 458178 271768 458234 271804
rect 460938 271768 460994 271824
rect 503626 271496 503682 271552
rect 418342 271360 418398 271416
rect 434718 271360 434774 271416
rect 445758 271380 445814 271416
rect 445758 271360 445760 271380
rect 445760 271360 445812 271380
rect 445812 271360 445814 271380
rect 503534 271360 503590 271416
rect 433338 271224 433394 271280
rect 437478 271224 437534 271280
rect 420918 271108 420974 271144
rect 420918 271088 420920 271108
rect 420920 271088 420972 271108
rect 420972 271088 420974 271108
rect 409878 270972 409934 271008
rect 409878 270952 409880 270972
rect 409880 270952 409932 270972
rect 409932 270952 409934 270972
rect 429198 270952 429254 271008
rect 437478 270952 437534 271008
rect 411350 270680 411406 270736
rect 404358 270544 404414 270600
rect 405738 270544 405794 270600
rect 407118 270544 407174 270600
rect 408498 270544 408554 270600
rect 409878 270544 409934 270600
rect 411258 270544 411314 270600
rect 413006 270544 413062 270600
rect 414018 270544 414074 270600
rect 415398 270544 415454 270600
rect 418158 270544 418214 270600
rect 418526 270544 418582 270600
rect 419538 270544 419594 270600
rect 420918 270544 420974 270600
rect 431958 270680 432014 270736
rect 436098 270564 436154 270600
rect 436098 270544 436100 270564
rect 436100 270544 436152 270564
rect 436152 270544 436154 270564
rect 500866 253308 500868 253328
rect 500868 253308 500920 253328
rect 500920 253308 500922 253328
rect 500866 253272 500922 253308
rect 499210 252728 499266 252784
rect 510894 252612 510950 252648
rect 510894 252592 510896 252612
rect 510896 252592 510948 252612
rect 510948 252592 510950 252612
rect 389178 251776 389234 251832
rect 416042 166776 416098 166832
rect 418434 166812 418436 166832
rect 418436 166812 418488 166832
rect 418488 166812 418490 166832
rect 418434 166776 418490 166812
rect 423402 166776 423458 166832
rect 425978 166796 426034 166832
rect 425978 166776 425980 166796
rect 425980 166776 426032 166796
rect 426032 166776 426034 166796
rect 470966 166776 471022 166832
rect 473450 166776 473506 166832
rect 475842 166776 475898 166832
rect 478418 166776 478474 166832
rect 480902 166776 480958 166832
rect 413558 166504 413614 166560
rect 408130 166232 408186 166288
rect 397458 165552 397514 165608
rect 401598 165552 401654 165608
rect 404358 165552 404414 165608
rect 410430 165552 410486 165608
rect 396170 164328 396226 164384
rect 396078 164192 396134 164248
rect 380898 146240 380954 146296
rect 395342 146104 395398 146160
rect 398838 164192 398894 164248
rect 400218 164192 400274 164248
rect 402978 164328 403034 164384
rect 403070 164192 403126 164248
rect 483386 166640 483442 166696
rect 485962 166640 486018 166696
rect 503258 166504 503314 166560
rect 428186 166252 428242 166288
rect 428186 166232 428188 166252
rect 428188 166232 428240 166252
rect 428240 166232 428242 166252
rect 415398 165552 415454 165608
rect 416870 165552 416926 165608
rect 418158 165552 418214 165608
rect 423770 165552 423826 165608
rect 426438 165552 426494 165608
rect 434626 165552 434682 165608
rect 411350 164328 411406 164384
rect 405738 164192 405794 164248
rect 407118 164192 407174 164248
rect 408498 164192 408554 164248
rect 409970 164192 410026 164248
rect 411258 164192 411314 164248
rect 412730 164192 412786 164248
rect 414018 164192 414074 164248
rect 420918 164872 420974 164928
rect 418250 164192 418306 164248
rect 419538 164192 419594 164248
rect 420918 164192 420974 164248
rect 423586 164192 423642 164248
rect 415398 146104 415454 146160
rect 425058 164192 425114 164248
rect 433338 164872 433394 164928
rect 433338 164600 433394 164656
rect 427726 164192 427782 164248
rect 423770 145832 423826 145888
rect 423678 145696 423734 145752
rect 429290 164328 429346 164384
rect 430670 164328 430726 164384
rect 429106 164192 429162 164248
rect 430578 164192 430634 164248
rect 431958 164192 432014 164248
rect 434810 165552 434866 165608
rect 437846 165552 437902 165608
rect 440238 165552 440294 165608
rect 442998 165552 443054 165608
rect 447322 165552 447378 165608
rect 449898 165552 449954 165608
rect 452658 165572 452714 165608
rect 452658 165552 452660 165572
rect 452660 165552 452712 165572
rect 452712 165552 452714 165572
rect 437754 165008 437810 165064
rect 434810 164192 434866 164248
rect 436098 164192 436154 164248
rect 455418 165552 455474 165608
rect 458362 165552 458418 165608
rect 445758 165028 445814 165064
rect 445758 165008 445760 165028
rect 445760 165008 445812 165028
rect 445812 165008 445814 165028
rect 440146 164192 440202 164248
rect 503626 164600 503682 164656
rect 429198 146240 429254 146296
rect 427818 145560 427874 145616
rect 510618 146104 510674 146160
rect 518898 459584 518954 459640
rect 519450 459584 519506 459640
rect 519358 400288 519414 400344
rect 518990 398112 519046 398168
rect 519174 396752 519230 396808
rect 519082 395256 519138 395312
rect 518898 291624 518954 291680
rect 518898 186360 518954 186416
rect 498658 144880 498714 144936
rect 499854 144880 499910 144936
rect 440238 144064 440294 144120
rect 396078 59764 396134 59800
rect 396078 59744 396080 59764
rect 396080 59744 396132 59764
rect 396132 59744 396134 59764
rect 397090 59744 397146 59800
rect 403070 59744 403126 59800
rect 413558 59744 413614 59800
rect 415858 59744 415914 59800
rect 419446 59744 419502 59800
rect 423494 59608 423550 59664
rect 503258 59608 503314 59664
rect 398194 59356 398250 59392
rect 398194 59336 398196 59356
rect 398196 59336 398248 59356
rect 398248 59336 398250 59356
rect 410706 59336 410762 59392
rect 416962 59336 417018 59392
rect 418158 59336 418214 59392
rect 421010 59336 421066 59392
rect 421746 59336 421802 59392
rect 425242 59336 425298 59392
rect 425978 59336 426034 59392
rect 428186 59336 428242 59392
rect 468482 59336 468538 59392
rect 398838 57840 398894 57896
rect 400402 57840 400458 57896
rect 401598 57840 401654 57896
rect 404082 57840 404138 57896
rect 404358 57840 404414 57896
rect 405830 57840 405886 57896
rect 407118 57840 407174 57896
rect 408314 57840 408370 57896
rect 408682 57840 408738 57896
rect 409878 57840 409934 57896
rect 411350 57840 411406 57896
rect 413466 57840 413522 57896
rect 414570 57840 414626 57896
rect 418434 57840 418490 57896
rect 422850 57840 422906 57896
rect 423678 57840 423734 57896
rect 426530 57840 426586 57896
rect 427634 57840 427690 57896
rect 427818 57840 427874 57896
rect 429658 57840 429714 57896
rect 430946 57840 431002 57896
rect 431958 57840 432014 57896
rect 433338 57840 433394 57896
rect 433522 57840 433578 57896
rect 435086 57840 435142 57896
rect 435914 57840 435970 57896
rect 438490 57840 438546 57896
rect 460938 57840 460994 57896
rect 465906 57840 465962 57896
rect 470874 57840 470930 57896
rect 475842 57876 475844 57896
rect 475844 57876 475896 57896
rect 475896 57876 475898 57896
rect 475842 57840 475898 57876
rect 480626 57860 480682 57896
rect 480626 57840 480628 57860
rect 480628 57840 480680 57860
rect 480680 57840 480682 57860
rect 411258 56888 411314 56944
rect 430578 57024 430634 57080
rect 433430 57432 433486 57488
rect 433706 57432 433762 57488
rect 433430 57024 433486 57080
rect 436098 57432 436154 57488
rect 483386 57840 483442 57896
rect 503350 57876 503352 57896
rect 503352 57876 503404 57896
rect 503404 57876 503406 57896
rect 503350 57840 503406 57876
rect 519266 394032 519322 394088
rect 519266 352824 519322 352880
rect 519082 288768 519138 288824
rect 518990 184728 519046 184784
rect 519174 287544 519230 287600
rect 519082 181872 519138 181928
rect 518990 79872 519046 79928
rect 580354 630808 580410 630864
rect 580262 577632 580318 577688
rect 578882 511264 578938 511320
rect 580262 458088 580318 458144
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 519450 352824 519506 352880
rect 519358 293800 519414 293856
rect 519266 246200 519322 246256
rect 519174 180648 519230 180704
rect 519082 75384 519138 75440
rect 519542 290264 519598 290320
rect 580170 351872 580226 351928
rect 580262 325216 580318 325272
rect 520186 288768 520242 288824
rect 519358 186360 519414 186416
rect 519266 139304 519322 139360
rect 580354 272176 580410 272232
rect 580262 232328 580318 232384
rect 580354 192480 580410 192536
rect 520186 184728 520242 184784
rect 519450 183368 519506 183424
rect 520094 183368 520150 183424
rect 519358 78240 519414 78296
rect 580262 152632 580318 152688
rect 520186 79872 520242 79928
rect 519450 76744 519506 76800
rect 519174 74160 519230 74216
rect 438858 57432 438914 57488
rect 438858 55120 438914 55176
rect 427818 54984 427874 55040
rect 580446 112784 580502 112840
rect 580354 72936 580410 72992
rect 580262 33088 580318 33144
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect 316677 647322 316743 647325
rect 423857 647322 423923 647325
rect 316677 647320 423923 647322
rect 316677 647264 316682 647320
rect 316738 647264 423862 647320
rect 423918 647264 423923 647320
rect 316677 647262 423923 647264
rect 316677 647259 316743 647262
rect 423857 647259 423923 647262
rect 54334 646172 54340 646236
rect 54404 646234 54410 646236
rect 333053 646234 333119 646237
rect 54404 646232 333119 646234
rect 54404 646176 333058 646232
rect 333114 646176 333119 646232
rect 54404 646174 333119 646176
rect 54404 646172 54410 646174
rect 333053 646171 333119 646174
rect 51574 646036 51580 646100
rect 51644 646098 51650 646100
rect 351085 646098 351151 646101
rect 51644 646096 351151 646098
rect 51644 646040 351090 646096
rect 351146 646040 351151 646096
rect 51644 646038 351151 646040
rect 51644 646036 51650 646038
rect 351085 646035 351151 646038
rect 53046 645900 53052 645964
rect 53116 645962 53122 645964
rect 410333 645962 410399 645965
rect 53116 645960 410399 645962
rect 53116 645904 410338 645960
rect 410394 645904 410399 645960
rect 53116 645902 410399 645904
rect 53116 645900 53122 645902
rect 410333 645899 410399 645902
rect -960 644996 480 645236
rect 321553 643650 321619 643653
rect 325006 643650 325066 644232
rect 583520 643908 584960 644148
rect 321553 643648 325066 643650
rect 321553 643592 321558 643648
rect 321614 643592 325066 643648
rect 321553 643590 325066 643592
rect 321553 643587 321619 643590
rect 237373 640794 237439 640797
rect 237373 640792 240242 640794
rect 237373 640736 237378 640792
rect 237434 640736 240242 640792
rect 237373 640734 240242 640736
rect 237373 640731 237439 640734
rect 57697 640658 57763 640661
rect 146293 640658 146359 640661
rect 57697 640656 60076 640658
rect 57697 640600 57702 640656
rect 57758 640600 60076 640656
rect 57697 640598 60076 640600
rect 146293 640656 150052 640658
rect 146293 640600 146298 640656
rect 146354 640600 150052 640656
rect 240182 640628 240242 640734
rect 146293 640598 150052 640600
rect 57697 640595 57763 640598
rect 146293 640595 146359 640598
rect 434805 640250 434871 640253
rect 433750 640248 434871 640250
rect 433750 640192 434810 640248
rect 434866 640192 434871 640248
rect 433750 640190 434871 640192
rect 433750 640152 433810 640190
rect 434805 640187 434871 640190
rect 122925 639978 122991 639981
rect 120796 639976 122991 639978
rect 120796 639920 122930 639976
rect 122986 639920 122991 639976
rect 120796 639918 122991 639920
rect 122925 639915 122991 639918
rect 210742 639434 210802 639948
rect 211245 639434 211311 639437
rect 210742 639432 211311 639434
rect 210742 639376 211250 639432
rect 211306 639376 211311 639432
rect 210742 639374 211311 639376
rect 300718 639434 300778 639948
rect 476062 639916 476068 639980
rect 476132 639978 476138 639980
rect 477125 639978 477191 639981
rect 476132 639976 477191 639978
rect 476132 639920 477130 639976
rect 477186 639920 477191 639976
rect 476132 639918 477191 639920
rect 476132 639916 476138 639918
rect 477125 639915 477191 639918
rect 488574 639916 488580 639980
rect 488644 639978 488650 639980
rect 488717 639978 488783 639981
rect 488644 639976 488783 639978
rect 488644 639920 488722 639976
rect 488778 639920 488783 639976
rect 488644 639918 488783 639920
rect 488644 639916 488650 639918
rect 488717 639915 488783 639918
rect 506606 639916 506612 639980
rect 506676 639978 506682 639980
rect 506749 639978 506815 639981
rect 506676 639976 506815 639978
rect 506676 639920 506754 639976
rect 506810 639920 506815 639976
rect 506676 639918 506815 639920
rect 506676 639916 506682 639918
rect 506749 639915 506815 639918
rect 456977 639706 457043 639709
rect 456977 639704 460092 639706
rect 456977 639648 456982 639704
rect 457038 639648 460092 639704
rect 456977 639646 460092 639648
rect 456977 639643 457043 639646
rect 300853 639434 300919 639437
rect 300718 639432 300919 639434
rect 300718 639376 300858 639432
rect 300914 639376 300919 639432
rect 300718 639374 300919 639376
rect 211245 639371 211311 639374
rect 300853 639371 300919 639374
rect 321553 639026 321619 639029
rect 325006 639026 325066 639472
rect 321553 639024 325066 639026
rect 321553 638968 321558 639024
rect 321614 638968 325066 639024
rect 321553 638966 325066 638968
rect 321553 638963 321619 638966
rect 59077 637938 59143 637941
rect 148593 637938 148659 637941
rect 59077 637936 59554 637938
rect 59077 637880 59082 637936
rect 59138 637926 59554 637936
rect 148593 637936 149530 637938
rect 59138 637880 60076 637926
rect 59077 637878 60076 637880
rect 59077 637875 59143 637878
rect 59494 637866 60076 637878
rect 148593 637880 148598 637936
rect 148654 637926 149530 637936
rect 148654 637880 150052 637926
rect 148593 637878 150052 637880
rect 148593 637875 148659 637878
rect 149470 637866 150052 637878
rect 239446 637810 240032 637870
rect 238201 637802 238267 637805
rect 239446 637802 239506 637810
rect 238201 637800 239506 637802
rect 238201 637744 238206 637800
rect 238262 637744 239506 637800
rect 238201 637742 239506 637744
rect 238201 637739 238267 637742
rect 123109 637258 123175 637261
rect 120796 637256 123175 637258
rect 120796 637200 123114 637256
rect 123170 637200 123175 637256
rect 120796 637198 123175 637200
rect 123109 637195 123175 637198
rect 210742 636714 210802 637228
rect 212625 636714 212691 636717
rect 210742 636712 212691 636714
rect 210742 636656 212630 636712
rect 212686 636656 212691 636712
rect 210742 636654 212691 636656
rect 300718 636714 300778 637228
rect 512177 636986 512243 636989
rect 509956 636984 512243 636986
rect 509956 636928 512182 636984
rect 512238 636928 512243 636984
rect 509956 636926 512243 636928
rect 512177 636923 512243 636926
rect 300945 636714 301011 636717
rect 300718 636712 301011 636714
rect 300718 636656 300950 636712
rect 301006 636656 301011 636712
rect 300718 636654 301011 636656
rect 212625 636651 212691 636654
rect 300945 636651 301011 636654
rect 436277 636034 436343 636037
rect 433750 636032 436343 636034
rect 433750 635976 436282 636032
rect 436338 635976 436343 636032
rect 433750 635974 436343 635976
rect 433750 635392 433810 635974
rect 436277 635971 436343 635974
rect 57789 634538 57855 634541
rect 147397 634538 147463 634541
rect 57789 634536 59554 634538
rect 57789 634480 57794 634536
rect 57850 634526 59554 634536
rect 147397 634536 149530 634538
rect 57850 634480 60076 634526
rect 57789 634478 60076 634480
rect 57789 634475 57855 634478
rect 59494 634466 60076 634478
rect 147397 634480 147402 634536
rect 147458 634526 149530 634536
rect 147458 634480 150052 634526
rect 147397 634478 150052 634480
rect 147397 634475 147463 634478
rect 149470 634466 150052 634478
rect 239446 634410 240032 634470
rect 237373 634402 237439 634405
rect 239446 634402 239506 634410
rect 237373 634400 239506 634402
rect 237373 634344 237378 634400
rect 237434 634344 239506 634400
rect 237373 634342 239506 634344
rect 237373 634339 237439 634342
rect 321553 634130 321619 634133
rect 325006 634130 325066 634712
rect 321553 634128 325066 634130
rect 321553 634072 321558 634128
rect 321614 634072 325066 634128
rect 321553 634070 325066 634072
rect 321553 634067 321619 634070
rect 121545 633858 121611 633861
rect 120796 633856 121611 633858
rect 120796 633800 121550 633856
rect 121606 633800 121611 633856
rect 120796 633798 121611 633800
rect 121545 633795 121611 633798
rect 210742 633450 210802 633828
rect 212717 633450 212783 633453
rect 210742 633448 212783 633450
rect 210742 633392 212722 633448
rect 212778 633392 212783 633448
rect 210742 633390 212783 633392
rect 300718 633450 300778 633828
rect 457713 633586 457779 633589
rect 457713 633584 460092 633586
rect 457713 633528 457718 633584
rect 457774 633528 460092 633584
rect 457713 633526 460092 633528
rect 457713 633523 457779 633526
rect 302233 633450 302299 633453
rect 300718 633448 302299 633450
rect 300718 633392 302238 633448
rect 302294 633392 302299 633448
rect 300718 633390 302299 633392
rect 212717 633387 212783 633390
rect 302233 633387 302299 633390
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 57605 631818 57671 631821
rect 146293 631818 146359 631821
rect 57605 631816 59554 631818
rect 57605 631760 57610 631816
rect 57666 631806 59554 631816
rect 146293 631816 149530 631818
rect 57666 631760 60076 631806
rect 57605 631758 60076 631760
rect 57605 631755 57671 631758
rect 59494 631746 60076 631758
rect 146293 631760 146298 631816
rect 146354 631806 149530 631816
rect 146354 631760 150052 631806
rect 146293 631758 150052 631760
rect 146293 631755 146359 631758
rect 149470 631746 150052 631758
rect 239446 631690 240032 631750
rect 237373 631682 237439 631685
rect 239446 631682 239506 631690
rect 237373 631680 239506 631682
rect 237373 631624 237378 631680
rect 237434 631624 239506 631680
rect 237373 631622 239506 631624
rect 237373 631619 237439 631622
rect 121821 631138 121887 631141
rect 120796 631136 121887 631138
rect 120796 631080 121826 631136
rect 121882 631080 121887 631136
rect 120796 631078 121887 631080
rect 121821 631075 121887 631078
rect 210742 630730 210802 631108
rect 211337 630730 211403 630733
rect 210742 630728 211403 630730
rect 210742 630672 211342 630728
rect 211398 630672 211403 630728
rect 210742 630670 211403 630672
rect 300718 630730 300778 631108
rect 433333 630866 433399 630869
rect 512085 630866 512151 630869
rect 433333 630864 433442 630866
rect 433333 630808 433338 630864
rect 433394 630808 433442 630864
rect 433333 630803 433442 630808
rect 509956 630864 512151 630866
rect 509956 630808 512090 630864
rect 512146 630808 512151 630864
rect 509956 630806 512151 630808
rect 512085 630803 512151 630806
rect 580349 630866 580415 630869
rect 583520 630866 584960 630956
rect 580349 630864 584960 630866
rect 580349 630808 580354 630864
rect 580410 630808 584960 630864
rect 580349 630806 584960 630808
rect 580349 630803 580415 630806
rect 301037 630730 301103 630733
rect 300718 630728 301103 630730
rect 300718 630672 301042 630728
rect 301098 630672 301103 630728
rect 300718 630670 301103 630672
rect 211337 630667 211403 630670
rect 301037 630667 301103 630670
rect 433382 630632 433442 630803
rect 583520 630716 584960 630806
rect 321553 629506 321619 629509
rect 325006 629506 325066 629952
rect 321553 629504 325066 629506
rect 321553 629448 321558 629504
rect 321614 629448 325066 629504
rect 321553 629446 325066 629448
rect 321553 629443 321619 629446
rect 58893 628418 58959 628421
rect 146293 628418 146359 628421
rect 58893 628416 59554 628418
rect 58893 628360 58898 628416
rect 58954 628406 59554 628416
rect 146293 628416 149530 628418
rect 58954 628360 60076 628406
rect 58893 628358 60076 628360
rect 58893 628355 58959 628358
rect 59494 628346 60076 628358
rect 146293 628360 146298 628416
rect 146354 628406 149530 628416
rect 146354 628360 150052 628406
rect 146293 628358 150052 628360
rect 146293 628355 146359 628358
rect 149470 628346 150052 628358
rect 239446 628290 240032 628350
rect 238293 628282 238359 628285
rect 239446 628282 239506 628290
rect 238293 628280 239506 628282
rect 238293 628224 238298 628280
rect 238354 628224 239506 628280
rect 238293 628222 239506 628224
rect 238293 628219 238359 628222
rect 121729 627738 121795 627741
rect 120796 627736 121795 627738
rect 120796 627680 121734 627736
rect 121790 627680 121795 627736
rect 120796 627678 121795 627680
rect 121729 627675 121795 627678
rect 210742 627194 210802 627708
rect 212533 627194 212599 627197
rect 210742 627192 212599 627194
rect 210742 627136 212538 627192
rect 212594 627136 212599 627192
rect 210742 627134 212599 627136
rect 300718 627194 300778 627708
rect 457621 627466 457687 627469
rect 457621 627464 460092 627466
rect 457621 627408 457626 627464
rect 457682 627408 460092 627464
rect 457621 627406 460092 627408
rect 457621 627403 457687 627406
rect 302325 627194 302391 627197
rect 300718 627192 302391 627194
rect 300718 627136 302330 627192
rect 302386 627136 302391 627192
rect 300718 627134 302391 627136
rect 212533 627131 212599 627134
rect 302325 627131 302391 627134
rect 436185 626514 436251 626517
rect 433750 626512 436251 626514
rect 433750 626456 436190 626512
rect 436246 626456 436251 626512
rect 433750 626454 436251 626456
rect 433750 625872 433810 626454
rect 436185 626451 436251 626454
rect 58525 625698 58591 625701
rect 147213 625698 147279 625701
rect 58525 625696 59554 625698
rect 58525 625640 58530 625696
rect 58586 625686 59554 625696
rect 147213 625696 149530 625698
rect 58586 625640 60076 625686
rect 58525 625638 60076 625640
rect 58525 625635 58591 625638
rect 59494 625626 60076 625638
rect 147213 625640 147218 625696
rect 147274 625686 149530 625696
rect 147274 625640 150052 625686
rect 147213 625638 150052 625640
rect 147213 625635 147279 625638
rect 149470 625626 150052 625638
rect 239446 625570 240032 625630
rect 237373 625562 237439 625565
rect 239446 625562 239506 625570
rect 237373 625560 239506 625562
rect 237373 625504 237378 625560
rect 237434 625504 239506 625560
rect 237373 625502 239506 625504
rect 237373 625499 237439 625502
rect 321553 625290 321619 625293
rect 321553 625288 325066 625290
rect 321553 625232 321558 625288
rect 321614 625232 325066 625288
rect 321553 625230 325066 625232
rect 321553 625227 321619 625230
rect 325006 625192 325066 625230
rect 123201 625018 123267 625021
rect 120796 625016 123267 625018
rect 120796 624960 123206 625016
rect 123262 624960 123267 625016
rect 120796 624958 123267 624960
rect 123201 624955 123267 624958
rect 210742 624474 210802 624988
rect 211521 624474 211587 624477
rect 210742 624472 211587 624474
rect 210742 624416 211526 624472
rect 211582 624416 211587 624472
rect 210742 624414 211587 624416
rect 300718 624474 300778 624988
rect 301129 624474 301195 624477
rect 300718 624472 301195 624474
rect 300718 624416 301134 624472
rect 301190 624416 301195 624472
rect 300718 624414 301195 624416
rect 211521 624411 211587 624414
rect 301129 624411 301195 624414
rect 511993 624066 512059 624069
rect 509956 624064 512059 624066
rect 509956 624008 511998 624064
rect 512054 624008 512059 624064
rect 509956 624006 512059 624008
rect 511993 624003 512059 624006
rect 58985 622298 59051 622301
rect 148685 622298 148751 622301
rect 58985 622296 59554 622298
rect 58985 622240 58990 622296
rect 59046 622286 59554 622296
rect 148685 622296 149530 622298
rect 59046 622240 60076 622286
rect 58985 622238 60076 622240
rect 58985 622235 59051 622238
rect 59494 622226 60076 622238
rect 148685 622240 148690 622296
rect 148746 622286 149530 622296
rect 148746 622240 150052 622286
rect 148685 622238 150052 622240
rect 148685 622235 148751 622238
rect 149470 622226 150052 622238
rect 239446 622170 240032 622230
rect 237373 622162 237439 622165
rect 239446 622162 239506 622170
rect 237373 622160 239506 622162
rect 237373 622104 237378 622160
rect 237434 622104 239506 622160
rect 237373 622102 239506 622104
rect 237373 622099 237439 622102
rect 436093 621754 436159 621757
rect 433750 621752 436159 621754
rect 433750 621696 436098 621752
rect 436154 621696 436159 621752
rect 433750 621694 436159 621696
rect 121913 621618 121979 621621
rect 120796 621616 121979 621618
rect 120796 621560 121918 621616
rect 121974 621560 121979 621616
rect 120796 621558 121979 621560
rect 121913 621555 121979 621558
rect 210742 621074 210802 621588
rect 211429 621074 211495 621077
rect 210742 621072 211495 621074
rect 210742 621016 211434 621072
rect 211490 621016 211495 621072
rect 210742 621014 211495 621016
rect 300718 621074 300778 621588
rect 433750 621112 433810 621694
rect 436093 621691 436159 621694
rect 457529 621346 457595 621349
rect 457529 621344 460092 621346
rect 457529 621288 457534 621344
rect 457590 621288 460092 621344
rect 457529 621286 460092 621288
rect 457529 621283 457595 621286
rect 302417 621074 302483 621077
rect 300718 621072 302483 621074
rect 300718 621016 302422 621072
rect 302478 621016 302483 621072
rect 300718 621014 302483 621016
rect 211429 621011 211495 621014
rect 302417 621011 302483 621014
rect 321553 619986 321619 619989
rect 325006 619986 325066 620432
rect 321553 619984 325066 619986
rect 321553 619928 321558 619984
rect 321614 619928 325066 619984
rect 321553 619926 325066 619928
rect 321553 619923 321619 619926
rect 59169 619578 59235 619581
rect 147305 619578 147371 619581
rect 238845 619578 238911 619581
rect 59169 619576 59554 619578
rect 59169 619520 59174 619576
rect 59230 619566 59554 619576
rect 147305 619576 149530 619578
rect 59230 619520 60076 619566
rect 59169 619518 60076 619520
rect 59169 619515 59235 619518
rect 59494 619506 60076 619518
rect 147305 619520 147310 619576
rect 147366 619566 149530 619576
rect 238845 619576 239506 619578
rect 147366 619520 150052 619566
rect 147305 619518 150052 619520
rect 147305 619515 147371 619518
rect 149470 619506 150052 619518
rect 238845 619520 238850 619576
rect 238906 619560 239506 619576
rect 238906 619520 240120 619560
rect 238845 619518 240120 619520
rect 238845 619515 238911 619518
rect 239446 619500 240120 619518
rect -960 619020 480 619260
rect 120766 618357 120826 618868
rect 120766 618352 120875 618357
rect 120766 618296 120814 618352
rect 120870 618296 120875 618352
rect 120766 618294 120875 618296
rect 210742 618354 210802 618868
rect 212809 618354 212875 618357
rect 210742 618352 212875 618354
rect 210742 618296 212814 618352
rect 212870 618296 212875 618352
rect 210742 618294 212875 618296
rect 300718 618354 300778 618868
rect 302601 618354 302667 618357
rect 300718 618352 302667 618354
rect 300718 618296 302606 618352
rect 302662 618296 302667 618352
rect 300718 618294 302667 618296
rect 120809 618291 120875 618294
rect 212809 618291 212875 618294
rect 302601 618291 302667 618294
rect 512085 617946 512151 617949
rect 509956 617944 512151 617946
rect 509956 617888 512090 617944
rect 512146 617888 512151 617944
rect 509956 617886 512151 617888
rect 512085 617883 512151 617886
rect 583520 617388 584960 617628
rect 57881 616178 57947 616181
rect 146201 616178 146267 616181
rect 238017 616178 238083 616181
rect 57881 616176 59554 616178
rect 57881 616120 57886 616176
rect 57942 616166 59554 616176
rect 146201 616176 149530 616178
rect 57942 616120 60076 616166
rect 57881 616118 60076 616120
rect 57881 616115 57947 616118
rect 59494 616106 60076 616118
rect 146201 616120 146206 616176
rect 146262 616166 149530 616176
rect 238017 616176 239506 616178
rect 146262 616120 150052 616166
rect 146201 616118 150052 616120
rect 146201 616115 146267 616118
rect 149470 616106 150052 616118
rect 238017 616120 238022 616176
rect 238078 616160 239506 616176
rect 238078 616120 240120 616160
rect 238017 616118 240120 616120
rect 238017 616115 238083 616118
rect 239446 616100 240120 616118
rect 433750 615906 433810 616352
rect 436737 615906 436803 615909
rect 433750 615904 436803 615906
rect 433750 615848 436742 615904
rect 436798 615848 436803 615904
rect 433750 615846 436803 615848
rect 436737 615843 436803 615846
rect 321553 615634 321619 615637
rect 325006 615634 325066 615672
rect 321553 615632 325066 615634
rect 321553 615576 321558 615632
rect 321614 615576 325066 615632
rect 321553 615574 325066 615576
rect 321553 615571 321619 615574
rect 123385 615498 123451 615501
rect 120796 615496 123451 615498
rect 120796 615440 123390 615496
rect 123446 615440 123451 615496
rect 120796 615438 123451 615440
rect 123385 615435 123451 615438
rect 210742 614954 210802 615468
rect 212993 614954 213059 614957
rect 210742 614952 213059 614954
rect 210742 614896 212998 614952
rect 213054 614896 213059 614952
rect 210742 614894 213059 614896
rect 300718 614954 300778 615468
rect 302509 614954 302575 614957
rect 300718 614952 302575 614954
rect 300718 614896 302514 614952
rect 302570 614896 302575 614952
rect 300718 614894 302575 614896
rect 212993 614891 213059 614894
rect 302509 614891 302575 614894
rect 457621 614546 457687 614549
rect 457621 614544 460092 614546
rect 457621 614488 457626 614544
rect 457682 614488 460092 614544
rect 457621 614486 460092 614488
rect 457621 614483 457687 614486
rect 57513 613458 57579 613461
rect 148501 613458 148567 613461
rect 57513 613456 59554 613458
rect 57513 613400 57518 613456
rect 57574 613446 59554 613456
rect 148501 613456 149530 613458
rect 57574 613400 60076 613446
rect 57513 613398 60076 613400
rect 57513 613395 57579 613398
rect 59494 613386 60076 613398
rect 148501 613400 148506 613456
rect 148562 613446 149530 613456
rect 148562 613400 150052 613446
rect 148501 613398 150052 613400
rect 148501 613395 148567 613398
rect 149470 613386 150052 613398
rect 239446 613330 240032 613390
rect 237373 613322 237439 613325
rect 239446 613322 239506 613330
rect 237373 613320 239506 613322
rect 237373 613264 237378 613320
rect 237434 613264 239506 613320
rect 237373 613262 239506 613264
rect 237373 613259 237439 613262
rect 212901 612914 212967 612917
rect 301221 612914 301287 612917
rect 210742 612912 212967 612914
rect 210742 612856 212906 612912
rect 212962 612856 212967 612912
rect 210742 612854 212967 612856
rect 123017 612778 123083 612781
rect 120796 612776 123083 612778
rect 120796 612720 123022 612776
rect 123078 612720 123083 612776
rect 210742 612748 210802 612854
rect 212901 612851 212967 612854
rect 300718 612912 301287 612914
rect 300718 612856 301226 612912
rect 301282 612856 301287 612912
rect 300718 612854 301287 612856
rect 300718 612748 300778 612854
rect 301221 612851 301287 612854
rect 120796 612718 123083 612720
rect 123017 612715 123083 612718
rect 512177 611826 512243 611829
rect 509956 611824 512243 611826
rect 509956 611768 512182 611824
rect 512238 611768 512243 611824
rect 509956 611766 512243 611768
rect 512177 611763 512243 611766
rect 433382 611421 433442 611592
rect 433333 611416 433442 611421
rect 433333 611360 433338 611416
rect 433394 611360 433442 611416
rect 433333 611358 433442 611360
rect 433333 611355 433399 611358
rect 321553 610330 321619 610333
rect 325006 610330 325066 610912
rect 321553 610328 325066 610330
rect 321553 610272 321558 610328
rect 321614 610272 325066 610328
rect 321553 610270 325066 610272
rect 321553 610267 321619 610270
rect 58801 610058 58867 610061
rect 146293 610058 146359 610061
rect 237373 610058 237439 610061
rect 58801 610056 59554 610058
rect 58801 610000 58806 610056
rect 58862 610046 59554 610056
rect 146293 610056 149530 610058
rect 58862 610000 60076 610046
rect 58801 609998 60076 610000
rect 58801 609995 58867 609998
rect 59494 609986 60076 609998
rect 146293 610000 146298 610056
rect 146354 610046 149530 610056
rect 237373 610056 239506 610058
rect 146354 610000 150052 610046
rect 146293 609998 150052 610000
rect 146293 609995 146359 609998
rect 149470 609986 150052 609998
rect 237373 610000 237378 610056
rect 237434 610040 239506 610056
rect 237434 610000 240120 610040
rect 237373 609998 240120 610000
rect 237373 609995 237439 609998
rect 239446 609980 240120 609998
rect 303153 609514 303219 609517
rect 300718 609512 303219 609514
rect 300718 609456 303158 609512
rect 303214 609456 303219 609512
rect 300718 609454 303219 609456
rect 124029 609378 124095 609381
rect 120796 609376 124095 609378
rect 120796 609320 124034 609376
rect 124090 609320 124095 609376
rect 300718 609348 300778 609454
rect 303153 609451 303219 609454
rect 120796 609318 124095 609320
rect 124029 609315 124095 609318
rect 210742 608834 210802 609348
rect 213821 608834 213887 608837
rect 210742 608832 213887 608834
rect 210742 608776 213826 608832
rect 213882 608776 213887 608832
rect 210742 608774 213887 608776
rect 213821 608771 213887 608774
rect 457529 608426 457595 608429
rect 457529 608424 460092 608426
rect 457529 608368 457534 608424
rect 457590 608368 460092 608424
rect 457529 608366 460092 608368
rect 457529 608363 457595 608366
rect 57421 607338 57487 607341
rect 147121 607338 147187 607341
rect 237373 607338 237439 607341
rect 57421 607336 59554 607338
rect 57421 607280 57426 607336
rect 57482 607326 59554 607336
rect 147121 607336 149530 607338
rect 57482 607280 60076 607326
rect 57421 607278 60076 607280
rect 57421 607275 57487 607278
rect 59494 607266 60076 607278
rect 147121 607280 147126 607336
rect 147182 607326 149530 607336
rect 237373 607336 239506 607338
rect 147182 607280 150052 607326
rect 147121 607278 150052 607280
rect 147121 607275 147187 607278
rect 149470 607266 150052 607278
rect 237373 607280 237378 607336
rect 237434 607320 239506 607336
rect 237434 607280 240120 607320
rect 237373 607278 240120 607280
rect 237373 607275 237439 607278
rect 239446 607260 240120 607278
rect 324221 606794 324287 606797
rect 324221 606792 325066 606794
rect 324221 606736 324226 606792
rect 324282 606736 325066 606792
rect 324221 606734 325066 606736
rect 324221 606731 324287 606734
rect 122005 606658 122071 606661
rect 120796 606656 122071 606658
rect 120796 606600 122010 606656
rect 122066 606600 122071 606656
rect 120796 606598 122071 606600
rect 122005 606595 122071 606598
rect 210742 606250 210802 606628
rect 211705 606250 211771 606253
rect 210742 606248 211771 606250
rect -960 605964 480 606204
rect 210742 606192 211710 606248
rect 211766 606192 211771 606248
rect 210742 606190 211771 606192
rect 300718 606250 300778 606628
rect 301313 606250 301379 606253
rect 300718 606248 301379 606250
rect 300718 606192 301318 606248
rect 301374 606192 301379 606248
rect 300718 606190 301379 606192
rect 211705 606187 211771 606190
rect 301313 606187 301379 606190
rect 325006 606152 325066 606734
rect 433750 606386 433810 606832
rect 436134 606386 436140 606388
rect 433750 606326 436140 606386
rect 436134 606324 436140 606326
rect 436204 606324 436210 606388
rect 511993 605706 512059 605709
rect 509956 605704 512059 605706
rect 509956 605648 511998 605704
rect 512054 605648 512059 605704
rect 509956 605646 512059 605648
rect 511993 605643 512059 605646
rect 583520 604060 584960 604300
rect 58617 603938 58683 603941
rect 148225 603938 148291 603941
rect 58617 603936 59554 603938
rect 58617 603880 58622 603936
rect 58678 603926 59554 603936
rect 148225 603936 149530 603938
rect 58678 603880 60076 603926
rect 58617 603878 60076 603880
rect 58617 603875 58683 603878
rect 59494 603866 60076 603878
rect 148225 603880 148230 603936
rect 148286 603926 149530 603936
rect 148286 603880 150052 603926
rect 148225 603878 150052 603880
rect 148225 603875 148291 603878
rect 149470 603866 150052 603878
rect 239446 603810 240032 603870
rect 237373 603802 237439 603805
rect 239446 603802 239506 603810
rect 237373 603800 239506 603802
rect 237373 603744 237378 603800
rect 237434 603744 239506 603800
rect 237373 603742 239506 603744
rect 237373 603739 237439 603742
rect 213085 603394 213151 603397
rect 302693 603394 302759 603397
rect 210742 603392 213151 603394
rect 210742 603336 213090 603392
rect 213146 603336 213151 603392
rect 210742 603334 213151 603336
rect 121085 603258 121151 603261
rect 120796 603256 121151 603258
rect 120796 603200 121090 603256
rect 121146 603200 121151 603256
rect 210742 603228 210802 603334
rect 213085 603331 213151 603334
rect 300718 603392 302759 603394
rect 300718 603336 302698 603392
rect 302754 603336 302759 603392
rect 300718 603334 302759 603336
rect 300718 603228 300778 603334
rect 302693 603331 302759 603334
rect 120796 603198 121151 603200
rect 121085 603195 121151 603198
rect 457437 602306 457503 602309
rect 457437 602304 460092 602306
rect 457437 602248 457442 602304
rect 457498 602248 460092 602304
rect 457437 602246 460092 602248
rect 457437 602243 457503 602246
rect 433382 601765 433442 602072
rect 433382 601760 433491 601765
rect 433382 601704 433430 601760
rect 433486 601704 433491 601760
rect 433382 601702 433491 601704
rect 433425 601699 433491 601702
rect 57329 601218 57395 601221
rect 147305 601218 147371 601221
rect 57329 601216 59554 601218
rect 57329 601160 57334 601216
rect 57390 601206 59554 601216
rect 147305 601216 149530 601218
rect 57390 601160 60076 601206
rect 57329 601158 60076 601160
rect 57329 601155 57395 601158
rect 59494 601146 60076 601158
rect 147305 601160 147310 601216
rect 147366 601206 149530 601216
rect 147366 601160 150052 601206
rect 147305 601158 150052 601160
rect 147305 601155 147371 601158
rect 149470 601146 150052 601158
rect 239446 601090 240032 601150
rect 237373 601082 237439 601085
rect 239446 601082 239506 601090
rect 237373 601080 239506 601082
rect 237373 601024 237378 601080
rect 237434 601024 239506 601080
rect 237373 601022 239506 601024
rect 237373 601019 237439 601022
rect 321553 600810 321619 600813
rect 325006 600810 325066 601392
rect 321553 600808 325066 600810
rect 321553 600752 321558 600808
rect 321614 600752 325066 600808
rect 321553 600750 325066 600752
rect 321553 600747 321619 600750
rect 211613 600674 211679 600677
rect 301405 600674 301471 600677
rect 210742 600672 211679 600674
rect 210742 600616 211618 600672
rect 211674 600616 211679 600672
rect 210742 600614 211679 600616
rect 122097 600538 122163 600541
rect 120796 600536 122163 600538
rect 120796 600480 122102 600536
rect 122158 600480 122163 600536
rect 210742 600508 210802 600614
rect 211613 600611 211679 600614
rect 300718 600672 301471 600674
rect 300718 600616 301410 600672
rect 301466 600616 301471 600672
rect 300718 600614 301471 600616
rect 300718 600508 300778 600614
rect 301405 600611 301471 600614
rect 120796 600478 122163 600480
rect 122097 600475 122163 600478
rect 512269 599586 512335 599589
rect 509956 599584 512335 599586
rect 509956 599528 512274 599584
rect 512330 599528 512335 599584
rect 509956 599526 512335 599528
rect 512269 599523 512335 599526
rect 58433 597818 58499 597821
rect 146293 597818 146359 597821
rect 58433 597816 59554 597818
rect 58433 597760 58438 597816
rect 58494 597806 59554 597816
rect 146293 597816 149530 597818
rect 58494 597760 60076 597806
rect 58433 597758 60076 597760
rect 58433 597755 58499 597758
rect 59494 597746 60076 597758
rect 146293 597760 146298 597816
rect 146354 597806 149530 597816
rect 146354 597760 150052 597806
rect 146293 597758 150052 597760
rect 146293 597755 146359 597758
rect 149470 597746 150052 597758
rect 239446 597690 240032 597750
rect 237373 597682 237439 597685
rect 239446 597682 239506 597690
rect 237373 597680 239506 597682
rect 237373 597624 237378 597680
rect 237434 597624 239506 597680
rect 237373 597622 239506 597624
rect 237373 597619 237439 597622
rect 122189 597138 122255 597141
rect 120796 597136 122255 597138
rect 120796 597080 122194 597136
rect 122250 597080 122255 597136
rect 120796 597078 122255 597080
rect 122189 597075 122255 597078
rect 210742 596730 210802 597108
rect 211797 596730 211863 596733
rect 210742 596728 211863 596730
rect 210742 596672 211802 596728
rect 211858 596672 211863 596728
rect 210742 596670 211863 596672
rect 300718 596730 300778 597108
rect 302969 596730 303035 596733
rect 300718 596728 303035 596730
rect 300718 596672 302974 596728
rect 303030 596672 303035 596728
rect 300718 596670 303035 596672
rect 433750 596730 433810 597312
rect 434805 596730 434871 596733
rect 433750 596728 434871 596730
rect 433750 596672 434810 596728
rect 434866 596672 434871 596728
rect 433750 596670 434871 596672
rect 211797 596667 211863 596670
rect 302969 596667 303035 596670
rect 434805 596667 434871 596670
rect 321553 596458 321619 596461
rect 325006 596458 325066 596632
rect 321553 596456 325066 596458
rect 321553 596400 321558 596456
rect 321614 596400 325066 596456
rect 321553 596398 325066 596400
rect 321553 596395 321619 596398
rect 457437 596186 457503 596189
rect 457437 596184 460092 596186
rect 457437 596128 457442 596184
rect 457498 596128 460092 596184
rect 457437 596126 460092 596128
rect 457437 596123 457503 596126
rect 59169 595098 59235 595101
rect 146937 595098 147003 595101
rect 59169 595096 59554 595098
rect 59169 595040 59174 595096
rect 59230 595086 59554 595096
rect 146937 595096 149530 595098
rect 59230 595040 60076 595086
rect 59169 595038 60076 595040
rect 59169 595035 59235 595038
rect 59494 595026 60076 595038
rect 146937 595040 146942 595096
rect 146998 595086 149530 595096
rect 146998 595040 150052 595086
rect 146937 595038 150052 595040
rect 146937 595035 147003 595038
rect 149470 595026 150052 595038
rect 239446 594970 240032 595030
rect 237373 594962 237439 594965
rect 239446 594962 239506 594970
rect 237373 594960 239506 594962
rect 237373 594904 237378 594960
rect 237434 594904 239506 594960
rect 237373 594902 239506 594904
rect 237373 594899 237439 594902
rect 123293 594418 123359 594421
rect 120796 594416 123359 594418
rect 120796 594360 123298 594416
rect 123354 594360 123359 594416
rect 120796 594358 123359 594360
rect 123293 594355 123359 594358
rect 210742 593874 210802 594388
rect 213269 593874 213335 593877
rect 210742 593872 213335 593874
rect 210742 593816 213274 593872
rect 213330 593816 213335 593872
rect 210742 593814 213335 593816
rect 300718 593874 300778 594388
rect 301497 593874 301563 593877
rect 300718 593872 301563 593874
rect 300718 593816 301502 593872
rect 301558 593816 301563 593872
rect 300718 593814 301563 593816
rect 213269 593811 213335 593814
rect 301497 593811 301563 593814
rect -960 592908 480 593148
rect 513281 592786 513347 592789
rect 509956 592784 513347 592786
rect 509956 592728 513286 592784
rect 513342 592728 513347 592784
rect 509956 592726 513347 592728
rect 513281 592723 513347 592726
rect 433750 592106 433810 592552
rect 436185 592106 436251 592109
rect 433750 592104 436251 592106
rect 433750 592048 436190 592104
rect 436246 592048 436251 592104
rect 433750 592046 436251 592048
rect 436185 592043 436251 592046
rect 57237 591698 57303 591701
rect 146293 591698 146359 591701
rect 57237 591696 59554 591698
rect 57237 591640 57242 591696
rect 57298 591686 59554 591696
rect 146293 591696 149530 591698
rect 57298 591640 60076 591686
rect 57237 591638 60076 591640
rect 57237 591635 57303 591638
rect 59494 591626 60076 591638
rect 146293 591640 146298 591696
rect 146354 591686 149530 591696
rect 146354 591640 150052 591686
rect 146293 591638 150052 591640
rect 146293 591635 146359 591638
rect 149470 591626 150052 591638
rect 239446 591570 240032 591630
rect 237373 591562 237439 591565
rect 239446 591562 239506 591570
rect 237373 591560 239506 591562
rect 237373 591504 237378 591560
rect 237434 591504 239506 591560
rect 237373 591502 239506 591504
rect 237373 591499 237439 591502
rect 321553 591290 321619 591293
rect 325006 591290 325066 591872
rect 321553 591288 325066 591290
rect 321553 591232 321558 591288
rect 321614 591232 325066 591288
rect 321553 591230 325066 591232
rect 321553 591227 321619 591230
rect 123477 591018 123543 591021
rect 120796 591016 123543 591018
rect 120796 590960 123482 591016
rect 123538 590960 123543 591016
rect 120796 590958 123543 590960
rect 123477 590955 123543 590958
rect 210742 590746 210802 590988
rect 213177 590746 213243 590749
rect 210742 590744 213243 590746
rect 210742 590688 213182 590744
rect 213238 590688 213243 590744
rect 210742 590686 213243 590688
rect 300718 590746 300778 590988
rect 583520 590868 584960 591108
rect 302877 590746 302943 590749
rect 300718 590744 302943 590746
rect 300718 590688 302882 590744
rect 302938 590688 302943 590744
rect 300718 590686 302943 590688
rect 213177 590683 213243 590686
rect 302877 590683 302943 590686
rect 58709 588978 58775 588981
rect 147029 588978 147095 588981
rect 58709 588976 59554 588978
rect 58709 588920 58714 588976
rect 58770 588966 59554 588976
rect 147029 588976 149530 588978
rect 58770 588920 60076 588966
rect 58709 588918 60076 588920
rect 58709 588915 58775 588918
rect 59494 588906 60076 588918
rect 147029 588920 147034 588976
rect 147090 588966 149530 588976
rect 147090 588920 150052 588966
rect 147029 588918 150052 588920
rect 147029 588915 147095 588918
rect 149470 588906 150052 588918
rect 239446 588850 240032 588910
rect 237373 588842 237439 588845
rect 239446 588842 239506 588850
rect 237373 588840 239506 588842
rect 237373 588784 237378 588840
rect 237434 588784 239506 588840
rect 237373 588782 239506 588784
rect 237373 588779 237439 588782
rect 122281 588298 122347 588301
rect 120796 588296 122347 588298
rect 120796 588240 122286 588296
rect 122342 588240 122347 588296
rect 120796 588238 122347 588240
rect 122281 588235 122347 588238
rect 210742 588026 210802 588268
rect 211889 588026 211955 588029
rect 210742 588024 211955 588026
rect 210742 587968 211894 588024
rect 211950 587968 211955 588024
rect 210742 587966 211955 587968
rect 300718 588026 300778 588268
rect 301589 588026 301655 588029
rect 300718 588024 301655 588026
rect 300718 587968 301594 588024
rect 301650 587968 301655 588024
rect 300718 587966 301655 587968
rect 211889 587963 211955 587966
rect 301589 587963 301655 587966
rect 433566 586805 433626 587112
rect 433517 586800 433626 586805
rect 433517 586744 433522 586800
rect 433578 586744 433626 586800
rect 433517 586742 433626 586744
rect 433517 586739 433583 586742
rect 321093 585850 321159 585853
rect 325006 585850 325066 586432
rect 321093 585848 325066 585850
rect 321093 585792 321098 585848
rect 321154 585792 325066 585848
rect 321093 585790 325066 585792
rect 321093 585787 321159 585790
rect 57145 585578 57211 585581
rect 149053 585578 149119 585581
rect 57145 585576 59554 585578
rect 57145 585520 57150 585576
rect 57206 585566 59554 585576
rect 149053 585576 149530 585578
rect 57206 585520 60076 585566
rect 57145 585518 60076 585520
rect 57145 585515 57211 585518
rect 59494 585506 60076 585518
rect 149053 585520 149058 585576
rect 149114 585566 149530 585576
rect 149114 585520 150052 585566
rect 149053 585518 150052 585520
rect 149053 585515 149119 585518
rect 149470 585506 150052 585518
rect 239446 585450 240032 585510
rect 237373 585442 237439 585445
rect 239446 585442 239506 585450
rect 237373 585440 239506 585442
rect 237373 585384 237378 585440
rect 237434 585384 239506 585440
rect 237373 585382 239506 585384
rect 237373 585379 237439 585382
rect 123109 584898 123175 584901
rect 120796 584896 123175 584898
rect 120796 584840 123114 584896
rect 123170 584840 123175 584896
rect 120796 584838 123175 584840
rect 123109 584835 123175 584838
rect 210742 584357 210802 584868
rect 210742 584352 210851 584357
rect 210742 584296 210790 584352
rect 210846 584296 210851 584352
rect 210742 584294 210851 584296
rect 300718 584354 300778 584868
rect 303061 584354 303127 584357
rect 300718 584352 303127 584354
rect 300718 584296 303066 584352
rect 303122 584296 303127 584352
rect 300718 584294 303127 584296
rect 210785 584291 210851 584294
rect 303061 584291 303127 584294
rect 57053 582858 57119 582861
rect 148961 582858 149027 582861
rect 57053 582856 59554 582858
rect 57053 582800 57058 582856
rect 57114 582846 59554 582856
rect 148961 582856 149530 582858
rect 57114 582800 60076 582846
rect 57053 582798 60076 582800
rect 57053 582795 57119 582798
rect 59494 582786 60076 582798
rect 148961 582800 148966 582856
rect 149022 582846 149530 582856
rect 149022 582800 150052 582846
rect 148961 582798 150052 582800
rect 148961 582795 149027 582798
rect 149470 582786 150052 582798
rect 239446 582730 240032 582790
rect 237373 582722 237439 582725
rect 239446 582722 239506 582730
rect 237373 582720 239506 582722
rect 237373 582664 237378 582720
rect 237434 582664 239506 582720
rect 237373 582662 239506 582664
rect 237373 582659 237439 582662
rect 321001 582314 321067 582317
rect 321001 582312 325066 582314
rect 321001 582256 321006 582312
rect 321062 582256 325066 582312
rect 321001 582254 325066 582256
rect 321001 582251 321067 582254
rect 120766 581637 120826 582148
rect 120717 581632 120826 581637
rect 120717 581576 120722 581632
rect 120778 581576 120826 581632
rect 120717 581574 120826 581576
rect 210742 581634 210802 582148
rect 300718 581637 300778 582148
rect 325006 581672 325066 582254
rect 433750 581770 433810 582352
rect 436277 581770 436343 581773
rect 433750 581768 436343 581770
rect 433750 581712 436282 581768
rect 436338 581712 436343 581768
rect 433750 581710 436343 581712
rect 436277 581707 436343 581710
rect 210877 581634 210943 581637
rect 210742 581632 210943 581634
rect 210742 581576 210882 581632
rect 210938 581576 210943 581632
rect 210742 581574 210943 581576
rect 120717 581571 120783 581574
rect 210877 581571 210943 581574
rect 300669 581632 300778 581637
rect 300669 581576 300674 581632
rect 300730 581576 300778 581632
rect 300669 581574 300778 581576
rect 300669 581571 300735 581574
rect -960 580002 480 580092
rect 3141 580002 3207 580005
rect -960 580000 3207 580002
rect -960 579944 3146 580000
rect 3202 579944 3207 580000
rect -960 579942 3207 579944
rect -960 579852 480 579942
rect 3141 579939 3207 579942
rect 580257 577690 580323 577693
rect 583520 577690 584960 577780
rect 580257 577688 584960 577690
rect 580257 577632 580262 577688
rect 580318 577632 584960 577688
rect 580257 577630 584960 577632
rect 580257 577627 580323 577630
rect 433750 577282 433810 577592
rect 583520 577540 584960 577630
rect 436369 577282 436435 577285
rect 433750 577280 436435 577282
rect 433750 577224 436374 577280
rect 436430 577224 436435 577280
rect 433750 577222 436435 577224
rect 436369 577219 436435 577222
rect 321829 576874 321895 576877
rect 325006 576874 325066 576912
rect 321829 576872 325066 576874
rect 321829 576816 321834 576872
rect 321890 576816 325066 576872
rect 321829 576814 325066 576816
rect 321829 576811 321895 576814
rect 433566 572661 433626 572832
rect 433566 572656 433675 572661
rect 433566 572600 433614 572656
rect 433670 572600 433675 572656
rect 433566 572598 433675 572600
rect 433609 572595 433675 572598
rect 321553 571706 321619 571709
rect 325006 571706 325066 572152
rect 321553 571704 325066 571706
rect 321553 571648 321558 571704
rect 321614 571648 325066 571704
rect 321553 571646 325066 571648
rect 321553 571643 321619 571646
rect 433750 567626 433810 568072
rect 436461 567626 436527 567629
rect 433750 567624 436527 567626
rect 433750 567568 436466 567624
rect 436522 567568 436527 567624
rect 433750 567566 436527 567568
rect 436461 567563 436527 567566
rect 321553 567354 321619 567357
rect 325006 567354 325066 567392
rect 321553 567352 325066 567354
rect 321553 567296 321558 567352
rect 321614 567296 325066 567352
rect 321553 567294 325066 567296
rect 321553 567291 321619 567294
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect 433750 563138 433810 563312
rect 436553 563138 436619 563141
rect 433750 563136 436619 563138
rect 433750 563080 436558 563136
rect 436614 563080 436619 563136
rect 433750 563078 436619 563080
rect 436553 563075 436619 563078
rect 321553 562866 321619 562869
rect 321553 562864 325066 562866
rect 321553 562808 321558 562864
rect 321614 562808 325066 562864
rect 321553 562806 325066 562808
rect 321553 562803 321619 562806
rect 325006 562632 325066 562806
rect 433750 558106 433810 558552
rect 436645 558106 436711 558109
rect 433750 558104 436711 558106
rect 433750 558048 436650 558104
rect 436706 558048 436711 558104
rect 433750 558046 436711 558048
rect 436645 558043 436711 558046
rect 321553 557834 321619 557837
rect 325006 557834 325066 557872
rect 321553 557832 325066 557834
rect 321553 557776 321558 557832
rect 321614 557776 325066 557832
rect 321553 557774 325066 557776
rect 321553 557771 321619 557774
rect 255129 555522 255195 555525
rect 323945 555522 324011 555525
rect 255129 555520 324011 555522
rect 255129 555464 255134 555520
rect 255190 555464 323950 555520
rect 324006 555464 324011 555520
rect 255129 555462 324011 555464
rect 255129 555459 255195 555462
rect 323945 555459 324011 555462
rect 298093 555386 298159 555389
rect 305637 555386 305703 555389
rect 298093 555384 305703 555386
rect 298093 555328 298098 555384
rect 298154 555328 305642 555384
rect 305698 555328 305703 555384
rect 298093 555326 305703 555328
rect 298093 555323 298159 555326
rect 305637 555323 305703 555326
rect 286685 555250 286751 555253
rect 322381 555250 322447 555253
rect 286685 555248 322447 555250
rect 286685 555192 286690 555248
rect 286746 555192 322386 555248
rect 322442 555192 322447 555248
rect 286685 555190 322447 555192
rect 286685 555187 286751 555190
rect 322381 555187 322447 555190
rect 241513 555114 241579 555117
rect 300577 555114 300643 555117
rect 241513 555112 300643 555114
rect 241513 555056 241518 555112
rect 241574 555056 300582 555112
rect 300638 555056 300643 555112
rect 241513 555054 300643 555056
rect 241513 555051 241579 555054
rect 300577 555051 300643 555054
rect 238661 554978 238727 554981
rect 300209 554978 300275 554981
rect 238661 554976 300275 554978
rect 238661 554920 238666 554976
rect 238722 554920 300214 554976
rect 300270 554920 300275 554976
rect 238661 554918 300275 554920
rect 238661 554915 238727 554918
rect 300209 554915 300275 554918
rect 285949 554842 286015 554845
rect 302877 554842 302943 554845
rect 285949 554840 302943 554842
rect 285949 554784 285954 554840
rect 286010 554784 302882 554840
rect 302938 554784 302943 554840
rect 285949 554782 302943 554784
rect 285949 554779 286015 554782
rect 302877 554779 302943 554782
rect -960 553740 480 553980
rect 249425 553890 249491 553893
rect 301957 553890 302023 553893
rect 249425 553888 302023 553890
rect 249425 553832 249430 553888
rect 249486 553832 301962 553888
rect 302018 553832 302023 553888
rect 249425 553830 302023 553832
rect 249425 553827 249491 553830
rect 301957 553827 302023 553830
rect 293125 553754 293191 553757
rect 316953 553754 317019 553757
rect 293125 553752 317019 553754
rect 293125 553696 293130 553752
rect 293186 553696 316958 553752
rect 317014 553696 317019 553752
rect 293125 553694 317019 553696
rect 293125 553691 293191 553694
rect 316953 553691 317019 553694
rect 293769 553618 293835 553621
rect 319805 553618 319871 553621
rect 293769 553616 319871 553618
rect 293769 553560 293774 553616
rect 293830 553560 319810 553616
rect 319866 553560 319871 553616
rect 293769 553558 319871 553560
rect 293769 553555 293835 553558
rect 319805 553555 319871 553558
rect 294505 553482 294571 553485
rect 319621 553482 319687 553485
rect 294505 553480 319687 553482
rect 294505 553424 294510 553480
rect 294566 553424 319626 553480
rect 319682 553424 319687 553480
rect 294505 553422 319687 553424
rect 433750 553482 433810 553792
rect 436093 553482 436159 553485
rect 433750 553480 436159 553482
rect 433750 553424 436098 553480
rect 436154 553424 436159 553480
rect 433750 553422 436159 553424
rect 294505 553419 294571 553422
rect 319621 553419 319687 553422
rect 436093 553419 436159 553422
rect 321553 553346 321619 553349
rect 321553 553344 325066 553346
rect 321553 553288 321558 553344
rect 321614 553288 325066 553344
rect 321553 553286 325066 553288
rect 321553 553283 321619 553286
rect 325006 553112 325066 553286
rect 583520 551020 584960 551260
rect 321645 548994 321711 548997
rect 321645 548992 325066 548994
rect 321645 548936 321650 548992
rect 321706 548936 325066 548992
rect 321645 548934 325066 548936
rect 321645 548931 321711 548934
rect 325006 548352 325066 548934
rect 433750 548450 433810 549032
rect 436829 548450 436895 548453
rect 433750 548448 436895 548450
rect 433750 548392 436834 548448
rect 436890 548392 436895 548448
rect 433750 548390 436895 548392
rect 436829 548387 436895 548390
rect 302233 545458 302299 545461
rect 299828 545456 302299 545458
rect 299828 545400 302238 545456
rect 302294 545400 302299 545456
rect 299828 545398 302299 545400
rect 302233 545395 302299 545398
rect 434897 544914 434963 544917
rect 433750 544912 434963 544914
rect 433750 544856 434902 544912
rect 434958 544856 434963 544912
rect 433750 544854 434963 544856
rect 433750 544272 433810 544854
rect 434897 544851 434963 544854
rect 321553 543690 321619 543693
rect 321553 543688 325066 543690
rect 321553 543632 321558 543688
rect 321614 543632 325066 543688
rect 321553 543630 325066 543632
rect 321553 543627 321619 543630
rect 325006 543592 325066 543630
rect -960 540684 480 540924
rect 321553 539338 321619 539341
rect 321553 539336 325066 539338
rect 321553 539280 321558 539336
rect 321614 539280 325066 539336
rect 321553 539278 325066 539280
rect 321553 539275 321619 539278
rect 325006 538832 325066 539278
rect 433750 538930 433810 539512
rect 434621 538930 434687 538933
rect 433750 538928 434687 538930
rect 433750 538872 434626 538928
rect 434682 538872 434687 538928
rect 433750 538870 434687 538872
rect 434621 538867 434687 538870
rect 583520 537692 584960 537932
rect 433425 534986 433491 534989
rect 433382 534984 433491 534986
rect 433382 534928 433430 534984
rect 433486 534928 433491 534984
rect 433382 534923 433491 534928
rect 433382 534752 433442 534923
rect 300577 534578 300643 534581
rect 436134 534578 436140 534580
rect 300577 534576 436140 534578
rect 300577 534520 300582 534576
rect 300638 534520 436140 534576
rect 300577 534518 436140 534520
rect 300577 534515 300643 534518
rect 436134 534516 436140 534518
rect 436204 534516 436210 534580
rect 301957 532674 302023 532677
rect 429193 532674 429259 532677
rect 301957 532672 429259 532674
rect 301957 532616 301962 532672
rect 302018 532616 429198 532672
rect 429254 532616 429259 532672
rect 301957 532614 429259 532616
rect 301957 532611 302023 532614
rect 429193 532611 429259 532614
rect 322749 532538 322815 532541
rect 360745 532538 360811 532541
rect 322749 532536 360811 532538
rect 322749 532480 322754 532536
rect 322810 532480 360750 532536
rect 360806 532480 360811 532536
rect 322749 532478 360811 532480
rect 322749 532475 322815 532478
rect 360745 532475 360811 532478
rect 323853 532402 323919 532405
rect 342713 532402 342779 532405
rect 323853 532400 342779 532402
rect 323853 532344 323858 532400
rect 323914 532344 342718 532400
rect 342774 532344 342779 532400
rect 323853 532342 342779 532344
rect 323853 532339 323919 532342
rect 342713 532339 342779 532342
rect 302417 530498 302483 530501
rect 299828 530496 302483 530498
rect 299828 530440 302422 530496
rect 302478 530440 302483 530496
rect 299828 530438 302483 530440
rect 302417 530435 302483 530438
rect 370630 529076 370636 529140
rect 370700 529138 370706 529140
rect 397453 529138 397519 529141
rect 370700 529136 397519 529138
rect 370700 529080 397458 529136
rect 397514 529080 397519 529136
rect 370700 529078 397519 529080
rect 370700 529076 370706 529078
rect 397453 529075 397519 529078
rect -960 527764 480 528004
rect 371734 526356 371740 526420
rect 371804 526418 371810 526420
rect 512085 526418 512151 526421
rect 371804 526416 512151 526418
rect 371804 526360 512090 526416
rect 512146 526360 512151 526416
rect 371804 526358 512151 526360
rect 371804 526356 371810 526358
rect 512085 526355 512151 526358
rect 583520 524364 584960 524604
rect 57697 523018 57763 523021
rect 57881 523018 57947 523021
rect 57697 523016 60076 523018
rect 57697 522960 57702 523016
rect 57758 522960 57886 523016
rect 57942 522960 60076 523016
rect 57697 522958 60076 522960
rect 57697 522955 57763 522958
rect 57881 522955 57947 522958
rect 302785 515538 302851 515541
rect 299828 515536 302851 515538
rect 299828 515480 302790 515536
rect 302846 515480 302851 515536
rect 299828 515478 302851 515480
rect 302785 515475 302851 515478
rect -960 514858 480 514948
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 578877 511322 578943 511325
rect 583520 511322 584960 511412
rect 578877 511320 584960 511322
rect 578877 511264 578882 511320
rect 578938 511264 584960 511320
rect 578877 511262 584960 511264
rect 578877 511259 578943 511262
rect 583520 511172 584960 511262
rect -960 501652 480 501892
rect 302877 500578 302943 500581
rect 299828 500576 302943 500578
rect 299828 500520 302882 500576
rect 302938 500520 302943 500576
rect 299828 500518 302943 500520
rect 302877 500515 302943 500518
rect 583520 497844 584960 498084
rect 363454 496028 363460 496092
rect 363524 496090 363530 496092
rect 476062 496090 476068 496092
rect 363524 496030 476068 496090
rect 363524 496028 363530 496030
rect 476062 496028 476068 496030
rect 476132 496028 476138 496092
rect 364926 493308 364932 493372
rect 364996 493370 365002 493372
rect 483013 493370 483079 493373
rect 364996 493368 483079 493370
rect 364996 493312 483018 493368
rect 483074 493312 483079 493368
rect 364996 493310 483079 493312
rect 364996 493308 365002 493310
rect 483013 493307 483079 493310
rect 208894 491812 208900 491876
rect 208964 491874 208970 491876
rect 488574 491874 488580 491876
rect 208964 491814 488580 491874
rect 208964 491812 208970 491814
rect 488574 491812 488580 491814
rect 488644 491812 488650 491876
rect 60222 491132 60228 491196
rect 60292 491194 60298 491196
rect 71589 491194 71655 491197
rect 60292 491192 71655 491194
rect 60292 491136 71594 491192
rect 71650 491136 71655 491192
rect 60292 491134 71655 491136
rect 60292 491132 60298 491134
rect 71589 491131 71655 491134
rect 71773 491194 71839 491197
rect 77753 491194 77819 491197
rect 71773 491192 77819 491194
rect 71773 491136 71778 491192
rect 71834 491136 77758 491192
rect 77814 491136 77819 491192
rect 71773 491134 77819 491136
rect 71773 491131 71839 491134
rect 77753 491131 77819 491134
rect 185669 491194 185735 491197
rect 198222 491194 198228 491196
rect 185669 491192 198228 491194
rect 185669 491136 185674 491192
rect 185730 491136 198228 491192
rect 185669 491134 198228 491136
rect 185669 491131 185735 491134
rect 198222 491132 198228 491134
rect 198292 491132 198298 491196
rect 213361 491194 213427 491197
rect 216622 491194 216628 491196
rect 213361 491192 216628 491194
rect 213361 491136 213366 491192
rect 213422 491136 216628 491192
rect 213361 491134 216628 491136
rect 213361 491131 213427 491134
rect 216622 491132 216628 491134
rect 216692 491132 216698 491196
rect 219934 491132 219940 491196
rect 220004 491194 220010 491196
rect 224861 491194 224927 491197
rect 220004 491192 224927 491194
rect 220004 491136 224866 491192
rect 224922 491136 224927 491192
rect 220004 491134 224927 491136
rect 220004 491132 220010 491134
rect 224861 491131 224927 491134
rect 234981 491194 235047 491197
rect 357934 491194 357940 491196
rect 234981 491192 357940 491194
rect 234981 491136 234986 491192
rect 235042 491136 357940 491192
rect 234981 491134 357940 491136
rect 234981 491131 235047 491134
rect 357934 491132 357940 491134
rect 358004 491132 358010 491196
rect 72233 491058 72299 491061
rect 77293 491058 77359 491061
rect 72233 491056 77359 491058
rect 72233 491000 72238 491056
rect 72294 491000 77298 491056
rect 77354 491000 77359 491056
rect 72233 490998 77359 491000
rect 72233 490995 72299 490998
rect 77293 490995 77359 490998
rect 184749 491058 184815 491061
rect 199326 491058 199332 491060
rect 184749 491056 199332 491058
rect 184749 491000 184754 491056
rect 184810 491000 199332 491056
rect 184749 490998 199332 491000
rect 184749 490995 184815 490998
rect 199326 490996 199332 490998
rect 199396 490996 199402 491060
rect 201585 491058 201651 491061
rect 202638 491058 202644 491060
rect 201585 491056 202644 491058
rect 201585 491000 201590 491056
rect 201646 491000 202644 491056
rect 201585 490998 202644 491000
rect 201585 490995 201651 490998
rect 202638 490996 202644 490998
rect 202708 490996 202714 491060
rect 205633 491058 205699 491061
rect 206686 491058 206692 491060
rect 205633 491056 206692 491058
rect 205633 491000 205638 491056
rect 205694 491000 206692 491056
rect 205633 490998 206692 491000
rect 205633 490995 205699 490998
rect 206686 490996 206692 490998
rect 206756 490996 206762 491060
rect 212073 491058 212139 491061
rect 216806 491058 216812 491060
rect 212073 491056 216812 491058
rect 212073 491000 212078 491056
rect 212134 491000 216812 491056
rect 212073 490998 216812 491000
rect 212073 490995 212139 490998
rect 216806 490996 216812 490998
rect 216876 490996 216882 491060
rect 236269 491058 236335 491061
rect 371918 491058 371924 491060
rect 236269 491056 371924 491058
rect 236269 491000 236274 491056
rect 236330 491000 371924 491056
rect 236269 490998 371924 491000
rect 236269 490995 236335 490998
rect 371918 490996 371924 490998
rect 371988 490996 371994 491060
rect 54886 490860 54892 490924
rect 54956 490922 54962 490924
rect 72049 490922 72115 490925
rect 54956 490920 72115 490922
rect 54956 490864 72054 490920
rect 72110 490864 72115 490920
rect 54956 490862 72115 490864
rect 54956 490860 54962 490862
rect 72049 490859 72115 490862
rect 179965 490922 180031 490925
rect 196566 490922 196572 490924
rect 179965 490920 196572 490922
rect 179965 490864 179970 490920
rect 180026 490864 196572 490920
rect 179965 490862 196572 490864
rect 179965 490859 180031 490862
rect 196566 490860 196572 490862
rect 196636 490860 196642 490924
rect 200757 490922 200823 490925
rect 201350 490922 201356 490924
rect 200757 490920 201356 490922
rect 200757 490864 200762 490920
rect 200818 490864 201356 490920
rect 200757 490862 201356 490864
rect 200757 490859 200823 490862
rect 201350 490860 201356 490862
rect 201420 490860 201426 490924
rect 204253 490922 204319 490925
rect 205214 490922 205220 490924
rect 204253 490920 205220 490922
rect 204253 490864 204258 490920
rect 204314 490864 205220 490920
rect 204253 490862 205220 490864
rect 204253 490859 204319 490862
rect 205214 490860 205220 490862
rect 205284 490860 205290 490924
rect 231485 490922 231551 490925
rect 367870 490922 367876 490924
rect 231485 490920 367876 490922
rect 231485 490864 231490 490920
rect 231546 490864 367876 490920
rect 231485 490862 367876 490864
rect 231485 490859 231551 490862
rect 367870 490860 367876 490862
rect 367940 490860 367946 490924
rect 55070 490724 55076 490788
rect 55140 490786 55146 490788
rect 73797 490786 73863 490789
rect 55140 490784 73863 490786
rect 55140 490728 73802 490784
rect 73858 490728 73863 490784
rect 55140 490726 73863 490728
rect 55140 490724 55146 490726
rect 73797 490723 73863 490726
rect 147765 490786 147831 490789
rect 197854 490786 197860 490788
rect 147765 490784 197860 490786
rect 147765 490728 147770 490784
rect 147826 490728 197860 490784
rect 147765 490726 197860 490728
rect 147765 490723 147831 490726
rect 197854 490724 197860 490726
rect 197924 490724 197930 490788
rect 219014 490724 219020 490788
rect 219084 490786 219090 490788
rect 226149 490786 226215 490789
rect 219084 490784 226215 490786
rect 219084 490728 226154 490784
rect 226210 490728 226215 490784
rect 219084 490726 226215 490728
rect 219084 490724 219090 490726
rect 226149 490723 226215 490726
rect 230565 490786 230631 490789
rect 367686 490786 367692 490788
rect 230565 490784 367692 490786
rect 230565 490728 230570 490784
rect 230626 490728 367692 490784
rect 230565 490726 367692 490728
rect 230565 490723 230631 490726
rect 367686 490724 367692 490726
rect 367756 490724 367762 490788
rect 46790 490588 46796 490652
rect 46860 490650 46866 490652
rect 66345 490650 66411 490653
rect 46860 490648 66411 490650
rect 46860 490592 66350 490648
rect 66406 490592 66411 490648
rect 46860 490590 66411 490592
rect 46860 490588 46866 490590
rect 66345 490587 66411 490590
rect 68921 490650 68987 490653
rect 78673 490650 78739 490653
rect 68921 490648 78739 490650
rect 68921 490592 68926 490648
rect 68982 490592 78678 490648
rect 78734 490592 78739 490648
rect 68921 490590 78739 490592
rect 68921 490587 68987 490590
rect 78673 490587 78739 490590
rect 146477 490650 146543 490653
rect 200614 490650 200620 490652
rect 146477 490648 200620 490650
rect 146477 490592 146482 490648
rect 146538 490592 200620 490648
rect 146477 490590 200620 490592
rect 146477 490587 146543 490590
rect 200614 490588 200620 490590
rect 200684 490588 200690 490652
rect 202873 490650 202939 490653
rect 212533 490650 212599 490653
rect 213310 490650 213316 490652
rect 202873 490648 209790 490650
rect 202873 490592 202878 490648
rect 202934 490592 209790 490648
rect 202873 490590 209790 490592
rect 202873 490587 202939 490590
rect 50889 490516 50955 490517
rect 50838 490514 50844 490516
rect 50798 490454 50844 490514
rect 50908 490512 50955 490516
rect 50950 490456 50955 490512
rect 50838 490452 50844 490454
rect 50908 490452 50955 490456
rect 52310 490452 52316 490516
rect 52380 490514 52386 490516
rect 74625 490514 74691 490517
rect 52380 490512 74691 490514
rect 52380 490456 74630 490512
rect 74686 490456 74691 490512
rect 52380 490454 74691 490456
rect 52380 490452 52386 490454
rect 50889 490451 50955 490452
rect 74625 490451 74691 490454
rect 145097 490514 145163 490517
rect 202086 490514 202092 490516
rect 145097 490512 202092 490514
rect 145097 490456 145102 490512
rect 145158 490456 202092 490512
rect 145097 490454 202092 490456
rect 145097 490451 145163 490454
rect 202086 490452 202092 490454
rect 202156 490452 202162 490516
rect 204253 490514 204319 490517
rect 205398 490514 205404 490516
rect 204253 490512 205404 490514
rect 204253 490456 204258 490512
rect 204314 490456 205404 490512
rect 204253 490454 205404 490456
rect 204253 490451 204319 490454
rect 205398 490452 205404 490454
rect 205468 490452 205474 490516
rect 209730 490514 209790 490590
rect 212533 490648 213316 490650
rect 212533 490592 212538 490648
rect 212594 490592 213316 490648
rect 212533 490590 213316 490592
rect 212533 490587 212599 490590
rect 213310 490588 213316 490590
rect 213380 490588 213386 490652
rect 218830 490588 218836 490652
rect 218900 490650 218906 490652
rect 225689 490650 225755 490653
rect 218900 490648 225755 490650
rect 218900 490592 225694 490648
rect 225750 490592 225755 490648
rect 218900 490590 225755 490592
rect 218900 490588 218906 490590
rect 225689 490587 225755 490590
rect 234061 490650 234127 490653
rect 374494 490650 374500 490652
rect 234061 490648 374500 490650
rect 234061 490592 234066 490648
rect 234122 490592 374500 490648
rect 234061 490590 374500 490592
rect 234061 490587 234127 490590
rect 374494 490588 374500 490590
rect 374564 490588 374570 490652
rect 217542 490514 217548 490516
rect 209730 490454 217548 490514
rect 217542 490452 217548 490454
rect 217612 490452 217618 490516
rect 219198 490452 219204 490516
rect 219268 490514 219274 490516
rect 226609 490514 226675 490517
rect 219268 490512 226675 490514
rect 219268 490456 226614 490512
rect 226670 490456 226675 490512
rect 219268 490454 226675 490456
rect 219268 490452 219274 490454
rect 226609 490451 226675 490454
rect 232313 490514 232379 490517
rect 375966 490514 375972 490516
rect 232313 490512 375972 490514
rect 232313 490456 232318 490512
rect 232374 490456 375972 490512
rect 232313 490454 375972 490456
rect 232313 490451 232379 490454
rect 375966 490452 375972 490454
rect 376036 490452 376042 490516
rect 59302 490316 59308 490380
rect 59372 490378 59378 490380
rect 68645 490378 68711 490381
rect 59372 490376 68711 490378
rect 59372 490320 68650 490376
rect 68706 490320 68711 490376
rect 59372 490318 68711 490320
rect 59372 490316 59378 490318
rect 68645 490315 68711 490318
rect 186957 490378 187023 490381
rect 198038 490378 198044 490380
rect 186957 490376 198044 490378
rect 186957 490320 186962 490376
rect 187018 490320 198044 490376
rect 186957 490318 198044 490320
rect 186957 490315 187023 490318
rect 198038 490316 198044 490318
rect 198108 490316 198114 490380
rect 200573 490378 200639 490381
rect 200982 490378 200988 490380
rect 200573 490376 200988 490378
rect 200573 490320 200578 490376
rect 200634 490320 200988 490376
rect 200573 490318 200988 490320
rect 200573 490315 200639 490318
rect 200982 490316 200988 490318
rect 201052 490316 201058 490380
rect 205633 490378 205699 490381
rect 206870 490378 206876 490380
rect 205633 490376 206876 490378
rect 205633 490320 205638 490376
rect 205694 490320 206876 490376
rect 205633 490318 206876 490320
rect 205633 490315 205699 490318
rect 206870 490316 206876 490318
rect 206940 490316 206946 490380
rect 208393 490378 208459 490381
rect 209630 490378 209636 490380
rect 208393 490376 209636 490378
rect 208393 490320 208398 490376
rect 208454 490320 209636 490376
rect 208393 490318 209636 490320
rect 208393 490315 208459 490318
rect 209630 490316 209636 490318
rect 209700 490316 209706 490380
rect 59118 490180 59124 490244
rect 59188 490242 59194 490244
rect 73337 490242 73403 490245
rect 59188 490240 73403 490242
rect 59188 490184 73342 490240
rect 73398 490184 73403 490240
rect 59188 490182 73403 490184
rect 59188 490180 59194 490182
rect 73337 490179 73403 490182
rect 197353 490242 197419 490245
rect 198406 490242 198412 490244
rect 197353 490240 198412 490242
rect 197353 490184 197358 490240
rect 197414 490184 198412 490240
rect 197353 490182 198412 490184
rect 197353 490179 197419 490182
rect 198406 490180 198412 490182
rect 198476 490180 198482 490244
rect 55622 490044 55628 490108
rect 55692 490106 55698 490108
rect 56317 490106 56383 490109
rect 55692 490104 56383 490106
rect 55692 490048 56322 490104
rect 56378 490048 56383 490104
rect 55692 490046 56383 490048
rect 55692 490044 55698 490046
rect 56317 490043 56383 490046
rect 149145 489154 149211 489157
rect 213126 489154 213132 489156
rect 149145 489152 213132 489154
rect 149145 489096 149150 489152
rect 149206 489096 213132 489152
rect 149145 489094 213132 489096
rect 149145 489091 149211 489094
rect 213126 489092 213132 489094
rect 213196 489092 213202 489156
rect 247309 489154 247375 489157
rect 378910 489154 378916 489156
rect 247309 489152 378916 489154
rect 247309 489096 247314 489152
rect 247370 489096 378916 489152
rect 247309 489094 378916 489096
rect 247309 489091 247375 489094
rect 378910 489092 378916 489094
rect 378980 489092 378986 489156
rect -960 488596 480 488836
rect 57094 488276 57100 488340
rect 57164 488338 57170 488340
rect 121361 488338 121427 488341
rect 57164 488336 121427 488338
rect 57164 488280 121366 488336
rect 121422 488280 121427 488336
rect 57164 488278 121427 488280
rect 57164 488276 57170 488278
rect 121361 488275 121427 488278
rect 49141 488202 49207 488205
rect 120441 488202 120507 488205
rect 49141 488200 120507 488202
rect 49141 488144 49146 488200
rect 49202 488144 120446 488200
rect 120502 488144 120507 488200
rect 49141 488142 120507 488144
rect 49141 488139 49207 488142
rect 120441 488139 120507 488142
rect 46657 488066 46723 488069
rect 120073 488066 120139 488069
rect 46657 488064 120139 488066
rect 46657 488008 46662 488064
rect 46718 488008 120078 488064
rect 120134 488008 120139 488064
rect 46657 488006 120139 488008
rect 46657 488003 46723 488006
rect 120073 488003 120139 488006
rect 46473 487930 46539 487933
rect 120901 487930 120967 487933
rect 46473 487928 120967 487930
rect 46473 487872 46478 487928
rect 46534 487872 120906 487928
rect 120962 487872 120967 487928
rect 46473 487870 120967 487872
rect 46473 487867 46539 487870
rect 120901 487867 120967 487870
rect 44030 487732 44036 487796
rect 44100 487794 44106 487796
rect 126605 487794 126671 487797
rect 44100 487792 126671 487794
rect 44100 487736 126610 487792
rect 126666 487736 126671 487792
rect 44100 487734 126671 487736
rect 44100 487732 44106 487734
rect 126605 487731 126671 487734
rect 228817 487794 228883 487797
rect 358118 487794 358124 487796
rect 228817 487792 358124 487794
rect 228817 487736 228822 487792
rect 228878 487736 358124 487792
rect 228817 487734 358124 487736
rect 228817 487731 228883 487734
rect 358118 487732 358124 487734
rect 358188 487732 358194 487796
rect 229277 486434 229343 486437
rect 378726 486434 378732 486436
rect 229277 486432 378732 486434
rect 229277 486376 229282 486432
rect 229338 486376 378732 486432
rect 229277 486374 378732 486376
rect 229277 486371 229343 486374
rect 378726 486372 378732 486374
rect 378796 486372 378802 486436
rect 41321 485618 41387 485621
rect 80789 485618 80855 485621
rect 41321 485616 80855 485618
rect 41321 485560 41326 485616
rect 41382 485560 80794 485616
rect 80850 485560 80855 485616
rect 41321 485558 80855 485560
rect 41321 485555 41387 485558
rect 80789 485555 80855 485558
rect 54753 485482 54819 485485
rect 117405 485482 117471 485485
rect 54753 485480 117471 485482
rect 54753 485424 54758 485480
rect 54814 485424 117410 485480
rect 117466 485424 117471 485480
rect 54753 485422 117471 485424
rect 54753 485419 54819 485422
rect 117405 485419 117471 485422
rect 48129 485346 48195 485349
rect 116485 485346 116551 485349
rect 48129 485344 116551 485346
rect 48129 485288 48134 485344
rect 48190 485288 116490 485344
rect 116546 485288 116551 485344
rect 48129 485286 116551 485288
rect 48129 485283 48195 485286
rect 116485 485283 116551 485286
rect 46565 485210 46631 485213
rect 118693 485210 118759 485213
rect 46565 485208 118759 485210
rect 46565 485152 46570 485208
rect 46626 485152 118698 485208
rect 118754 485152 118759 485208
rect 46565 485150 118759 485152
rect 46565 485147 46631 485150
rect 118693 485147 118759 485150
rect 43989 485074 44055 485077
rect 118233 485074 118299 485077
rect 43989 485072 118299 485074
rect 43989 485016 43994 485072
rect 44050 485016 118238 485072
rect 118294 485016 118299 485072
rect 43989 485014 118299 485016
rect 43989 485011 44055 485014
rect 118233 485011 118299 485014
rect 152641 485074 152707 485077
rect 209814 485074 209820 485076
rect 152641 485072 209820 485074
rect 152641 485016 152646 485072
rect 152702 485016 209820 485072
rect 152641 485014 209820 485016
rect 152641 485011 152707 485014
rect 209814 485012 209820 485014
rect 209884 485012 209890 485076
rect 229737 485074 229803 485077
rect 376150 485074 376156 485076
rect 229737 485072 376156 485074
rect 229737 485016 229742 485072
rect 229798 485016 376156 485072
rect 229737 485014 376156 485016
rect 229737 485011 229803 485014
rect 376150 485012 376156 485014
rect 376220 485012 376226 485076
rect 583520 484516 584960 484756
rect 158805 483850 158871 483853
rect 207974 483850 207980 483852
rect 158805 483848 207980 483850
rect 158805 483792 158810 483848
rect 158866 483792 207980 483848
rect 158805 483790 207980 483792
rect 158805 483787 158871 483790
rect 207974 483788 207980 483790
rect 208044 483788 208050 483852
rect 151261 483714 151327 483717
rect 211654 483714 211660 483716
rect 151261 483712 211660 483714
rect 151261 483656 151266 483712
rect 151322 483656 211660 483712
rect 151261 483654 211660 483656
rect 151261 483651 151327 483654
rect 211654 483652 211660 483654
rect 211724 483652 211730 483716
rect 228357 483714 228423 483717
rect 360694 483714 360700 483716
rect 228357 483712 360700 483714
rect 228357 483656 228362 483712
rect 228418 483656 360700 483712
rect 228357 483654 360700 483656
rect 228357 483651 228423 483654
rect 360694 483652 360700 483654
rect 360764 483652 360770 483716
rect 57462 482428 57468 482492
rect 57532 482490 57538 482492
rect 128445 482490 128511 482493
rect 57532 482488 128511 482490
rect 57532 482432 128450 482488
rect 128506 482432 128511 482488
rect 57532 482430 128511 482432
rect 57532 482428 57538 482430
rect 128445 482427 128511 482430
rect 155677 482490 155743 482493
rect 211838 482490 211844 482492
rect 155677 482488 211844 482490
rect 155677 482432 155682 482488
rect 155738 482432 211844 482488
rect 155677 482430 211844 482432
rect 155677 482427 155743 482430
rect 211838 482428 211844 482430
rect 211908 482428 211914 482492
rect 47710 482292 47716 482356
rect 47780 482354 47786 482356
rect 125317 482354 125383 482357
rect 47780 482352 125383 482354
rect 47780 482296 125322 482352
rect 125378 482296 125383 482352
rect 47780 482294 125383 482296
rect 47780 482292 47786 482294
rect 125317 482291 125383 482294
rect 156137 482354 156203 482357
rect 214046 482354 214052 482356
rect 156137 482352 214052 482354
rect 156137 482296 156142 482352
rect 156198 482296 214052 482352
rect 156137 482294 214052 482296
rect 156137 482291 156203 482294
rect 214046 482292 214052 482294
rect 214116 482292 214122 482356
rect 235441 482354 235507 482357
rect 372654 482354 372660 482356
rect 235441 482352 372660 482354
rect 235441 482296 235446 482352
rect 235502 482296 372660 482352
rect 235441 482294 372660 482296
rect 235441 482291 235507 482294
rect 372654 482292 372660 482294
rect 372724 482292 372730 482356
rect 44950 482156 44956 482220
rect 45020 482218 45026 482220
rect 124029 482218 124095 482221
rect 45020 482216 124095 482218
rect 45020 482160 124034 482216
rect 124090 482160 124095 482216
rect 45020 482158 124095 482160
rect 45020 482156 45026 482158
rect 124029 482155 124095 482158
rect 146937 482218 147003 482221
rect 202270 482218 202276 482220
rect 146937 482216 202276 482218
rect 146937 482160 146942 482216
rect 146998 482160 202276 482216
rect 146937 482158 202276 482160
rect 146937 482155 147003 482158
rect 202270 482156 202276 482158
rect 202340 482156 202346 482220
rect 210366 482156 210372 482220
rect 210436 482218 210442 482220
rect 511993 482218 512059 482221
rect 210436 482216 512059 482218
rect 210436 482160 511998 482216
rect 512054 482160 512059 482216
rect 210436 482158 512059 482160
rect 210436 482156 210442 482158
rect 511993 482155 512059 482158
rect 253473 481130 253539 481133
rect 379462 481130 379468 481132
rect 253473 481128 379468 481130
rect 253473 481072 253478 481128
rect 253534 481072 379468 481128
rect 253473 481070 379468 481072
rect 253473 481067 253539 481070
rect 379462 481068 379468 481070
rect 379532 481068 379538 481132
rect 150433 480994 150499 480997
rect 215886 480994 215892 480996
rect 150433 480992 215892 480994
rect 150433 480936 150438 480992
rect 150494 480936 215892 480992
rect 150433 480934 215892 480936
rect 150433 480931 150499 480934
rect 215886 480932 215892 480934
rect 215956 480932 215962 480996
rect 223941 480994 224007 480997
rect 376334 480994 376340 480996
rect 223941 480992 376340 480994
rect 223941 480936 223946 480992
rect 224002 480936 376340 480992
rect 223941 480934 376340 480936
rect 223941 480931 224007 480934
rect 376334 480932 376340 480934
rect 376404 480932 376410 480996
rect 204846 480796 204852 480860
rect 204916 480858 204922 480860
rect 457529 480858 457595 480861
rect 204916 480856 457595 480858
rect 204916 480800 457534 480856
rect 457590 480800 457595 480856
rect 204916 480798 457595 480800
rect 204916 480796 204922 480798
rect 457529 480795 457595 480798
rect 145557 479498 145623 479501
rect 216070 479498 216076 479500
rect 145557 479496 216076 479498
rect 145557 479440 145562 479496
rect 145618 479440 216076 479496
rect 145557 479438 216076 479440
rect 145557 479435 145623 479438
rect 216070 479436 216076 479438
rect 216140 479436 216146 479500
rect 235901 479498 235967 479501
rect 378174 479498 378180 479500
rect 235901 479496 378180 479498
rect 235901 479440 235906 479496
rect 235962 479440 378180 479496
rect 235901 479438 378180 479440
rect 235901 479435 235967 479438
rect 378174 479436 378180 479438
rect 378244 479436 378250 479500
rect 158345 478138 158411 478141
rect 208342 478138 208348 478140
rect 158345 478136 208348 478138
rect 158345 478080 158350 478136
rect 158406 478080 208348 478136
rect 158345 478078 208348 478080
rect 158345 478075 158411 478078
rect 208342 478076 208348 478078
rect 208412 478076 208418 478140
rect 255681 478138 255747 478141
rect 359406 478138 359412 478140
rect 255681 478136 359412 478138
rect 255681 478080 255686 478136
rect 255742 478080 359412 478136
rect 255681 478078 359412 478080
rect 255681 478075 255747 478078
rect 359406 478076 359412 478078
rect 359476 478076 359482 478140
rect 157057 476914 157123 476917
rect 213862 476914 213868 476916
rect 157057 476912 213868 476914
rect 157057 476856 157062 476912
rect 157118 476856 213868 476912
rect 157057 476854 213868 476856
rect 157057 476851 157123 476854
rect 213862 476852 213868 476854
rect 213932 476852 213938 476916
rect 148685 476778 148751 476781
rect 206134 476778 206140 476780
rect 148685 476776 206140 476778
rect 148685 476720 148690 476776
rect 148746 476720 206140 476776
rect 148685 476718 206140 476720
rect 148685 476715 148751 476718
rect 206134 476716 206140 476718
rect 206204 476716 206210 476780
rect 234521 476778 234587 476781
rect 360142 476778 360148 476780
rect 234521 476776 360148 476778
rect 234521 476720 234526 476776
rect 234582 476720 360148 476776
rect 234521 476718 360148 476720
rect 234521 476715 234587 476718
rect 360142 476716 360148 476718
rect 360212 476716 360218 476780
rect -960 475540 480 475780
rect 252553 475554 252619 475557
rect 377254 475554 377260 475556
rect 252553 475552 377260 475554
rect 252553 475496 252558 475552
rect 252614 475496 377260 475552
rect 252553 475494 377260 475496
rect 252553 475491 252619 475494
rect 377254 475492 377260 475494
rect 377324 475492 377330 475556
rect 153929 475418 153995 475421
rect 215334 475418 215340 475420
rect 153929 475416 215340 475418
rect 153929 475360 153934 475416
rect 153990 475360 215340 475416
rect 153929 475358 215340 475360
rect 153929 475355 153995 475358
rect 215334 475356 215340 475358
rect 215404 475356 215410 475420
rect 231025 475418 231091 475421
rect 372102 475418 372108 475420
rect 231025 475416 372108 475418
rect 231025 475360 231030 475416
rect 231086 475360 372108 475416
rect 231025 475358 372108 475360
rect 231025 475355 231091 475358
rect 372102 475356 372108 475358
rect 372172 475356 372178 475420
rect 165797 474466 165863 474469
rect 216254 474466 216260 474468
rect 165797 474464 216260 474466
rect 165797 474408 165802 474464
rect 165858 474408 216260 474464
rect 165797 474406 216260 474408
rect 165797 474403 165863 474406
rect 216254 474404 216260 474406
rect 216324 474404 216330 474468
rect 146017 474330 146083 474333
rect 203190 474330 203196 474332
rect 146017 474328 203196 474330
rect 146017 474272 146022 474328
rect 146078 474272 203196 474328
rect 146017 474270 203196 474272
rect 146017 474267 146083 474270
rect 203190 474268 203196 474270
rect 203260 474268 203266 474332
rect 151721 474194 151787 474197
rect 214230 474194 214236 474196
rect 151721 474192 214236 474194
rect 151721 474136 151726 474192
rect 151782 474136 214236 474192
rect 151721 474134 214236 474136
rect 151721 474131 151787 474134
rect 214230 474132 214236 474134
rect 214300 474132 214306 474196
rect 122189 474058 122255 474061
rect 196750 474058 196756 474060
rect 122189 474056 196756 474058
rect 122189 474000 122194 474056
rect 122250 474000 196756 474056
rect 122189 473998 196756 474000
rect 122189 473995 122255 473998
rect 196750 473996 196756 473998
rect 196820 473996 196826 474060
rect 230105 474058 230171 474061
rect 370446 474058 370452 474060
rect 230105 474056 370452 474058
rect 230105 474000 230110 474056
rect 230166 474000 370452 474056
rect 230105 473998 370452 474000
rect 230105 473995 230171 473998
rect 370446 473996 370452 473998
rect 370516 473996 370522 474060
rect 366357 472698 366423 472701
rect 506606 472698 506612 472700
rect 366357 472696 506612 472698
rect 366357 472640 366362 472696
rect 366418 472640 506612 472696
rect 366357 472638 506612 472640
rect 366357 472635 366423 472638
rect 506606 472636 506612 472638
rect 506676 472636 506682 472700
rect 172881 472562 172947 472565
rect 202454 472562 202460 472564
rect 172881 472560 202460 472562
rect 172881 472504 172886 472560
rect 172942 472504 202460 472560
rect 172881 472502 202460 472504
rect 172881 472499 172947 472502
rect 202454 472500 202460 472502
rect 202524 472500 202530 472564
rect 233693 472562 233759 472565
rect 378358 472562 378364 472564
rect 233693 472560 378364 472562
rect 233693 472504 233698 472560
rect 233754 472504 378364 472560
rect 233693 472502 378364 472504
rect 233693 472499 233759 472502
rect 378358 472500 378364 472502
rect 378428 472500 378434 472564
rect 173341 471882 173407 471885
rect 203006 471882 203012 471884
rect 173341 471880 203012 471882
rect 173341 471824 173346 471880
rect 173402 471824 203012 471880
rect 173341 471822 203012 471824
rect 173341 471819 173407 471822
rect 203006 471820 203012 471822
rect 203076 471820 203082 471884
rect 44766 471684 44772 471748
rect 44836 471746 44842 471748
rect 65885 471746 65951 471749
rect 44836 471744 65951 471746
rect 44836 471688 65890 471744
rect 65946 471688 65951 471744
rect 44836 471686 65951 471688
rect 44836 471684 44842 471686
rect 65885 471683 65951 471686
rect 172421 471746 172487 471749
rect 205030 471746 205036 471748
rect 172421 471744 205036 471746
rect 172421 471688 172426 471744
rect 172482 471688 205036 471744
rect 172421 471686 205036 471688
rect 172421 471683 172487 471686
rect 205030 471684 205036 471686
rect 205100 471684 205106 471748
rect 57830 471548 57836 471612
rect 57900 471610 57906 471612
rect 91001 471610 91067 471613
rect 57900 471608 91067 471610
rect 57900 471552 91006 471608
rect 91062 471552 91067 471608
rect 57900 471550 91067 471552
rect 57900 471548 57906 471550
rect 91001 471547 91067 471550
rect 182541 471610 182607 471613
rect 217174 471610 217180 471612
rect 182541 471608 217180 471610
rect 182541 471552 182546 471608
rect 182602 471552 217180 471608
rect 182541 471550 217180 471552
rect 182541 471547 182607 471550
rect 217174 471548 217180 471550
rect 217244 471548 217250 471612
rect 59905 471474 59971 471477
rect 92749 471474 92815 471477
rect 59905 471472 92815 471474
rect 59905 471416 59910 471472
rect 59966 471416 92754 471472
rect 92810 471416 92815 471472
rect 59905 471414 92815 471416
rect 59905 471411 59971 471414
rect 92749 471411 92815 471414
rect 162761 471474 162827 471477
rect 202413 471474 202479 471477
rect 162761 471472 202479 471474
rect 162761 471416 162766 471472
rect 162822 471416 202418 471472
rect 202474 471416 202479 471472
rect 162761 471414 202479 471416
rect 162761 471411 162827 471414
rect 202413 471411 202479 471414
rect 295333 471474 295399 471477
rect 359590 471474 359596 471476
rect 295333 471472 359596 471474
rect 295333 471416 295338 471472
rect 295394 471416 359596 471472
rect 295333 471414 359596 471416
rect 295333 471411 295399 471414
rect 359590 471412 359596 471414
rect 359660 471412 359666 471476
rect 56225 471338 56291 471341
rect 90541 471338 90607 471341
rect 56225 471336 90607 471338
rect 56225 471280 56230 471336
rect 56286 471280 90546 471336
rect 90602 471280 90607 471336
rect 56225 471278 90607 471280
rect 56225 471275 56291 471278
rect 90541 471275 90607 471278
rect 160553 471338 160619 471341
rect 202229 471338 202295 471341
rect 160553 471336 202295 471338
rect 160553 471280 160558 471336
rect 160614 471280 202234 471336
rect 202290 471280 202295 471336
rect 160553 471278 202295 471280
rect 160553 471275 160619 471278
rect 202229 471275 202295 471278
rect 297541 471338 297607 471341
rect 377438 471338 377444 471340
rect 297541 471336 377444 471338
rect 297541 471280 297546 471336
rect 297602 471280 377444 471336
rect 297541 471278 377444 471280
rect 297541 471275 297607 471278
rect 377438 471276 377444 471278
rect 377508 471276 377514 471340
rect 583520 471324 584960 471564
rect 47894 471140 47900 471204
rect 47964 471202 47970 471204
rect 82629 471202 82695 471205
rect 47964 471200 82695 471202
rect 47964 471144 82634 471200
rect 82690 471144 82695 471200
rect 47964 471142 82695 471144
rect 47964 471140 47970 471142
rect 82629 471139 82695 471142
rect 163589 471202 163655 471205
rect 209221 471202 209287 471205
rect 163589 471200 209287 471202
rect 163589 471144 163594 471200
rect 163650 471144 209226 471200
rect 209282 471144 209287 471200
rect 163589 471142 209287 471144
rect 163589 471139 163655 471142
rect 209221 471139 209287 471142
rect 296161 471202 296227 471205
rect 377622 471202 377628 471204
rect 296161 471200 377628 471202
rect 296161 471144 296166 471200
rect 296222 471144 377628 471200
rect 296161 471142 377628 471144
rect 296161 471139 296227 471142
rect 377622 471140 377628 471142
rect 377692 471140 377698 471204
rect 58934 469780 58940 469844
rect 59004 469842 59010 469844
rect 69841 469842 69907 469845
rect 59004 469840 69907 469842
rect 59004 469784 69846 469840
rect 69902 469784 69907 469840
rect 59004 469782 69907 469784
rect 59004 469780 59010 469782
rect 69841 469779 69907 469782
rect 181253 469026 181319 469029
rect 199510 469026 199516 469028
rect 181253 469024 199516 469026
rect 181253 468968 181258 469024
rect 181314 468968 199516 469024
rect 181253 468966 199516 468968
rect 181253 468963 181319 468966
rect 199510 468964 199516 468966
rect 199580 468964 199586 469028
rect 48078 468828 48084 468892
rect 48148 468890 48154 468892
rect 70669 468890 70735 468893
rect 48148 468888 70735 468890
rect 48148 468832 70674 468888
rect 70730 468832 70735 468888
rect 48148 468830 70735 468832
rect 48148 468828 48154 468830
rect 70669 468827 70735 468830
rect 161841 468890 161907 468893
rect 200798 468890 200804 468892
rect 161841 468888 200804 468890
rect 161841 468832 161846 468888
rect 161902 468832 200804 468888
rect 161841 468830 200804 468832
rect 161841 468827 161907 468830
rect 200798 468828 200804 468830
rect 200868 468828 200874 468892
rect 46606 468692 46612 468756
rect 46676 468754 46682 468756
rect 70301 468754 70367 468757
rect 46676 468752 70367 468754
rect 46676 468696 70306 468752
rect 70362 468696 70367 468752
rect 46676 468694 70367 468696
rect 46676 468692 46682 468694
rect 70301 468691 70367 468694
rect 169845 468754 169911 468757
rect 210550 468754 210556 468756
rect 169845 468752 210556 468754
rect 169845 468696 169850 468752
rect 169906 468696 210556 468752
rect 169845 468694 210556 468696
rect 169845 468691 169911 468694
rect 210550 468692 210556 468694
rect 210620 468692 210626 468756
rect 53598 468556 53604 468620
rect 53668 468618 53674 468620
rect 79961 468618 80027 468621
rect 53668 468616 80027 468618
rect 53668 468560 79966 468616
rect 80022 468560 80027 468616
rect 53668 468558 80027 468560
rect 53668 468556 53674 468558
rect 79961 468555 80027 468558
rect 154849 468618 154915 468621
rect 218973 468618 219039 468621
rect 154849 468616 219039 468618
rect 154849 468560 154854 468616
rect 154910 468560 218978 468616
rect 219034 468560 219039 468616
rect 154849 468558 219039 468560
rect 154849 468555 154915 468558
rect 218973 468555 219039 468558
rect 50654 468420 50660 468484
rect 50724 468482 50730 468484
rect 80421 468482 80487 468485
rect 50724 468480 80487 468482
rect 50724 468424 80426 468480
rect 80482 468424 80487 468480
rect 50724 468422 80487 468424
rect 50724 468420 50730 468422
rect 80421 468419 80487 468422
rect 147305 468482 147371 468485
rect 218789 468482 218855 468485
rect 147305 468480 218855 468482
rect 147305 468424 147310 468480
rect 147366 468424 218794 468480
rect 218850 468424 218855 468480
rect 147305 468422 218855 468424
rect 147305 468419 147371 468422
rect 218789 468419 218855 468422
rect 276381 468482 276447 468485
rect 359774 468482 359780 468484
rect 276381 468480 359780 468482
rect 276381 468424 276386 468480
rect 276442 468424 359780 468480
rect 276381 468422 359780 468424
rect 276381 468419 276447 468422
rect 359774 468420 359780 468422
rect 359844 468420 359850 468484
rect 58750 467060 58756 467124
rect 58820 467122 58826 467124
rect 68093 467122 68159 467125
rect 58820 467120 68159 467122
rect 58820 467064 68098 467120
rect 68154 467064 68159 467120
rect 58820 467062 68159 467064
rect 58820 467060 58826 467062
rect 68093 467059 68159 467062
rect 171133 467122 171199 467125
rect 206318 467122 206324 467124
rect 171133 467120 206324 467122
rect 171133 467064 171138 467120
rect 171194 467064 206324 467120
rect 171133 467062 206324 467064
rect 171133 467059 171199 467062
rect 206318 467060 206324 467062
rect 206388 467060 206394 467124
rect 178033 466578 178099 466581
rect 178350 466578 178356 466580
rect 178033 466576 178356 466578
rect 178033 466520 178038 466576
rect 178094 466520 178356 466576
rect 178033 466518 178356 466520
rect 178033 466515 178099 466518
rect 178350 466516 178356 466518
rect 178420 466516 178426 466580
rect 179413 466578 179479 466581
rect 190913 466580 190979 466581
rect 338481 466580 338547 466581
rect 339769 466580 339835 466581
rect 350993 466580 351059 466581
rect 179638 466578 179644 466580
rect 179413 466576 179644 466578
rect 179413 466520 179418 466576
rect 179474 466520 179644 466576
rect 179413 466518 179644 466520
rect 179413 466515 179479 466518
rect 179638 466516 179644 466518
rect 179708 466516 179714 466580
rect 190862 466578 190868 466580
rect 190822 466518 190868 466578
rect 190932 466576 190979 466580
rect 338430 466578 338436 466580
rect 190974 466520 190979 466576
rect 190862 466516 190868 466518
rect 190932 466516 190979 466520
rect 338390 466518 338436 466578
rect 338500 466576 338547 466580
rect 339718 466578 339724 466580
rect 338542 466520 338547 466576
rect 338430 466516 338436 466518
rect 338500 466516 338547 466520
rect 339678 466518 339724 466578
rect 339788 466576 339835 466580
rect 350942 466578 350948 466580
rect 339830 466520 339835 466576
rect 339718 466516 339724 466518
rect 339788 466516 339835 466520
rect 350902 466518 350948 466578
rect 351012 466576 351059 466580
rect 351054 466520 351059 466576
rect 350942 466516 350948 466518
rect 351012 466516 351059 466520
rect 190913 466515 190979 466516
rect 338481 466515 338547 466516
rect 339769 466515 339835 466516
rect 350993 466515 351059 466516
rect 498469 466580 498535 466581
rect 499757 466580 499823 466581
rect 510889 466580 510955 466581
rect 498469 466576 498516 466580
rect 498580 466578 498586 466580
rect 498469 466520 498474 466576
rect 498469 466516 498516 466520
rect 498580 466518 498626 466578
rect 499757 466576 499804 466580
rect 499868 466578 499874 466580
rect 510838 466578 510844 466580
rect 499757 466520 499762 466576
rect 498580 466516 498586 466518
rect 499757 466516 499804 466520
rect 499868 466518 499914 466578
rect 510798 466518 510844 466578
rect 510908 466576 510955 466580
rect 510950 466520 510955 466576
rect 499868 466516 499874 466518
rect 510838 466516 510844 466518
rect 510908 466516 510955 466520
rect 498469 466515 498535 466516
rect 499757 466515 499823 466516
rect 510889 466515 510955 466516
rect 53414 466380 53420 466444
rect 53484 466442 53490 466444
rect 75085 466442 75151 466445
rect 53484 466440 75151 466442
rect 53484 466384 75090 466440
rect 75146 466384 75151 466440
rect 53484 466382 75151 466384
rect 53484 466380 53490 466382
rect 75085 466379 75151 466382
rect 54702 466244 54708 466308
rect 54772 466306 54778 466308
rect 76005 466306 76071 466309
rect 54772 466304 76071 466306
rect 54772 466248 76010 466304
rect 76066 466248 76071 466304
rect 54772 466246 76071 466248
rect 54772 466244 54778 466246
rect 76005 466243 76071 466246
rect 53230 466108 53236 466172
rect 53300 466170 53306 466172
rect 76833 466170 76899 466173
rect 53300 466168 76899 466170
rect 53300 466112 76838 466168
rect 76894 466112 76899 466168
rect 53300 466110 76899 466112
rect 53300 466108 53306 466110
rect 76833 466107 76899 466110
rect 180057 466170 180123 466173
rect 198958 466170 198964 466172
rect 180057 466168 198964 466170
rect 180057 466112 180062 466168
rect 180118 466112 198964 466168
rect 180057 466110 198964 466112
rect 180057 466107 180123 466110
rect 198958 466108 198964 466110
rect 199028 466108 199034 466172
rect 51942 465972 51948 466036
rect 52012 466034 52018 466036
rect 76465 466034 76531 466037
rect 52012 466032 76531 466034
rect 52012 465976 76470 466032
rect 76526 465976 76531 466032
rect 52012 465974 76531 465976
rect 52012 465972 52018 465974
rect 76465 465971 76531 465974
rect 167177 466034 167243 466037
rect 208158 466034 208164 466036
rect 167177 466032 208164 466034
rect 167177 465976 167182 466032
rect 167238 465976 208164 466032
rect 167177 465974 208164 465976
rect 167177 465971 167243 465974
rect 208158 465972 208164 465974
rect 208228 465972 208234 466036
rect 52126 465836 52132 465900
rect 52196 465898 52202 465900
rect 78213 465898 78279 465901
rect 52196 465896 78279 465898
rect 52196 465840 78218 465896
rect 78274 465840 78279 465896
rect 52196 465838 78279 465840
rect 52196 465836 52202 465838
rect 78213 465835 78279 465838
rect 168925 465898 168991 465901
rect 219065 465898 219131 465901
rect 168925 465896 219131 465898
rect 168925 465840 168930 465896
rect 168986 465840 219070 465896
rect 219126 465840 219131 465896
rect 168925 465838 219131 465840
rect 168925 465835 168991 465838
rect 219065 465835 219131 465838
rect 298369 465898 298435 465901
rect 377806 465898 377812 465900
rect 298369 465896 377812 465898
rect 298369 465840 298374 465896
rect 298430 465840 377812 465896
rect 298369 465838 377812 465840
rect 298369 465835 298435 465838
rect 377806 465836 377812 465838
rect 377876 465836 377882 465900
rect 48630 465700 48636 465764
rect 48700 465762 48706 465764
rect 79041 465762 79107 465765
rect 48700 465760 79107 465762
rect 48700 465704 79046 465760
rect 79102 465704 79107 465760
rect 48700 465702 79107 465704
rect 48700 465700 48706 465702
rect 79041 465699 79107 465702
rect 107745 465762 107811 465765
rect 198774 465762 198780 465764
rect 107745 465760 198780 465762
rect 107745 465704 107750 465760
rect 107806 465704 198780 465760
rect 107745 465702 198780 465704
rect 107745 465699 107811 465702
rect 198774 465700 198780 465702
rect 198844 465700 198850 465764
rect 224401 465762 224467 465765
rect 373257 465762 373323 465765
rect 224401 465760 373323 465762
rect 224401 465704 224406 465760
rect 224462 465704 373262 465760
rect 373318 465704 373323 465760
rect 224401 465702 373323 465704
rect 224401 465699 224467 465702
rect 373257 465699 373323 465702
rect 58566 465564 58572 465628
rect 58636 465626 58642 465628
rect 69381 465626 69447 465629
rect 58636 465624 69447 465626
rect 58636 465568 69386 465624
rect 69442 465568 69447 465624
rect 58636 465566 69447 465568
rect 58636 465564 58642 465566
rect 69381 465563 69447 465566
rect 50470 465156 50476 465220
rect 50540 465218 50546 465220
rect 50705 465218 50771 465221
rect 50540 465216 50771 465218
rect 50540 465160 50710 465216
rect 50766 465160 50771 465216
rect 50540 465158 50771 465160
rect 50540 465156 50546 465158
rect 50705 465155 50771 465158
rect 57646 464340 57652 464404
rect 57716 464402 57722 464404
rect 92289 464402 92355 464405
rect 57716 464400 92355 464402
rect 57716 464344 92294 464400
rect 92350 464344 92355 464400
rect 57716 464342 92355 464344
rect 57716 464340 57722 464342
rect 92289 464339 92355 464342
rect 183461 464402 183527 464405
rect 205173 464402 205239 464405
rect 183461 464400 205239 464402
rect 183461 464344 183466 464400
rect 183522 464344 205178 464400
rect 205234 464344 205239 464400
rect 183461 464342 205239 464344
rect 183461 464339 183527 464342
rect 205173 464339 205239 464342
rect -960 462634 480 462724
rect 3601 462634 3667 462637
rect -960 462632 3667 462634
rect -960 462576 3606 462632
rect 3662 462576 3667 462632
rect -960 462574 3667 462576
rect -960 462484 480 462574
rect 3601 462571 3667 462574
rect 196558 460186 196618 460190
rect 198733 460186 198799 460189
rect 196558 460184 198799 460186
rect 196558 460128 198738 460184
rect 198794 460128 198799 460184
rect 196558 460126 198799 460128
rect 356562 460186 356622 460190
rect 359365 460186 359431 460189
rect 356562 460184 359431 460186
rect 356562 460128 359370 460184
rect 359426 460128 359431 460184
rect 356562 460126 359431 460128
rect 198733 460123 198799 460126
rect 359365 460123 359431 460126
rect 516558 459642 516618 460190
rect 518893 459642 518959 459645
rect 519445 459642 519511 459645
rect 516558 459640 519511 459642
rect 516558 459584 518898 459640
rect 518954 459584 519450 459640
rect 519506 459584 519511 459640
rect 516558 459582 519511 459584
rect 518893 459579 518959 459582
rect 519445 459579 519511 459582
rect 580257 458146 580323 458149
rect 583520 458146 584960 458236
rect 580257 458144 584960 458146
rect 580257 458088 580262 458144
rect 580318 458088 584960 458144
rect 580257 458086 584960 458088
rect 580257 458083 580323 458086
rect 583520 457996 584960 458086
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect 57789 417890 57855 417893
rect 60002 417890 60062 417894
rect 57789 417888 60062 417890
rect 57789 417832 57794 417888
rect 57850 417832 60062 417888
rect 57789 417830 60062 417832
rect 216765 417890 216831 417893
rect 217777 417890 217843 417893
rect 219390 417890 220064 417924
rect 216765 417888 220064 417890
rect 216765 417832 216770 417888
rect 216826 417832 217782 417888
rect 217838 417864 220064 417888
rect 377029 417890 377095 417893
rect 379470 417890 380052 417924
rect 377029 417888 380052 417890
rect 217838 417832 219450 417864
rect 216765 417830 219450 417832
rect 377029 417832 377034 417888
rect 377090 417864 380052 417888
rect 377090 417832 379530 417864
rect 377029 417830 379530 417832
rect 57789 417827 57855 417830
rect 216765 417827 216831 417830
rect 217777 417827 217843 417830
rect 377029 417827 377095 417830
rect 57237 417618 57303 417621
rect 57237 417616 60062 417618
rect 57237 417560 57242 417616
rect 57298 417560 60062 417616
rect 57237 417558 60062 417560
rect 57237 417555 57303 417558
rect 60002 416942 60062 417558
rect 216857 416938 216923 416941
rect 217869 416938 217935 416941
rect 219390 416938 220064 416972
rect 216857 416936 220064 416938
rect 216857 416880 216862 416936
rect 216918 416880 217874 416936
rect 217930 416912 220064 416936
rect 377765 416938 377831 416941
rect 378041 416938 378107 416941
rect 379470 416938 380052 416972
rect 377765 416936 380052 416938
rect 217930 416880 219450 416912
rect 216857 416878 219450 416880
rect 377765 416880 377770 416936
rect 377826 416880 378046 416936
rect 378102 416912 380052 416936
rect 378102 416880 379530 416912
rect 377765 416878 379530 416880
rect 216857 416875 216923 416878
rect 217869 416875 217935 416878
rect 377765 416875 377831 416878
rect 378041 416875 378107 416878
rect 57789 414218 57855 414221
rect 60002 414218 60062 414766
rect 216857 414762 216923 414765
rect 219390 414762 220064 414796
rect 216857 414760 220064 414762
rect 216857 414704 216862 414760
rect 216918 414736 220064 414760
rect 377765 414762 377831 414765
rect 379470 414762 380052 414796
rect 377765 414760 380052 414762
rect 216918 414704 219450 414736
rect 216857 414702 219450 414704
rect 377765 414704 377770 414760
rect 377826 414736 380052 414760
rect 377826 414704 379530 414736
rect 377765 414702 379530 414704
rect 216857 414699 216923 414702
rect 377765 414699 377831 414702
rect 57789 414216 60062 414218
rect 57789 414160 57794 414216
rect 57850 414160 60062 414216
rect 57789 414158 60062 414160
rect 57789 414155 57855 414158
rect 57789 413266 57855 413269
rect 60002 413266 60062 413814
rect 216673 413810 216739 413813
rect 219390 413810 220064 413844
rect 216673 413808 220064 413810
rect 216673 413752 216678 413808
rect 216734 413784 220064 413808
rect 377673 413810 377739 413813
rect 379470 413810 380052 413844
rect 377673 413808 380052 413810
rect 216734 413752 219450 413784
rect 216673 413750 219450 413752
rect 377673 413752 377678 413808
rect 377734 413784 380052 413808
rect 377734 413752 379530 413784
rect 377673 413750 379530 413752
rect 216673 413747 216739 413750
rect 377673 413747 377739 413750
rect 57789 413264 60062 413266
rect 57789 413208 57794 413264
rect 57850 413208 60062 413264
rect 57789 413206 60062 413208
rect 57789 413203 57855 413206
rect 57789 411498 57855 411501
rect 60002 411498 60062 412046
rect 217685 412042 217751 412045
rect 219390 412042 220064 412076
rect 217685 412040 220064 412042
rect 217685 411984 217690 412040
rect 217746 412016 220064 412040
rect 377029 412042 377095 412045
rect 377489 412042 377555 412045
rect 379470 412042 380052 412076
rect 377029 412040 380052 412042
rect 217746 411984 219450 412016
rect 217685 411982 219450 411984
rect 377029 411984 377034 412040
rect 377090 411984 377494 412040
rect 377550 412016 380052 412040
rect 377550 411984 379530 412016
rect 377029 411982 379530 411984
rect 217685 411979 217751 411982
rect 377029 411979 377095 411982
rect 377489 411979 377555 411982
rect 57789 411496 60062 411498
rect 57789 411440 57794 411496
rect 57850 411440 60062 411496
rect 57789 411438 60062 411440
rect 57789 411435 57855 411438
rect -960 410546 480 410636
rect 2957 410546 3023 410549
rect -960 410544 3023 410546
rect -960 410488 2962 410544
rect 3018 410488 3023 410544
rect -960 410486 3023 410488
rect -960 410396 480 410486
rect 2957 410483 3023 410486
rect 57789 410410 57855 410413
rect 60002 410410 60062 410958
rect 217225 410954 217291 410957
rect 219390 410954 220064 410988
rect 217225 410952 220064 410954
rect 217225 410896 217230 410952
rect 217286 410928 220064 410952
rect 377397 410954 377463 410957
rect 379470 410954 380052 410988
rect 377397 410952 380052 410954
rect 217286 410896 219450 410928
rect 217225 410894 219450 410896
rect 377397 410896 377402 410952
rect 377458 410928 380052 410952
rect 377458 410896 379530 410928
rect 377397 410894 379530 410896
rect 217225 410891 217291 410894
rect 377397 410891 377463 410894
rect 359958 410484 359964 410548
rect 360028 410546 360034 410548
rect 376753 410546 376819 410549
rect 360028 410544 376819 410546
rect 360028 410488 376758 410544
rect 376814 410488 376819 410544
rect 360028 410486 376819 410488
rect 360028 410484 360034 410486
rect 376753 410483 376819 410486
rect 57789 410408 60062 410410
rect 57789 410352 57794 410408
rect 57850 410352 60062 410408
rect 57789 410350 60062 410352
rect 57789 410347 57855 410350
rect 57789 408642 57855 408645
rect 60002 408642 60062 409190
rect 216765 409186 216831 409189
rect 219390 409186 220064 409220
rect 216765 409184 220064 409186
rect 216765 409128 216770 409184
rect 216826 409160 220064 409184
rect 377397 409186 377463 409189
rect 377949 409186 378015 409189
rect 379470 409186 380052 409220
rect 377397 409184 380052 409186
rect 216826 409128 219450 409160
rect 216765 409126 219450 409128
rect 377397 409128 377402 409184
rect 377458 409128 377954 409184
rect 378010 409160 380052 409184
rect 378010 409128 379530 409160
rect 377397 409126 379530 409128
rect 216765 409123 216831 409126
rect 377397 409123 377463 409126
rect 377949 409123 378015 409126
rect 57789 408640 60062 408642
rect 57789 408584 57794 408640
rect 57850 408584 60062 408640
rect 57789 408582 60062 408584
rect 57789 408579 57855 408582
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect 196558 400346 196618 400350
rect 198917 400346 198983 400349
rect 196558 400344 198983 400346
rect 196558 400288 198922 400344
rect 198978 400288 198983 400344
rect 196558 400286 198983 400288
rect 356562 400346 356622 400350
rect 359089 400346 359155 400349
rect 356562 400344 359155 400346
rect 356562 400288 359094 400344
rect 359150 400288 359155 400344
rect 356562 400286 359155 400288
rect 516558 400346 516618 400350
rect 519353 400346 519419 400349
rect 516558 400344 519419 400346
rect 516558 400288 519358 400344
rect 519414 400288 519419 400344
rect 516558 400286 519419 400288
rect 198917 400283 198983 400286
rect 359089 400283 359155 400286
rect 519353 400283 519419 400286
rect 196558 398306 196618 398718
rect 199561 398306 199627 398309
rect 196558 398304 199627 398306
rect 196558 398248 199566 398304
rect 199622 398248 199627 398304
rect 196558 398246 199627 398248
rect 199561 398243 199627 398246
rect 356562 398170 356622 398718
rect 358997 398170 359063 398173
rect 356562 398168 359063 398170
rect 356562 398112 359002 398168
rect 359058 398112 359063 398168
rect 356562 398110 359063 398112
rect 516558 398170 516618 398718
rect 518985 398170 519051 398173
rect 516558 398168 519051 398170
rect 516558 398112 518990 398168
rect 519046 398112 519051 398168
rect 516558 398110 519051 398112
rect 358997 398107 359063 398110
rect 518985 398107 519051 398110
rect -960 397340 480 397580
rect 196558 397354 196618 397358
rect 199193 397354 199259 397357
rect 199469 397354 199535 397357
rect 196558 397352 199535 397354
rect 196558 397296 199198 397352
rect 199254 397296 199474 397352
rect 199530 397296 199535 397352
rect 196558 397294 199535 397296
rect 199193 397291 199259 397294
rect 199469 397291 199535 397294
rect 356562 396810 356622 397358
rect 359733 396810 359799 396813
rect 356562 396808 359799 396810
rect 356562 396752 359738 396808
rect 359794 396752 359799 396808
rect 356562 396750 359799 396752
rect 516558 396810 516618 397358
rect 519169 396810 519235 396813
rect 516558 396808 519235 396810
rect 516558 396752 519174 396808
rect 519230 396752 519235 396808
rect 516558 396750 519235 396752
rect 359733 396747 359799 396750
rect 519169 396747 519235 396750
rect 198641 396674 198707 396677
rect 216806 396674 216812 396676
rect 198641 396672 216812 396674
rect 198641 396616 198646 396672
rect 198702 396616 216812 396672
rect 198641 396614 216812 396616
rect 198641 396611 198707 396614
rect 216806 396612 216812 396614
rect 216876 396612 216882 396676
rect 196558 395314 196618 395862
rect 198917 395314 198983 395317
rect 196558 395312 198983 395314
rect 196558 395256 198922 395312
rect 198978 395256 198983 395312
rect 196558 395254 198983 395256
rect 356562 395314 356622 395862
rect 359917 395314 359983 395317
rect 356562 395312 359983 395314
rect 356562 395256 359922 395312
rect 359978 395256 359983 395312
rect 356562 395254 359983 395256
rect 516558 395314 516618 395862
rect 519077 395314 519143 395317
rect 516558 395312 519143 395314
rect 516558 395256 519082 395312
rect 519138 395256 519143 395312
rect 516558 395254 519143 395256
rect 198917 395251 198983 395254
rect 359917 395251 359983 395254
rect 519077 395251 519143 395254
rect 196558 394634 196618 394638
rect 199837 394634 199903 394637
rect 196558 394632 199903 394634
rect 196558 394576 199842 394632
rect 199898 394576 199903 394632
rect 196558 394574 199903 394576
rect 199837 394571 199903 394574
rect 356562 394090 356622 394638
rect 359825 394090 359891 394093
rect 356562 394088 359891 394090
rect 356562 394032 359830 394088
rect 359886 394032 359891 394088
rect 356562 394030 359891 394032
rect 516558 394090 516618 394638
rect 519261 394090 519327 394093
rect 516558 394088 519327 394090
rect 516558 394032 519266 394088
rect 519322 394032 519327 394088
rect 516558 394030 519327 394032
rect 359825 394027 359891 394030
rect 519261 394027 519327 394030
rect 57697 391642 57763 391645
rect 57697 391640 60062 391642
rect 57697 391584 57702 391640
rect 57758 391584 60062 391640
rect 583520 391628 584960 391868
rect 57697 391582 60062 391584
rect 57697 391579 57763 391582
rect 60002 390966 60062 391582
rect 216949 390962 217015 390965
rect 219390 390962 220064 390996
rect 216949 390960 220064 390962
rect 216949 390904 216954 390960
rect 217010 390936 220064 390960
rect 376845 390962 376911 390965
rect 379470 390962 380052 390996
rect 376845 390960 380052 390962
rect 217010 390904 219450 390936
rect 216949 390902 219450 390904
rect 376845 390904 376850 390960
rect 376906 390936 380052 390960
rect 376906 390904 379530 390936
rect 376845 390902 379530 390904
rect 216949 390899 217015 390902
rect 376845 390899 376911 390902
rect 57462 390628 57468 390692
rect 57532 390690 57538 390692
rect 58341 390690 58407 390693
rect 57532 390688 58407 390690
rect 57532 390632 58346 390688
rect 58402 390632 58407 390688
rect 57532 390630 58407 390632
rect 57532 390628 57538 390630
rect 58341 390627 58407 390630
rect 57421 389330 57487 389333
rect 59494 389330 60032 389364
rect 57421 389328 60032 389330
rect 57421 389272 57426 389328
rect 57482 389304 60032 389328
rect 216673 389330 216739 389333
rect 219390 389330 220064 389364
rect 216673 389328 220064 389330
rect 57482 389272 59554 389304
rect 57421 389270 59554 389272
rect 216673 389272 216678 389328
rect 216734 389304 220064 389328
rect 376937 389330 377003 389333
rect 379470 389330 380052 389364
rect 376937 389328 380052 389330
rect 216734 389272 219450 389304
rect 216673 389270 219450 389272
rect 376937 389272 376942 389328
rect 376998 389304 380052 389328
rect 376998 389272 379530 389304
rect 376937 389270 379530 389272
rect 57421 389267 57487 389270
rect 216673 389267 216739 389270
rect 376937 389267 377003 389270
rect 57237 389058 57303 389061
rect 60002 389058 60062 389062
rect 57237 389056 60062 389058
rect 57237 389000 57242 389056
rect 57298 389000 60062 389056
rect 57237 388998 60062 389000
rect 216949 389058 217015 389061
rect 219390 389058 220064 389092
rect 216949 389056 220064 389058
rect 216949 389000 216954 389056
rect 217010 389032 220064 389056
rect 376937 389058 377003 389061
rect 379470 389058 380052 389092
rect 376937 389056 380052 389058
rect 217010 389000 219450 389032
rect 216949 388998 219450 389000
rect 376937 389000 376942 389056
rect 376998 389032 380052 389056
rect 376998 389000 379530 389032
rect 376937 388998 379530 389000
rect 57237 388995 57303 388998
rect 216949 388995 217015 388998
rect 376937 388995 377003 388998
rect 53230 388452 53236 388516
rect 53300 388514 53306 388516
rect 53741 388514 53807 388517
rect 53300 388512 53807 388514
rect 53300 388456 53746 388512
rect 53802 388456 53807 388512
rect 53300 388454 53807 388456
rect 53300 388452 53306 388454
rect 53741 388451 53807 388454
rect -960 384284 480 384524
rect 55489 381034 55555 381037
rect 55622 381034 55628 381036
rect 55489 381032 55628 381034
rect 55489 380976 55494 381032
rect 55550 380976 55628 381032
rect 55489 380974 55628 380976
rect 55489 380971 55555 380974
rect 55622 380972 55628 380974
rect 55692 380972 55698 381036
rect 198406 380972 198412 381036
rect 198476 381034 198482 381036
rect 198549 381034 198615 381037
rect 198476 381032 198615 381034
rect 198476 380976 198554 381032
rect 198610 380976 198615 381032
rect 198476 380974 198615 380976
rect 198476 380972 198482 380974
rect 198549 380971 198615 380974
rect 200982 380972 200988 381036
rect 201052 381034 201058 381036
rect 201401 381034 201467 381037
rect 201052 381032 201467 381034
rect 201052 380976 201406 381032
rect 201462 380976 201467 381032
rect 201052 380974 201467 380976
rect 201052 380972 201058 380974
rect 201401 380971 201467 380974
rect 413553 380900 413619 380901
rect 421097 380900 421163 380901
rect 425973 380900 426039 380901
rect 433609 380900 433675 380901
rect 84208 380836 84214 380900
rect 84278 380898 84284 380900
rect 323360 380898 323366 380900
rect 84278 380838 209790 380898
rect 84278 380836 84284 380838
rect 83120 380700 83126 380764
rect 83190 380762 83196 380764
rect 207013 380762 207079 380765
rect 83190 380760 207079 380762
rect 83190 380704 207018 380760
rect 207074 380704 207079 380760
rect 83190 380702 207079 380704
rect 209730 380762 209790 380838
rect 219390 380838 323366 380898
rect 211245 380762 211311 380765
rect 213637 380762 213703 380765
rect 209730 380760 213703 380762
rect 209730 380704 211250 380760
rect 211306 380704 213642 380760
rect 213698 380704 213703 380760
rect 209730 380702 213703 380704
rect 83190 380700 83196 380702
rect 207013 380699 207079 380702
rect 211245 380699 211311 380702
rect 213637 380699 213703 380702
rect 217542 380700 217548 380764
rect 217612 380762 217618 380764
rect 219390 380762 219450 380838
rect 323360 380836 323366 380838
rect 323430 380836 323436 380900
rect 413553 380896 413598 380900
rect 413662 380898 413668 380900
rect 421072 380898 421078 380900
rect 413553 380840 413558 380896
rect 413553 380836 413598 380840
rect 413662 380838 413710 380898
rect 421006 380838 421078 380898
rect 421142 380896 421163 380900
rect 425968 380898 425974 380900
rect 421158 380840 421163 380896
rect 413662 380836 413668 380838
rect 421072 380836 421078 380838
rect 421142 380836 421163 380840
rect 425882 380838 425974 380898
rect 425968 380836 425974 380838
rect 426038 380836 426044 380900
rect 433584 380898 433590 380900
rect 433518 380838 433590 380898
rect 433654 380896 433675 380900
rect 433670 380840 433675 380896
rect 433584 380836 433590 380838
rect 433654 380836 433675 380840
rect 413553 380835 413619 380836
rect 421097 380835 421163 380836
rect 425973 380835 426039 380836
rect 433609 380835 433675 380836
rect 436001 380900 436067 380901
rect 436001 380896 436038 380900
rect 436102 380898 436108 380900
rect 436001 380840 436006 380896
rect 436001 380836 436038 380840
rect 436102 380838 436158 380898
rect 436102 380836 436108 380838
rect 436001 380835 436067 380836
rect 217612 380702 219450 380762
rect 235993 380764 236059 380765
rect 237097 380764 237163 380765
rect 243077 380764 243143 380765
rect 248229 380764 248295 380765
rect 254485 380764 254551 380765
rect 255865 380764 255931 380765
rect 313457 380764 313523 380765
rect 438485 380764 438551 380765
rect 440877 380764 440943 380765
rect 443453 380764 443519 380765
rect 448237 380764 448303 380765
rect 235993 380760 236054 380764
rect 235993 380704 235998 380760
rect 217612 380700 217618 380702
rect 235993 380700 236054 380704
rect 236118 380762 236124 380764
rect 236118 380702 236150 380762
rect 237097 380760 237142 380764
rect 237206 380762 237212 380764
rect 237097 380704 237102 380760
rect 236118 380700 236124 380702
rect 237097 380700 237142 380704
rect 237206 380702 237254 380762
rect 243077 380760 243126 380764
rect 243190 380762 243196 380764
rect 243077 380704 243082 380760
rect 237206 380700 237212 380702
rect 243077 380700 243126 380704
rect 243190 380702 243234 380762
rect 248229 380760 248294 380764
rect 248229 380704 248234 380760
rect 248290 380704 248294 380760
rect 243190 380700 243196 380702
rect 248229 380700 248294 380704
rect 248358 380762 248364 380764
rect 248358 380702 248386 380762
rect 254485 380760 254550 380764
rect 254485 380704 254490 380760
rect 254546 380704 254550 380760
rect 248358 380700 248364 380702
rect 254485 380700 254550 380704
rect 254614 380762 254620 380764
rect 254614 380702 254642 380762
rect 255865 380760 255910 380764
rect 255974 380762 255980 380764
rect 313432 380762 313438 380764
rect 255865 380704 255870 380760
rect 254614 380700 254620 380702
rect 255865 380700 255910 380704
rect 255974 380702 256022 380762
rect 313366 380702 313438 380762
rect 313502 380760 313523 380764
rect 438480 380762 438486 380764
rect 313518 380704 313523 380760
rect 255974 380700 255980 380702
rect 313432 380700 313438 380702
rect 313502 380700 313523 380704
rect 438394 380702 438486 380762
rect 438480 380700 438486 380702
rect 438550 380700 438556 380764
rect 440877 380760 440934 380764
rect 440998 380762 441004 380764
rect 440877 380704 440882 380760
rect 440877 380700 440934 380704
rect 440998 380702 441034 380762
rect 443453 380760 443518 380764
rect 443453 380704 443458 380760
rect 443514 380704 443518 380760
rect 440998 380700 441004 380702
rect 443453 380700 443518 380704
rect 443582 380762 443588 380764
rect 443582 380702 443610 380762
rect 448237 380760 448278 380764
rect 448342 380762 448348 380764
rect 448237 380704 448242 380760
rect 443582 380700 443588 380702
rect 448237 380700 448278 380704
rect 448342 380702 448394 380762
rect 448342 380700 448348 380702
rect 235993 380699 236059 380700
rect 237097 380699 237163 380700
rect 243077 380699 243143 380700
rect 248229 380699 248295 380700
rect 254485 380699 254551 380700
rect 255865 380699 255931 380700
rect 313457 380699 313523 380700
rect 438485 380699 438551 380700
rect 440877 380699 440943 380700
rect 443453 380699 443519 380700
rect 448237 380699 448303 380700
rect 94544 380564 94550 380628
rect 94614 380626 94620 380628
rect 212625 380626 212691 380629
rect 258073 380628 258139 380629
rect 261753 380628 261819 380629
rect 270953 380628 271019 380629
rect 315849 380628 315915 380629
rect 404169 380628 404235 380629
rect 405457 380628 405523 380629
rect 413461 380628 413527 380629
rect 445937 380628 446003 380629
rect 503345 380628 503411 380629
rect 256992 380626 256998 380628
rect 94614 380624 212691 380626
rect 94614 380568 212630 380624
rect 212686 380568 212691 380624
rect 94614 380566 212691 380568
rect 94614 380564 94620 380566
rect 212625 380563 212691 380566
rect 219390 380566 256998 380626
rect 212993 380490 213059 380493
rect 103470 380488 213059 380490
rect 103470 380432 212998 380488
rect 213054 380432 213059 380488
rect 103470 380430 213059 380432
rect 95918 380292 95924 380356
rect 95988 380354 95994 380356
rect 103470 380354 103530 380430
rect 212993 380427 213059 380430
rect 95988 380294 103530 380354
rect 110965 380356 111031 380357
rect 113541 380356 113607 380357
rect 115933 380356 115999 380357
rect 118325 380356 118391 380357
rect 120993 380356 121059 380357
rect 110965 380352 111012 380356
rect 111076 380354 111082 380356
rect 110965 380296 110970 380352
rect 95988 380292 95994 380294
rect 110965 380292 111012 380296
rect 111076 380294 111122 380354
rect 113541 380352 113588 380356
rect 113652 380354 113658 380356
rect 113541 380296 113546 380352
rect 111076 380292 111082 380294
rect 113541 380292 113588 380296
rect 113652 380294 113698 380354
rect 115933 380352 115980 380356
rect 116044 380354 116050 380356
rect 115933 380296 115938 380352
rect 113652 380292 113658 380294
rect 115933 380292 115980 380296
rect 116044 380294 116090 380354
rect 118325 380352 118372 380356
rect 118436 380354 118442 380356
rect 120942 380354 120948 380356
rect 118325 380296 118330 380352
rect 116044 380292 116050 380294
rect 118325 380292 118372 380296
rect 118436 380294 118482 380354
rect 120902 380294 120948 380354
rect 121012 380352 121059 380356
rect 121054 380296 121059 380352
rect 118436 380292 118442 380294
rect 120942 380292 120948 380294
rect 121012 380292 121059 380296
rect 110965 380291 111031 380292
rect 113541 380291 113607 380292
rect 115933 380291 115999 380292
rect 118325 380291 118391 380292
rect 120993 380291 121059 380292
rect 123477 380356 123543 380357
rect 128353 380356 128419 380357
rect 135897 380356 135963 380357
rect 143625 380356 143691 380357
rect 148593 380356 148659 380357
rect 155953 380356 156019 380357
rect 158529 380356 158595 380357
rect 160921 380356 160987 380357
rect 163497 380356 163563 380357
rect 166073 380356 166139 380357
rect 123477 380352 123524 380356
rect 123588 380354 123594 380356
rect 128302 380354 128308 380356
rect 123477 380296 123482 380352
rect 123477 380292 123524 380296
rect 123588 380294 123634 380354
rect 128262 380294 128308 380354
rect 128372 380352 128419 380356
rect 135846 380354 135852 380356
rect 128414 380296 128419 380352
rect 123588 380292 123594 380294
rect 128302 380292 128308 380294
rect 128372 380292 128419 380296
rect 135806 380294 135852 380354
rect 135916 380352 135963 380356
rect 143574 380354 143580 380356
rect 135958 380296 135963 380352
rect 135846 380292 135852 380294
rect 135916 380292 135963 380296
rect 143534 380294 143580 380354
rect 143644 380352 143691 380356
rect 148542 380354 148548 380356
rect 143686 380296 143691 380352
rect 143574 380292 143580 380294
rect 143644 380292 143691 380296
rect 148502 380294 148548 380354
rect 148612 380352 148659 380356
rect 155902 380354 155908 380356
rect 148654 380296 148659 380352
rect 148542 380292 148548 380294
rect 148612 380292 148659 380296
rect 155862 380294 155908 380354
rect 155972 380352 156019 380356
rect 158478 380354 158484 380356
rect 156014 380296 156019 380352
rect 155902 380292 155908 380294
rect 155972 380292 156019 380296
rect 158438 380294 158484 380354
rect 158548 380352 158595 380356
rect 160870 380354 160876 380356
rect 158590 380296 158595 380352
rect 158478 380292 158484 380294
rect 158548 380292 158595 380296
rect 160830 380294 160876 380354
rect 160940 380352 160987 380356
rect 163446 380354 163452 380356
rect 160982 380296 160987 380352
rect 160870 380292 160876 380294
rect 160940 380292 160987 380296
rect 163406 380294 163452 380354
rect 163516 380352 163563 380356
rect 166022 380354 166028 380356
rect 163558 380296 163563 380352
rect 163446 380292 163452 380294
rect 163516 380292 163563 380296
rect 165982 380294 166028 380354
rect 166092 380352 166139 380356
rect 166134 380296 166139 380352
rect 166022 380292 166028 380294
rect 166092 380292 166139 380296
rect 123477 380291 123543 380292
rect 128353 380291 128419 380292
rect 135897 380291 135963 380292
rect 143625 380291 143691 380292
rect 148593 380291 148659 380292
rect 155953 380291 156019 380292
rect 158529 380291 158595 380292
rect 160921 380291 160987 380292
rect 163497 380291 163563 380292
rect 166073 380291 166139 380292
rect 207013 380354 207079 380357
rect 215293 380354 215359 380357
rect 207013 380352 215359 380354
rect 207013 380296 207018 380352
rect 207074 380296 215298 380352
rect 215354 380296 215359 380352
rect 207013 380294 215359 380296
rect 207013 380291 207079 380294
rect 215293 380291 215359 380294
rect 99373 380218 99439 380221
rect 204713 380218 204779 380221
rect 99373 380216 204779 380218
rect 99373 380160 99378 380216
rect 99434 380160 204718 380216
rect 204774 380160 204779 380216
rect 99373 380158 204779 380160
rect 99373 380155 99439 380158
rect 204713 380155 204779 380158
rect 205909 380218 205975 380221
rect 216622 380218 216628 380220
rect 205909 380216 216628 380218
rect 205909 380160 205914 380216
rect 205970 380160 216628 380216
rect 205909 380158 216628 380160
rect 205909 380155 205975 380158
rect 216622 380156 216628 380158
rect 216692 380218 216698 380220
rect 219390 380218 219450 380566
rect 256992 380564 256998 380566
rect 257062 380564 257068 380628
rect 258073 380624 258086 380628
rect 258150 380626 258156 380628
rect 258073 380568 258078 380624
rect 258073 380564 258086 380568
rect 258150 380566 258230 380626
rect 258150 380564 258156 380566
rect 261752 380564 261758 380628
rect 261822 380626 261828 380628
rect 261822 380566 261910 380626
rect 270953 380624 271006 380628
rect 271070 380626 271076 380628
rect 270953 380568 270958 380624
rect 261822 380564 261828 380566
rect 270953 380564 271006 380568
rect 271070 380566 271110 380626
rect 315849 380624 315886 380628
rect 315950 380626 315956 380628
rect 315849 380568 315854 380624
rect 271070 380564 271076 380566
rect 315849 380564 315886 380568
rect 315950 380566 316006 380626
rect 404169 380624 404214 380628
rect 404278 380626 404284 380628
rect 405432 380626 405438 380628
rect 404169 380568 404174 380624
rect 315950 380564 315956 380566
rect 404169 380564 404214 380568
rect 404278 380566 404326 380626
rect 405366 380566 405438 380626
rect 405502 380624 405523 380628
rect 413456 380626 413462 380628
rect 405518 380568 405523 380624
rect 404278 380564 404284 380566
rect 405432 380564 405438 380566
rect 405502 380564 405523 380568
rect 413370 380566 413462 380626
rect 413456 380564 413462 380566
rect 413526 380564 413532 380628
rect 445937 380624 445966 380628
rect 446030 380626 446036 380628
rect 445937 380568 445942 380624
rect 445937 380564 445966 380568
rect 446030 380566 446094 380626
rect 503345 380624 503358 380628
rect 503422 380626 503428 380628
rect 503345 380568 503350 380624
rect 446030 380564 446036 380566
rect 503345 380564 503358 380568
rect 503422 380566 503502 380626
rect 503422 380564 503428 380566
rect 258073 380563 258139 380564
rect 261753 380563 261819 380564
rect 270953 380563 271019 380564
rect 315849 380563 315915 380564
rect 404169 380563 404235 380564
rect 405457 380563 405523 380564
rect 413461 380563 413527 380564
rect 445937 380563 446003 380564
rect 503345 380563 503411 380564
rect 244273 380492 244339 380493
rect 244222 380490 244228 380492
rect 244182 380430 244228 380490
rect 244292 380488 244339 380492
rect 244334 380432 244339 380488
rect 244222 380428 244228 380430
rect 244292 380428 244339 380432
rect 244273 380427 244339 380428
rect 220721 380354 220787 380357
rect 247534 380354 247540 380356
rect 220721 380352 247540 380354
rect 220721 380296 220726 380352
rect 220782 380296 247540 380352
rect 220721 380294 247540 380296
rect 220721 380291 220787 380294
rect 247534 380292 247540 380294
rect 247604 380292 247610 380356
rect 216692 380158 219450 380218
rect 216692 380156 216698 380158
rect 359590 380156 359596 380220
rect 359660 380218 359666 380220
rect 380893 380218 380959 380221
rect 427486 380218 427492 380220
rect 359660 380216 427492 380218
rect 359660 380160 380898 380216
rect 380954 380160 427492 380216
rect 359660 380158 427492 380160
rect 359660 380156 359666 380158
rect 380893 380155 380959 380158
rect 427486 380156 427492 380158
rect 427556 380156 427562 380220
rect 214373 380082 214439 380085
rect 259494 380082 259500 380084
rect 214373 380080 259500 380082
rect 214373 380024 214378 380080
rect 214434 380024 259500 380080
rect 214373 380022 259500 380024
rect 214373 380019 214439 380022
rect 259494 380020 259500 380022
rect 259564 380020 259570 380084
rect 204713 379946 204779 379949
rect 208301 379946 208367 379949
rect 204713 379944 208367 379946
rect 204713 379888 204718 379944
rect 204774 379888 208306 379944
rect 208362 379888 208367 379944
rect 204713 379886 208367 379888
rect 204713 379883 204779 379886
rect 208301 379883 208367 379886
rect 212993 379810 213059 379813
rect 217961 379810 218027 379813
rect 212993 379808 218027 379810
rect 212993 379752 212998 379808
rect 213054 379752 217966 379808
rect 218022 379752 218027 379808
rect 212993 379750 218027 379752
rect 212993 379747 213059 379750
rect 217961 379747 218027 379750
rect 217317 379676 217383 379677
rect 217317 379672 217364 379676
rect 217428 379674 217434 379676
rect 217317 379616 217322 379672
rect 217317 379612 217364 379616
rect 217428 379614 217474 379674
rect 217428 379612 217434 379614
rect 217317 379611 217383 379612
rect 51942 379476 51948 379540
rect 52012 379538 52018 379540
rect 52177 379538 52243 379541
rect 52012 379536 52243 379538
rect 52012 379480 52182 379536
rect 52238 379480 52243 379536
rect 52012 379478 52243 379480
rect 52012 379476 52018 379478
rect 52177 379475 52243 379478
rect 209814 379476 209820 379540
rect 209884 379538 209890 379540
rect 211061 379538 211127 379541
rect 209884 379536 211127 379538
rect 209884 379480 211066 379536
rect 211122 379480 211127 379536
rect 209884 379478 211127 379480
rect 209884 379476 209890 379478
rect 211061 379475 211127 379478
rect 218830 379476 218836 379540
rect 218900 379538 218906 379540
rect 219341 379538 219407 379541
rect 218900 379536 219407 379538
rect 218900 379480 219346 379536
rect 219402 379480 219407 379536
rect 218900 379478 219407 379480
rect 218900 379476 218906 379478
rect 219341 379475 219407 379478
rect 360142 379476 360148 379540
rect 360212 379538 360218 379540
rect 361481 379538 361547 379541
rect 360212 379536 361547 379538
rect 360212 379480 361486 379536
rect 361542 379480 361547 379536
rect 360212 379478 361547 379480
rect 360212 379476 360218 379478
rect 361481 379475 361547 379478
rect 371601 379538 371667 379541
rect 378225 379538 378291 379541
rect 371601 379536 378291 379538
rect 371601 379480 371606 379536
rect 371662 379480 378230 379536
rect 378286 379480 378291 379536
rect 371601 379478 378291 379480
rect 371601 379475 371667 379478
rect 378225 379475 378291 379478
rect 46105 379402 46171 379405
rect 77201 379404 77267 379405
rect 77150 379402 77156 379404
rect 46105 379400 77034 379402
rect 46105 379344 46110 379400
rect 46166 379344 77034 379400
rect 46105 379342 77034 379344
rect 77110 379342 77156 379402
rect 77220 379400 77267 379404
rect 77262 379344 77267 379400
rect 46105 379339 46171 379342
rect 47669 379266 47735 379269
rect 76833 379266 76899 379269
rect 47669 379264 76899 379266
rect 47669 379208 47674 379264
rect 47730 379208 76838 379264
rect 76894 379208 76899 379264
rect 47669 379206 76899 379208
rect 76974 379266 77034 379342
rect 77150 379340 77156 379342
rect 77220 379340 77267 379344
rect 77201 379339 77267 379340
rect 80421 379404 80487 379405
rect 85481 379404 85547 379405
rect 86585 379404 86651 379405
rect 80421 379400 80468 379404
rect 80532 379402 80538 379404
rect 85430 379402 85436 379404
rect 80421 379344 80426 379400
rect 80421 379340 80468 379344
rect 80532 379342 80578 379402
rect 85390 379342 85436 379402
rect 85500 379400 85547 379404
rect 86534 379402 86540 379404
rect 85542 379344 85547 379400
rect 80532 379340 80538 379342
rect 85430 379340 85436 379342
rect 85500 379340 85547 379344
rect 86494 379342 86540 379402
rect 86604 379400 86651 379404
rect 86646 379344 86651 379400
rect 86534 379340 86540 379342
rect 86604 379340 86651 379344
rect 80421 379339 80487 379340
rect 85481 379339 85547 379340
rect 86585 379339 86651 379340
rect 88333 379404 88399 379405
rect 88793 379404 88859 379405
rect 88333 379400 88380 379404
rect 88444 379402 88450 379404
rect 88742 379402 88748 379404
rect 88333 379344 88338 379400
rect 88333 379340 88380 379344
rect 88444 379342 88490 379402
rect 88702 379342 88748 379402
rect 88812 379400 88859 379404
rect 88854 379344 88859 379400
rect 88444 379340 88450 379342
rect 88742 379340 88748 379342
rect 88812 379340 88859 379344
rect 88333 379339 88399 379340
rect 88793 379339 88859 379340
rect 90725 379404 90791 379405
rect 91369 379404 91435 379405
rect 90725 379400 90772 379404
rect 90836 379402 90842 379404
rect 91318 379402 91324 379404
rect 90725 379344 90730 379400
rect 90725 379340 90772 379344
rect 90836 379342 90882 379402
rect 91278 379342 91324 379402
rect 91388 379400 91435 379404
rect 91430 379344 91435 379400
rect 90836 379340 90842 379342
rect 91318 379340 91324 379342
rect 91388 379340 91435 379344
rect 90725 379339 90791 379340
rect 91369 379339 91435 379340
rect 92381 379404 92447 379405
rect 92381 379400 92428 379404
rect 92492 379402 92498 379404
rect 92381 379344 92386 379400
rect 92381 379340 92428 379344
rect 92492 379342 92538 379402
rect 92492 379340 92498 379342
rect 93342 379340 93348 379404
rect 93412 379402 93418 379404
rect 93577 379402 93643 379405
rect 93412 379400 93643 379402
rect 93412 379344 93582 379400
rect 93638 379344 93643 379400
rect 93412 379342 93643 379344
rect 93412 379340 93418 379342
rect 92381 379339 92447 379340
rect 93577 379339 93643 379342
rect 96061 379404 96127 379405
rect 98453 379404 98519 379405
rect 101029 379404 101095 379405
rect 96061 379400 96108 379404
rect 96172 379402 96178 379404
rect 96061 379344 96066 379400
rect 96061 379340 96108 379344
rect 96172 379342 96218 379402
rect 98453 379400 98500 379404
rect 98564 379402 98570 379404
rect 98453 379344 98458 379400
rect 96172 379340 96178 379342
rect 98453 379340 98500 379344
rect 98564 379342 98610 379402
rect 101029 379400 101076 379404
rect 101140 379402 101146 379404
rect 101029 379344 101034 379400
rect 98564 379340 98570 379342
rect 101029 379340 101076 379344
rect 101140 379342 101186 379402
rect 101140 379340 101146 379342
rect 103278 379340 103284 379404
rect 103348 379402 103354 379404
rect 103513 379402 103579 379405
rect 103348 379400 103579 379402
rect 103348 379344 103518 379400
rect 103574 379344 103579 379400
rect 103348 379342 103579 379344
rect 103348 379340 103354 379342
rect 96061 379339 96127 379340
rect 98453 379339 98519 379340
rect 101029 379339 101095 379340
rect 103513 379339 103579 379342
rect 105353 379402 105419 379405
rect 108205 379404 108271 379405
rect 108849 379404 108915 379405
rect 109769 379404 109835 379405
rect 111241 379404 111307 379405
rect 112345 379404 112411 379405
rect 113449 379404 113515 379405
rect 105854 379402 105860 379404
rect 105353 379400 105860 379402
rect 105353 379344 105358 379400
rect 105414 379344 105860 379400
rect 105353 379342 105860 379344
rect 105353 379339 105419 379342
rect 105854 379340 105860 379342
rect 105924 379340 105930 379404
rect 108205 379400 108252 379404
rect 108316 379402 108322 379404
rect 108798 379402 108804 379404
rect 108205 379344 108210 379400
rect 108205 379340 108252 379344
rect 108316 379342 108362 379402
rect 108758 379342 108804 379402
rect 108868 379400 108915 379404
rect 109718 379402 109724 379404
rect 108910 379344 108915 379400
rect 108316 379340 108322 379342
rect 108798 379340 108804 379342
rect 108868 379340 108915 379344
rect 109678 379342 109724 379402
rect 109788 379400 109835 379404
rect 111190 379402 111196 379404
rect 109830 379344 109835 379400
rect 109718 379340 109724 379342
rect 109788 379340 109835 379344
rect 111150 379342 111196 379402
rect 111260 379400 111307 379404
rect 112294 379402 112300 379404
rect 111302 379344 111307 379400
rect 111190 379340 111196 379342
rect 111260 379340 111307 379344
rect 112254 379342 112300 379402
rect 112364 379400 112411 379404
rect 113398 379402 113404 379404
rect 112406 379344 112411 379400
rect 112294 379340 112300 379342
rect 112364 379340 112411 379344
rect 113358 379342 113404 379402
rect 113468 379400 113515 379404
rect 113510 379344 113515 379400
rect 113398 379340 113404 379342
rect 113468 379340 113515 379344
rect 108205 379339 108271 379340
rect 108849 379339 108915 379340
rect 109769 379339 109835 379340
rect 111241 379339 111307 379340
rect 112345 379339 112411 379340
rect 113449 379339 113515 379340
rect 114461 379404 114527 379405
rect 115841 379404 115907 379405
rect 117129 379404 117195 379405
rect 141049 379404 141115 379405
rect 146017 379404 146083 379405
rect 150985 379404 151051 379405
rect 153561 379404 153627 379405
rect 114461 379400 114508 379404
rect 114572 379402 114578 379404
rect 115790 379402 115796 379404
rect 114461 379344 114466 379400
rect 114461 379340 114508 379344
rect 114572 379342 114618 379402
rect 115750 379342 115796 379402
rect 115860 379400 115907 379404
rect 117078 379402 117084 379404
rect 115902 379344 115907 379400
rect 114572 379340 114578 379342
rect 115790 379340 115796 379342
rect 115860 379340 115907 379344
rect 117038 379342 117084 379402
rect 117148 379400 117195 379404
rect 140998 379402 141004 379404
rect 117190 379344 117195 379400
rect 117078 379340 117084 379342
rect 117148 379340 117195 379344
rect 140958 379342 141004 379402
rect 141068 379400 141115 379404
rect 145966 379402 145972 379404
rect 141110 379344 141115 379400
rect 140998 379340 141004 379342
rect 141068 379340 141115 379344
rect 145926 379342 145972 379402
rect 146036 379400 146083 379404
rect 150934 379402 150940 379404
rect 146078 379344 146083 379400
rect 145966 379340 145972 379342
rect 146036 379340 146083 379344
rect 150894 379342 150940 379402
rect 151004 379400 151051 379404
rect 153510 379402 153516 379404
rect 151046 379344 151051 379400
rect 150934 379340 150940 379342
rect 151004 379340 151051 379344
rect 153470 379342 153516 379402
rect 153580 379400 153627 379404
rect 153622 379344 153627 379400
rect 153510 379340 153516 379342
rect 153580 379340 153627 379344
rect 114461 379339 114527 379340
rect 115841 379339 115907 379340
rect 117129 379339 117195 379340
rect 141049 379339 141115 379340
rect 146017 379339 146083 379340
rect 150985 379339 151051 379340
rect 153561 379339 153627 379340
rect 212993 379402 213059 379405
rect 220077 379402 220143 379405
rect 220721 379402 220787 379405
rect 212993 379400 220787 379402
rect 212993 379344 212998 379400
rect 213054 379344 220082 379400
rect 220138 379344 220726 379400
rect 220782 379344 220787 379400
rect 212993 379342 220787 379344
rect 212993 379339 213059 379342
rect 220077 379339 220143 379342
rect 220721 379339 220787 379342
rect 239581 379404 239647 379405
rect 239581 379400 239628 379404
rect 239692 379402 239698 379404
rect 244917 379402 244983 379405
rect 245326 379402 245332 379404
rect 239581 379344 239586 379400
rect 239581 379340 239628 379344
rect 239692 379342 239738 379402
rect 244917 379400 245332 379402
rect 244917 379344 244922 379400
rect 244978 379344 245332 379400
rect 244917 379342 245332 379344
rect 239692 379340 239698 379342
rect 239581 379339 239647 379340
rect 244917 379339 244983 379342
rect 245326 379340 245332 379342
rect 245396 379340 245402 379404
rect 246205 379402 246271 379405
rect 248597 379404 248663 379405
rect 250069 379404 250135 379405
rect 251173 379404 251239 379405
rect 252277 379404 252343 379405
rect 253381 379404 253447 379405
rect 263869 379404 263935 379405
rect 246430 379402 246436 379404
rect 246205 379400 246436 379402
rect 246205 379344 246210 379400
rect 246266 379344 246436 379400
rect 246205 379342 246436 379344
rect 246205 379339 246271 379342
rect 246430 379340 246436 379342
rect 246500 379340 246506 379404
rect 248597 379400 248644 379404
rect 248708 379402 248714 379404
rect 248597 379344 248602 379400
rect 248597 379340 248644 379344
rect 248708 379342 248754 379402
rect 250069 379400 250116 379404
rect 250180 379402 250186 379404
rect 250069 379344 250074 379400
rect 248708 379340 248714 379342
rect 250069 379340 250116 379344
rect 250180 379342 250226 379402
rect 251173 379400 251220 379404
rect 251284 379402 251290 379404
rect 251173 379344 251178 379400
rect 250180 379340 250186 379342
rect 251173 379340 251220 379344
rect 251284 379342 251330 379402
rect 252277 379400 252324 379404
rect 252388 379402 252394 379404
rect 252277 379344 252282 379400
rect 251284 379340 251290 379342
rect 252277 379340 252324 379344
rect 252388 379342 252434 379402
rect 253381 379400 253428 379404
rect 253492 379402 253498 379404
rect 253381 379344 253386 379400
rect 252388 379340 252394 379342
rect 253381 379340 253428 379344
rect 253492 379342 253538 379402
rect 263869 379400 263916 379404
rect 263980 379402 263986 379404
rect 264973 379402 265039 379405
rect 265198 379402 265204 379404
rect 263869 379344 263874 379400
rect 253492 379340 253498 379342
rect 263869 379340 263916 379344
rect 263980 379342 264026 379402
rect 264973 379400 265204 379402
rect 264973 379344 264978 379400
rect 265034 379344 265204 379400
rect 264973 379342 265204 379344
rect 263980 379340 263986 379342
rect 248597 379339 248663 379340
rect 250069 379339 250135 379340
rect 251173 379339 251239 379340
rect 252277 379339 252343 379340
rect 253381 379339 253447 379340
rect 263869 379339 263935 379340
rect 264973 379339 265039 379342
rect 265198 379340 265204 379342
rect 265268 379340 265274 379404
rect 268285 379402 268351 379405
rect 269757 379404 269823 379405
rect 271045 379404 271111 379405
rect 272149 379404 272215 379405
rect 273253 379404 273319 379405
rect 275737 379404 275803 379405
rect 268694 379402 268700 379404
rect 268285 379400 268700 379402
rect 268285 379344 268290 379400
rect 268346 379344 268700 379400
rect 268285 379342 268700 379344
rect 268285 379339 268351 379342
rect 268694 379340 268700 379342
rect 268764 379340 268770 379404
rect 269757 379400 269804 379404
rect 269868 379402 269874 379404
rect 269757 379344 269762 379400
rect 269757 379340 269804 379344
rect 269868 379342 269914 379402
rect 271045 379400 271092 379404
rect 271156 379402 271162 379404
rect 271045 379344 271050 379400
rect 269868 379340 269874 379342
rect 271045 379340 271092 379344
rect 271156 379342 271202 379402
rect 272149 379400 272196 379404
rect 272260 379402 272266 379404
rect 272149 379344 272154 379400
rect 271156 379340 271162 379342
rect 272149 379340 272196 379344
rect 272260 379342 272306 379402
rect 273253 379400 273300 379404
rect 273364 379402 273370 379404
rect 275686 379402 275692 379404
rect 273253 379344 273258 379400
rect 272260 379340 272266 379342
rect 273253 379340 273300 379344
rect 273364 379342 273410 379402
rect 275646 379342 275692 379402
rect 275756 379400 275803 379404
rect 275798 379344 275803 379400
rect 273364 379340 273370 379342
rect 275686 379340 275692 379342
rect 275756 379340 275803 379344
rect 269757 379339 269823 379340
rect 271045 379339 271111 379340
rect 272149 379339 272215 379340
rect 273253 379339 273319 379340
rect 275737 379339 275803 379340
rect 285949 379404 286015 379405
rect 285949 379400 285996 379404
rect 286060 379402 286066 379404
rect 287697 379402 287763 379405
rect 288198 379402 288204 379404
rect 285949 379344 285954 379400
rect 285949 379340 285996 379344
rect 286060 379342 286106 379402
rect 287697 379400 288204 379402
rect 287697 379344 287702 379400
rect 287758 379344 288204 379400
rect 287697 379342 288204 379344
rect 286060 379340 286066 379342
rect 285949 379339 286015 379340
rect 287697 379339 287763 379342
rect 288198 379340 288204 379342
rect 288268 379340 288274 379404
rect 290181 379402 290247 379405
rect 293309 379404 293375 379405
rect 295885 379404 295951 379405
rect 290958 379402 290964 379404
rect 290181 379400 290964 379402
rect 290181 379344 290186 379400
rect 290242 379344 290964 379400
rect 290181 379342 290964 379344
rect 290181 379339 290247 379342
rect 290958 379340 290964 379342
rect 291028 379340 291034 379404
rect 293309 379400 293356 379404
rect 293420 379402 293426 379404
rect 293309 379344 293314 379400
rect 293309 379340 293356 379344
rect 293420 379342 293466 379402
rect 295885 379400 295932 379404
rect 295996 379402 296002 379404
rect 298093 379402 298159 379405
rect 305821 379404 305887 379405
rect 298502 379402 298508 379404
rect 295885 379344 295890 379400
rect 293420 379340 293426 379342
rect 295885 379340 295932 379344
rect 295996 379342 296042 379402
rect 298093 379400 298508 379402
rect 298093 379344 298098 379400
rect 298154 379344 298508 379400
rect 298093 379342 298508 379344
rect 295996 379340 296002 379342
rect 293309 379339 293375 379340
rect 295885 379339 295951 379340
rect 298093 379339 298159 379342
rect 298502 379340 298508 379342
rect 298572 379340 298578 379404
rect 305821 379400 305868 379404
rect 305932 379402 305938 379404
rect 307845 379402 307911 379405
rect 310973 379404 311039 379405
rect 308438 379402 308444 379404
rect 305821 379344 305826 379400
rect 305821 379340 305868 379344
rect 305932 379342 305978 379402
rect 307845 379400 308444 379402
rect 307845 379344 307850 379400
rect 307906 379344 308444 379400
rect 307845 379342 308444 379344
rect 305932 379340 305938 379342
rect 305821 379339 305887 379340
rect 307845 379339 307911 379342
rect 308438 379340 308444 379342
rect 308508 379340 308514 379404
rect 310973 379400 311020 379404
rect 311084 379402 311090 379404
rect 317781 379402 317847 379405
rect 320909 379404 320975 379405
rect 325877 379404 325943 379405
rect 396073 379404 396139 379405
rect 318374 379402 318380 379404
rect 310973 379344 310978 379400
rect 310973 379340 311020 379344
rect 311084 379342 311130 379402
rect 317781 379400 318380 379402
rect 317781 379344 317786 379400
rect 317842 379344 318380 379400
rect 317781 379342 318380 379344
rect 311084 379340 311090 379342
rect 310973 379339 311039 379340
rect 317781 379339 317847 379342
rect 318374 379340 318380 379342
rect 318444 379340 318450 379404
rect 320909 379400 320956 379404
rect 321020 379402 321026 379404
rect 320909 379344 320914 379400
rect 320909 379340 320956 379344
rect 321020 379342 321066 379402
rect 325877 379400 325924 379404
rect 325988 379402 325994 379404
rect 396022 379402 396028 379404
rect 325877 379344 325882 379400
rect 321020 379340 321026 379342
rect 325877 379340 325924 379344
rect 325988 379342 326034 379402
rect 395982 379342 396028 379402
rect 396092 379400 396139 379404
rect 396134 379344 396139 379400
rect 325988 379340 325994 379342
rect 396022 379340 396028 379342
rect 396092 379340 396139 379344
rect 320909 379339 320975 379340
rect 325877 379339 325943 379340
rect 396073 379339 396139 379340
rect 396349 379402 396415 379405
rect 398189 379404 398255 379405
rect 399477 379404 399543 379405
rect 397126 379402 397132 379404
rect 396349 379400 397132 379402
rect 396349 379344 396354 379400
rect 396410 379344 397132 379400
rect 396349 379342 397132 379344
rect 396349 379339 396415 379342
rect 397126 379340 397132 379342
rect 397196 379340 397202 379404
rect 398189 379400 398236 379404
rect 398300 379402 398306 379404
rect 398189 379344 398194 379400
rect 398189 379340 398236 379344
rect 398300 379342 398346 379402
rect 399477 379400 399524 379404
rect 399588 379402 399594 379404
rect 405825 379402 405891 379405
rect 407573 379404 407639 379405
rect 408309 379404 408375 379405
rect 406510 379402 406516 379404
rect 399477 379344 399482 379400
rect 398300 379340 398306 379342
rect 399477 379340 399524 379344
rect 399588 379342 399634 379402
rect 405825 379400 406516 379402
rect 405825 379344 405830 379400
rect 405886 379344 406516 379400
rect 405825 379342 406516 379344
rect 399588 379340 399594 379342
rect 398189 379339 398255 379340
rect 399477 379339 399543 379340
rect 405825 379339 405891 379342
rect 406510 379340 406516 379342
rect 406580 379340 406586 379404
rect 407573 379400 407620 379404
rect 407684 379402 407690 379404
rect 407573 379344 407578 379400
rect 407573 379340 407620 379344
rect 407684 379342 407730 379402
rect 408309 379400 408356 379404
rect 408420 379402 408426 379404
rect 410333 379402 410399 379405
rect 411253 379404 411319 379405
rect 412357 379404 412423 379405
rect 420637 379404 420703 379405
rect 428181 379404 428247 379405
rect 431125 379404 431191 379405
rect 434253 379404 434319 379405
rect 437933 379404 437999 379405
rect 450997 379404 451063 379405
rect 410742 379402 410748 379404
rect 408309 379344 408314 379400
rect 407684 379340 407690 379342
rect 408309 379340 408356 379344
rect 408420 379342 408466 379402
rect 410333 379400 410748 379402
rect 410333 379344 410338 379400
rect 410394 379344 410748 379400
rect 410333 379342 410748 379344
rect 408420 379340 408426 379342
rect 407573 379339 407639 379340
rect 408309 379339 408375 379340
rect 410333 379339 410399 379342
rect 410742 379340 410748 379342
rect 410812 379340 410818 379404
rect 411253 379400 411300 379404
rect 411364 379402 411370 379404
rect 411253 379344 411258 379400
rect 411253 379340 411300 379344
rect 411364 379342 411410 379402
rect 412357 379400 412404 379404
rect 412468 379402 412474 379404
rect 412357 379344 412362 379400
rect 411364 379340 411370 379342
rect 412357 379340 412404 379344
rect 412468 379342 412514 379402
rect 420637 379400 420684 379404
rect 420748 379402 420754 379404
rect 420637 379344 420642 379400
rect 412468 379340 412474 379342
rect 420637 379340 420684 379344
rect 420748 379342 420794 379402
rect 428181 379400 428228 379404
rect 428292 379402 428298 379404
rect 428181 379344 428186 379400
rect 420748 379340 420754 379342
rect 428181 379340 428228 379344
rect 428292 379342 428338 379402
rect 431125 379400 431172 379404
rect 431236 379402 431242 379404
rect 431125 379344 431130 379400
rect 428292 379340 428298 379342
rect 431125 379340 431172 379344
rect 431236 379342 431282 379402
rect 434253 379400 434300 379404
rect 434364 379402 434370 379404
rect 434253 379344 434258 379400
rect 431236 379340 431242 379342
rect 434253 379340 434300 379344
rect 434364 379342 434410 379402
rect 437933 379400 437980 379404
rect 438044 379402 438050 379404
rect 437933 379344 437938 379400
rect 434364 379340 434370 379342
rect 437933 379340 437980 379344
rect 438044 379342 438090 379402
rect 450997 379400 451044 379404
rect 451108 379402 451114 379404
rect 453021 379402 453087 379405
rect 453430 379402 453436 379404
rect 450997 379344 451002 379400
rect 438044 379340 438050 379342
rect 450997 379340 451044 379344
rect 451108 379342 451154 379402
rect 453021 379400 453436 379402
rect 453021 379344 453026 379400
rect 453082 379344 453436 379400
rect 453021 379342 453436 379344
rect 451108 379340 451114 379342
rect 411253 379339 411319 379340
rect 412357 379339 412423 379340
rect 420637 379339 420703 379340
rect 428181 379339 428247 379340
rect 431125 379339 431191 379340
rect 434253 379339 434319 379340
rect 437933 379339 437999 379340
rect 450997 379339 451063 379340
rect 453021 379339 453087 379342
rect 453430 379340 453436 379342
rect 453500 379340 453506 379404
rect 455597 379402 455663 379405
rect 460933 379404 460999 379405
rect 463509 379404 463575 379405
rect 473445 379404 473511 379405
rect 455822 379402 455828 379404
rect 455597 379400 455828 379402
rect 455597 379344 455602 379400
rect 455658 379344 455828 379400
rect 455597 379342 455828 379344
rect 455597 379339 455663 379342
rect 455822 379340 455828 379342
rect 455892 379340 455898 379404
rect 460933 379400 460980 379404
rect 461044 379402 461050 379404
rect 460933 379344 460938 379400
rect 460933 379340 460980 379344
rect 461044 379342 461090 379402
rect 463509 379400 463556 379404
rect 463620 379402 463626 379404
rect 463509 379344 463514 379400
rect 461044 379340 461050 379342
rect 463509 379340 463556 379344
rect 463620 379342 463666 379402
rect 473445 379400 473492 379404
rect 473556 379402 473562 379404
rect 480621 379402 480687 379405
rect 485957 379404 486023 379405
rect 480846 379402 480852 379404
rect 473445 379344 473450 379400
rect 463620 379340 463626 379342
rect 473445 379340 473492 379344
rect 473556 379342 473602 379402
rect 480621 379400 480852 379402
rect 480621 379344 480626 379400
rect 480682 379344 480852 379400
rect 480621 379342 480852 379344
rect 473556 379340 473562 379342
rect 460933 379339 460999 379340
rect 463509 379339 463575 379340
rect 473445 379339 473511 379340
rect 480621 379339 480687 379342
rect 480846 379340 480852 379342
rect 480916 379340 480922 379404
rect 485957 379400 486004 379404
rect 486068 379402 486074 379404
rect 485957 379344 485962 379400
rect 485957 379340 486004 379344
rect 486068 379342 486114 379402
rect 486068 379340 486074 379342
rect 503294 379340 503300 379404
rect 503364 379402 503370 379404
rect 503621 379402 503687 379405
rect 503364 379400 503687 379402
rect 503364 379344 503626 379400
rect 503682 379344 503687 379400
rect 503364 379342 503687 379344
rect 503364 379340 503370 379342
rect 485957 379339 486023 379340
rect 503621 379339 503687 379342
rect 78254 379266 78260 379268
rect 76974 379206 78260 379266
rect 47669 379203 47735 379206
rect 76833 379203 76899 379206
rect 78254 379204 78260 379206
rect 78324 379204 78330 379268
rect 81750 379204 81756 379268
rect 81820 379204 81826 379268
rect 90030 379204 90036 379268
rect 90100 379266 90106 379268
rect 90817 379266 90883 379269
rect 90100 379264 90883 379266
rect 90100 379208 90822 379264
rect 90878 379208 90883 379264
rect 90100 379206 90883 379208
rect 90100 379204 90106 379206
rect 44766 379068 44772 379132
rect 44836 379130 44842 379132
rect 47485 379130 47551 379133
rect 81758 379130 81818 379204
rect 90817 379203 90883 379206
rect 93485 379266 93551 379269
rect 99465 379268 99531 379269
rect 102961 379268 103027 379269
rect 93710 379266 93716 379268
rect 93485 379264 93716 379266
rect 93485 379208 93490 379264
rect 93546 379208 93716 379264
rect 93485 379206 93716 379208
rect 93485 379203 93551 379206
rect 93710 379204 93716 379206
rect 93780 379204 93786 379268
rect 99414 379266 99420 379268
rect 99374 379206 99420 379266
rect 99484 379264 99531 379268
rect 102910 379266 102916 379268
rect 99526 379208 99531 379264
rect 99414 379204 99420 379206
rect 99484 379204 99531 379208
rect 102870 379206 102916 379266
rect 102980 379264 103027 379268
rect 103022 379208 103027 379264
rect 102910 379204 102916 379206
rect 102980 379204 103027 379208
rect 104014 379204 104020 379268
rect 104084 379266 104090 379268
rect 104249 379266 104315 379269
rect 104084 379264 104315 379266
rect 104084 379208 104254 379264
rect 104310 379208 104315 379264
rect 104084 379206 104315 379208
rect 104084 379204 104090 379206
rect 99465 379203 99531 379204
rect 102961 379203 103027 379204
rect 104249 379203 104315 379206
rect 118182 379204 118188 379268
rect 118252 379266 118258 379268
rect 213821 379266 213887 379269
rect 238201 379268 238267 379269
rect 276105 379268 276171 379269
rect 277025 379268 277091 379269
rect 238150 379266 238156 379268
rect 118252 379264 213887 379266
rect 118252 379208 213826 379264
rect 213882 379208 213887 379264
rect 118252 379206 213887 379208
rect 238110 379206 238156 379266
rect 238220 379264 238267 379268
rect 274398 379266 274404 379268
rect 238262 379208 238267 379264
rect 118252 379204 118258 379206
rect 213821 379203 213887 379206
rect 238150 379204 238156 379206
rect 238220 379204 238267 379208
rect 238201 379203 238267 379204
rect 238710 379206 274404 379266
rect 204253 379130 204319 379133
rect 205725 379130 205791 379133
rect 44836 379128 204319 379130
rect 44836 379072 47490 379128
rect 47546 379072 204258 379128
rect 204314 379072 204319 379128
rect 44836 379070 204319 379072
rect 44836 379068 44842 379070
rect 47485 379067 47551 379070
rect 204253 379067 204319 379070
rect 204486 379128 205791 379130
rect 204486 379072 205730 379128
rect 205786 379072 205791 379128
rect 204486 379070 205791 379072
rect 78254 378932 78260 378996
rect 78324 378994 78330 378996
rect 204486 378994 204546 379070
rect 205725 379067 205791 379070
rect 207013 379130 207079 379133
rect 219985 379130 220051 379133
rect 238710 379130 238770 379206
rect 274398 379204 274404 379206
rect 274468 379204 274474 379268
rect 276054 379266 276060 379268
rect 276014 379206 276060 379266
rect 276124 379264 276171 379268
rect 276974 379266 276980 379268
rect 276166 379208 276171 379264
rect 276054 379204 276060 379206
rect 276124 379204 276171 379208
rect 276934 379206 276980 379266
rect 277044 379264 277091 379268
rect 277086 379208 277091 379264
rect 276974 379204 276980 379206
rect 277044 379204 277091 379208
rect 276105 379203 276171 379204
rect 277025 379203 277091 379204
rect 278405 379268 278471 379269
rect 280797 379268 280863 379269
rect 278405 379264 278452 379268
rect 278516 379266 278522 379268
rect 278405 379208 278410 379264
rect 278405 379204 278452 379208
rect 278516 379206 278562 379266
rect 280797 379264 280844 379268
rect 280908 379266 280914 379268
rect 283097 379266 283163 379269
rect 300853 379268 300919 379269
rect 402973 379268 403039 379269
rect 414565 379268 414631 379269
rect 415853 379268 415919 379269
rect 416037 379268 416103 379269
rect 283414 379266 283420 379268
rect 280797 379208 280802 379264
rect 278516 379204 278522 379206
rect 280797 379204 280844 379208
rect 280908 379206 280954 379266
rect 283097 379264 283420 379266
rect 283097 379208 283102 379264
rect 283158 379208 283420 379264
rect 283097 379206 283420 379208
rect 280908 379204 280914 379206
rect 278405 379203 278471 379204
rect 280797 379203 280863 379204
rect 283097 379203 283163 379206
rect 283414 379204 283420 379206
rect 283484 379204 283490 379268
rect 300853 379264 300900 379268
rect 300964 379266 300970 379268
rect 300853 379208 300858 379264
rect 300853 379204 300900 379208
rect 300964 379206 301010 379266
rect 300964 379204 300970 379206
rect 401726 379204 401732 379268
rect 401796 379204 401802 379268
rect 402973 379264 403020 379268
rect 403084 379266 403090 379268
rect 402973 379208 402978 379264
rect 402973 379204 403020 379208
rect 403084 379206 403130 379266
rect 414565 379264 414612 379268
rect 414676 379266 414682 379268
rect 415853 379266 415900 379268
rect 414565 379208 414570 379264
rect 403084 379204 403090 379206
rect 414565 379204 414612 379208
rect 414676 379206 414722 379266
rect 415808 379264 415900 379266
rect 415808 379208 415858 379264
rect 415808 379206 415900 379208
rect 414676 379204 414682 379206
rect 415853 379204 415900 379206
rect 415964 379204 415970 379268
rect 416037 379264 416084 379268
rect 416148 379266 416154 379268
rect 422845 379266 422911 379269
rect 423438 379266 423444 379268
rect 416037 379208 416042 379264
rect 416037 379204 416084 379208
rect 416148 379206 416194 379266
rect 422845 379264 423444 379266
rect 422845 379208 422850 379264
rect 422906 379208 423444 379264
rect 422845 379206 423444 379208
rect 416148 379204 416154 379206
rect 300853 379203 300919 379204
rect 343449 379132 343515 379133
rect 278078 379130 278084 379132
rect 207013 379128 238770 379130
rect 207013 379072 207018 379128
rect 207074 379072 219990 379128
rect 220046 379072 238770 379128
rect 207013 379070 238770 379072
rect 273302 379070 278084 379130
rect 207013 379067 207079 379070
rect 219985 379067 220051 379070
rect 78324 378934 204546 378994
rect 204713 378994 204779 378997
rect 209865 378994 209931 378997
rect 212993 378994 213059 378997
rect 204713 378992 213059 378994
rect 204713 378936 204718 378992
rect 204774 378936 209870 378992
rect 209926 378936 212998 378992
rect 213054 378936 213059 378992
rect 204713 378934 213059 378936
rect 78324 378932 78330 378934
rect 204713 378931 204779 378934
rect 209865 378931 209931 378934
rect 212993 378931 213059 378934
rect 213821 378994 213887 378997
rect 273302 378994 273362 379070
rect 277350 378997 277410 379070
rect 278078 379068 278084 379070
rect 278148 379068 278154 379132
rect 343398 379130 343404 379132
rect 343358 379070 343404 379130
rect 343468 379128 343515 379132
rect 343510 379072 343515 379128
rect 343398 379068 343404 379070
rect 343468 379068 343515 379072
rect 343449 379067 343515 379068
rect 369853 379130 369919 379133
rect 371049 379130 371115 379133
rect 400438 379130 400444 379132
rect 369853 379128 400444 379130
rect 369853 379072 369858 379128
rect 369914 379072 371054 379128
rect 371110 379072 400444 379128
rect 369853 379070 400444 379072
rect 369853 379067 369919 379070
rect 371049 379067 371115 379070
rect 400438 379068 400444 379070
rect 400508 379068 400514 379132
rect 213821 378992 273362 378994
rect 213821 378936 213826 378992
rect 213882 378936 273362 378992
rect 213821 378934 273362 378936
rect 273437 378996 273503 378997
rect 273437 378992 273484 378996
rect 273548 378994 273554 378996
rect 273437 378936 273442 378992
rect 213821 378931 213887 378934
rect 273437 378932 273484 378936
rect 273548 378934 273594 378994
rect 277301 378992 277410 378997
rect 277301 378936 277306 378992
rect 277362 378936 277410 378992
rect 277301 378934 277410 378936
rect 302509 378994 302575 378997
rect 303470 378994 303476 378996
rect 302509 378992 303476 378994
rect 302509 378936 302514 378992
rect 302570 378936 303476 378992
rect 302509 378934 303476 378936
rect 273548 378932 273554 378934
rect 273437 378931 273503 378932
rect 277301 378931 277367 378934
rect 302509 378931 302575 378934
rect 303470 378932 303476 378934
rect 303540 378932 303546 378996
rect 343214 378932 343220 378996
rect 343284 378994 343290 378996
rect 343541 378994 343607 378997
rect 401734 378994 401794 379204
rect 402973 379203 403039 379204
rect 414565 379203 414631 379204
rect 415853 379203 415919 379204
rect 416037 379203 416103 379204
rect 422845 379203 422911 379206
rect 423438 379204 423444 379206
rect 423508 379204 423514 379268
rect 419349 379132 419415 379133
rect 419349 379128 419396 379132
rect 419460 379130 419466 379132
rect 465073 379130 465139 379133
rect 465942 379130 465948 379132
rect 419349 379072 419354 379128
rect 419349 379068 419396 379072
rect 419460 379070 419506 379130
rect 465073 379128 465948 379130
rect 465073 379072 465078 379128
rect 465134 379072 465948 379128
rect 465073 379070 465948 379072
rect 419460 379068 419466 379070
rect 419349 379067 419415 379068
rect 465073 379067 465139 379070
rect 465942 379068 465948 379070
rect 466012 379068 466018 379132
rect 343284 378992 343607 378994
rect 343284 378936 343546 378992
rect 343602 378936 343607 378992
rect 343284 378934 343607 378936
rect 343284 378932 343290 378934
rect 343541 378931 343607 378934
rect 373950 378934 401794 378994
rect 470869 378996 470935 378997
rect 470869 378992 470916 378996
rect 470980 378994 470986 378996
rect 470869 378936 470874 378992
rect 76833 378858 76899 378861
rect 79542 378858 79548 378860
rect 76833 378856 79548 378858
rect 76833 378800 76838 378856
rect 76894 378800 79548 378856
rect 76833 378798 79548 378800
rect 76833 378795 76899 378798
rect 79542 378796 79548 378798
rect 79612 378858 79618 378860
rect 210325 378858 210391 378861
rect 79612 378856 210391 378858
rect 79612 378800 210330 378856
rect 210386 378800 210391 378856
rect 79612 378798 210391 378800
rect 79612 378796 79618 378798
rect 210325 378795 210391 378798
rect 250621 378860 250687 378861
rect 250621 378856 250668 378860
rect 250732 378858 250738 378860
rect 253197 378858 253263 378861
rect 372337 378858 372403 378861
rect 373950 378858 374010 378934
rect 470869 378932 470916 378936
rect 470980 378934 471026 378994
rect 470980 378932 470986 378934
rect 470869 378931 470935 378932
rect 250621 378800 250626 378856
rect 250621 378796 250668 378800
rect 250732 378798 250778 378858
rect 253197 378856 374010 378858
rect 253197 378800 253202 378856
rect 253258 378800 372342 378856
rect 372398 378800 374010 378856
rect 253197 378798 374010 378800
rect 250732 378796 250738 378798
rect 250621 378795 250687 378796
rect 253197 378795 253263 378798
rect 372337 378795 372403 378798
rect 377622 378796 377628 378860
rect 377692 378858 377698 378860
rect 381077 378858 381143 378861
rect 429694 378858 429700 378860
rect 377692 378856 429700 378858
rect 377692 378800 381082 378856
rect 381138 378800 429700 378856
rect 377692 378798 429700 378800
rect 377692 378796 377698 378798
rect 381077 378795 381143 378798
rect 429694 378796 429700 378798
rect 429764 378796 429770 378860
rect 467925 378858 467991 378861
rect 468518 378858 468524 378860
rect 467925 378856 468524 378858
rect 467925 378800 467930 378856
rect 467986 378800 468524 378856
rect 467925 378798 468524 378800
rect 467925 378795 467991 378798
rect 468518 378796 468524 378798
rect 468588 378796 468594 378860
rect 474733 378858 474799 378861
rect 475878 378858 475884 378860
rect 474733 378856 475884 378858
rect 474733 378800 474738 378856
rect 474794 378800 475884 378856
rect 474733 378798 475884 378800
rect 474733 378795 474799 378798
rect 475878 378796 475884 378798
rect 475948 378796 475954 378860
rect 477493 378858 477559 378861
rect 483381 378860 483447 378861
rect 478454 378858 478460 378860
rect 477493 378856 478460 378858
rect 477493 378800 477498 378856
rect 477554 378800 478460 378856
rect 477493 378798 478460 378800
rect 477493 378795 477559 378798
rect 478454 378796 478460 378798
rect 478524 378796 478530 378860
rect 483381 378856 483428 378860
rect 483492 378858 483498 378860
rect 483381 378800 483386 378856
rect 483381 378796 483428 378800
rect 483492 378798 483538 378858
rect 483492 378796 483498 378798
rect 483381 378795 483447 378796
rect 80421 378722 80487 378725
rect 220905 378722 220971 378725
rect 240542 378722 240548 378724
rect 80421 378720 240548 378722
rect 80421 378664 80426 378720
rect 80482 378664 220910 378720
rect 220966 378664 240548 378720
rect 80421 378662 240548 378664
rect 80421 378659 80487 378662
rect 220905 378659 220971 378662
rect 240542 378660 240548 378662
rect 240612 378722 240618 378724
rect 369853 378722 369919 378725
rect 240612 378720 369919 378722
rect 240612 378664 369858 378720
rect 369914 378664 369919 378720
rect 240612 378662 369919 378664
rect 240612 378660 240618 378662
rect 369853 378659 369919 378662
rect 377438 378660 377444 378724
rect 377508 378722 377514 378724
rect 381169 378722 381235 378725
rect 433374 378722 433380 378724
rect 377508 378720 433380 378722
rect 377508 378664 381174 378720
rect 381230 378664 433380 378720
rect 377508 378662 433380 378664
rect 377508 378660 377514 378662
rect 381169 378659 381235 378662
rect 433374 378660 433380 378662
rect 433444 378660 433450 378724
rect 76046 378524 76052 378588
rect 76116 378586 76122 378588
rect 77109 378586 77175 378589
rect 97073 378588 97139 378589
rect 97022 378586 97028 378588
rect 76116 378584 77175 378586
rect 76116 378528 77114 378584
rect 77170 378528 77175 378584
rect 76116 378526 77175 378528
rect 96982 378526 97028 378586
rect 97092 378584 97139 378588
rect 97134 378528 97139 378584
rect 76116 378524 76122 378526
rect 77109 378523 77175 378526
rect 97022 378524 97028 378526
rect 97092 378524 97139 378528
rect 98126 378524 98132 378588
rect 98196 378586 98202 378588
rect 98545 378586 98611 378589
rect 101857 378588 101923 378589
rect 107561 378588 107627 378589
rect 101806 378586 101812 378588
rect 98196 378584 98611 378586
rect 98196 378528 98550 378584
rect 98606 378528 98611 378584
rect 98196 378526 98611 378528
rect 101766 378526 101812 378586
rect 101876 378584 101923 378588
rect 107510 378586 107516 378588
rect 101918 378528 101923 378584
rect 98196 378524 98202 378526
rect 97073 378523 97139 378524
rect 98545 378523 98611 378526
rect 101806 378524 101812 378526
rect 101876 378524 101923 378528
rect 107470 378526 107516 378586
rect 107580 378584 107627 378588
rect 107622 378528 107627 378584
rect 107510 378524 107516 378526
rect 107580 378524 107627 378528
rect 119102 378524 119108 378588
rect 119172 378586 119178 378588
rect 204805 378586 204871 378589
rect 119172 378584 204871 378586
rect 119172 378528 204810 378584
rect 204866 378528 204871 378584
rect 119172 378526 204871 378528
rect 119172 378524 119178 378526
rect 101857 378523 101923 378524
rect 107561 378523 107627 378524
rect 204805 378523 204871 378526
rect 208342 378524 208348 378588
rect 208412 378586 208418 378588
rect 209681 378586 209747 378589
rect 208412 378584 209747 378586
rect 208412 378528 209686 378584
rect 209742 378528 209747 378584
rect 208412 378526 209747 378528
rect 208412 378524 208418 378526
rect 209681 378523 209747 378526
rect 220721 378586 220787 378589
rect 258349 378588 258415 378589
rect 260557 378588 260623 378589
rect 260925 378588 260991 378589
rect 262765 378588 262831 378589
rect 263593 378588 263659 378589
rect 220721 378584 258090 378586
rect 220721 378528 220726 378584
rect 220782 378528 258090 378584
rect 220721 378526 258090 378528
rect 220721 378523 220787 378526
rect 125961 378452 126027 378453
rect 125910 378450 125916 378452
rect 125870 378390 125916 378450
rect 125980 378448 126027 378452
rect 126022 378392 126027 378448
rect 125910 378388 125916 378390
rect 125980 378388 126027 378392
rect 125961 378387 126027 378388
rect 131021 378452 131087 378453
rect 133505 378452 133571 378453
rect 138473 378452 138539 378453
rect 131021 378448 131068 378452
rect 131132 378450 131138 378452
rect 133454 378450 133460 378452
rect 131021 378392 131026 378448
rect 131021 378388 131068 378392
rect 131132 378390 131178 378450
rect 133414 378390 133460 378450
rect 133524 378448 133571 378452
rect 138422 378450 138428 378452
rect 133566 378392 133571 378448
rect 131132 378388 131138 378390
rect 133454 378388 133460 378390
rect 133524 378388 133571 378392
rect 138382 378390 138428 378450
rect 138492 378448 138539 378452
rect 138534 378392 138539 378448
rect 138422 378388 138428 378390
rect 138492 378388 138539 378392
rect 131021 378387 131087 378388
rect 133505 378387 133571 378388
rect 138473 378387 138539 378388
rect 182357 378450 182423 378453
rect 183502 378450 183508 378452
rect 182357 378448 183508 378450
rect 182357 378392 182362 378448
rect 182418 378392 183508 378448
rect 182357 378390 183508 378392
rect 182357 378387 182423 378390
rect 183502 378388 183508 378390
rect 183572 378388 183578 378452
rect 204253 378450 204319 378453
rect 208117 378450 208183 378453
rect 241830 378450 241836 378452
rect 204253 378448 241836 378450
rect 204253 378392 204258 378448
rect 204314 378392 208122 378448
rect 208178 378392 241836 378448
rect 204253 378390 241836 378392
rect 204253 378387 204319 378390
rect 208117 378387 208183 378390
rect 241830 378388 241836 378390
rect 241900 378450 241906 378452
rect 253197 378450 253263 378453
rect 241900 378448 253263 378450
rect 241900 378392 253202 378448
rect 253258 378392 253263 378448
rect 241900 378390 253263 378392
rect 241900 378388 241906 378390
rect 253197 378387 253263 378390
rect 253381 378450 253447 378453
rect 255957 378452 256023 378453
rect 253606 378450 253612 378452
rect 253381 378448 253612 378450
rect 253381 378392 253386 378448
rect 253442 378392 253612 378448
rect 253381 378390 253612 378392
rect 253381 378387 253447 378390
rect 253606 378388 253612 378390
rect 253676 378388 253682 378452
rect 255957 378448 256004 378452
rect 256068 378450 256074 378452
rect 258030 378450 258090 378526
rect 258349 378584 258396 378588
rect 258460 378586 258466 378588
rect 258349 378528 258354 378584
rect 258349 378524 258396 378528
rect 258460 378526 258506 378586
rect 260557 378584 260604 378588
rect 260668 378586 260674 378588
rect 260557 378528 260562 378584
rect 258460 378524 258466 378526
rect 260557 378524 260604 378528
rect 260668 378526 260714 378586
rect 260925 378584 260972 378588
rect 261036 378586 261042 378588
rect 260925 378528 260930 378584
rect 260668 378524 260674 378526
rect 260925 378524 260972 378528
rect 261036 378526 261082 378586
rect 262765 378584 262812 378588
rect 262876 378586 262882 378588
rect 263542 378586 263548 378588
rect 262765 378528 262770 378584
rect 261036 378524 261042 378526
rect 262765 378524 262812 378528
rect 262876 378526 262922 378586
rect 263502 378526 263548 378586
rect 263612 378584 263659 378588
rect 263654 378528 263659 378584
rect 262876 378524 262882 378526
rect 263542 378524 263548 378526
rect 263612 378524 263659 378528
rect 258349 378523 258415 378524
rect 260557 378523 260623 378524
rect 260925 378523 260991 378524
rect 262765 378523 262831 378524
rect 263593 378523 263659 378524
rect 265893 378588 265959 378589
rect 266353 378588 266419 378589
rect 265893 378584 265940 378588
rect 266004 378586 266010 378588
rect 266302 378586 266308 378588
rect 265893 378528 265898 378584
rect 265893 378524 265940 378528
rect 266004 378526 266050 378586
rect 266262 378526 266308 378586
rect 266372 378584 266419 378588
rect 266414 378528 266419 378584
rect 266004 378524 266010 378526
rect 266302 378524 266308 378526
rect 266372 378524 266419 378528
rect 265893 378523 265959 378524
rect 266353 378523 266419 378524
rect 267549 378588 267615 378589
rect 267549 378584 267596 378588
rect 267660 378586 267666 378588
rect 268009 378586 268075 378589
rect 408677 378588 408743 378589
rect 418429 378588 418495 378589
rect 421741 378588 421807 378589
rect 268326 378586 268332 378588
rect 267549 378528 267554 378584
rect 267549 378524 267596 378528
rect 267660 378526 267706 378586
rect 268009 378584 268332 378586
rect 268009 378528 268014 378584
rect 268070 378528 268332 378584
rect 268009 378526 268332 378528
rect 267660 378524 267666 378526
rect 267549 378523 267615 378524
rect 268009 378523 268075 378526
rect 268326 378524 268332 378526
rect 268396 378524 268402 378588
rect 408677 378584 408724 378588
rect 408788 378586 408794 378588
rect 408677 378528 408682 378584
rect 408677 378524 408724 378528
rect 408788 378526 408834 378586
rect 418429 378584 418476 378588
rect 418540 378586 418546 378588
rect 418429 378528 418434 378584
rect 408788 378524 408794 378526
rect 418429 378524 418476 378528
rect 418540 378526 418586 378586
rect 421741 378584 421788 378588
rect 421852 378586 421858 378588
rect 430665 378586 430731 378589
rect 430982 378586 430988 378588
rect 421741 378528 421746 378584
rect 418540 378524 418546 378526
rect 421741 378524 421788 378528
rect 421852 378526 421898 378586
rect 430665 378584 430988 378586
rect 430665 378528 430670 378584
rect 430726 378528 430988 378584
rect 430665 378526 430988 378528
rect 421852 378524 421858 378526
rect 408677 378523 408743 378524
rect 418429 378523 418495 378524
rect 421741 378523 421807 378524
rect 430665 378523 430731 378526
rect 430982 378524 430988 378526
rect 431052 378524 431058 378588
rect 436185 378586 436251 378589
rect 436870 378586 436876 378588
rect 436185 378584 436876 378586
rect 436185 378528 436190 378584
rect 436246 378528 436876 378584
rect 436185 378526 436876 378528
rect 436185 378523 436251 378526
rect 436870 378524 436876 378526
rect 436940 378524 436946 378588
rect 274633 378450 274699 378453
rect 255957 378392 255962 378448
rect 255957 378388 256004 378392
rect 256068 378390 256114 378450
rect 258030 378448 274699 378450
rect 258030 378392 274638 378448
rect 274694 378392 274699 378448
rect 258030 378390 274699 378392
rect 256068 378388 256074 378390
rect 255957 378387 256023 378388
rect 274633 378387 274699 378390
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 100753 378316 100819 378317
rect 100702 378314 100708 378316
rect 100662 378254 100708 378314
rect 100772 378312 100819 378316
rect 100814 378256 100819 378312
rect 100702 378252 100708 378254
rect 100772 378252 100819 378256
rect 100753 378251 100819 378252
rect 182265 378314 182331 378317
rect 182817 378314 182883 378317
rect 183134 378314 183140 378316
rect 182265 378312 183140 378314
rect 182265 378256 182270 378312
rect 182326 378256 182822 378312
rect 182878 378256 183140 378312
rect 182265 378254 183140 378256
rect 182265 378251 182331 378254
rect 182817 378251 182883 378254
rect 183134 378252 183140 378254
rect 183204 378252 183210 378316
rect 205541 378314 205607 378317
rect 276013 378314 276079 378317
rect 205541 378312 276079 378314
rect 205541 378256 205546 378312
rect 205602 378256 276018 378312
rect 276074 378256 276079 378312
rect 205541 378254 276079 378256
rect 205541 378251 205607 378254
rect 276013 378251 276079 378254
rect 422569 378314 422635 378317
rect 422886 378314 422892 378316
rect 422569 378312 422892 378314
rect 422569 378256 422574 378312
rect 422630 378256 422892 378312
rect 422569 378254 422892 378256
rect 422569 378251 422635 378254
rect 422886 378252 422892 378254
rect 422956 378252 422962 378316
rect 583520 378300 584960 378390
rect 87638 378116 87644 378180
rect 87708 378178 87714 378180
rect 204713 378178 204779 378181
rect 87708 378176 204779 378178
rect 87708 378120 204718 378176
rect 204774 378120 204779 378176
rect 87708 378118 204779 378120
rect 87708 378116 87714 378118
rect 204713 378115 204779 378118
rect 210969 378178 211035 378181
rect 212441 378178 212507 378181
rect 278998 378178 279004 378180
rect 210969 378176 279004 378178
rect 210969 378120 210974 378176
rect 211030 378120 212446 378176
rect 212502 378120 279004 378176
rect 210969 378118 279004 378120
rect 210969 378115 211035 378118
rect 212441 378115 212507 378118
rect 278998 378116 279004 378118
rect 279068 378178 279074 378180
rect 280061 378178 280127 378181
rect 279068 378176 280127 378178
rect 279068 378120 280066 378176
rect 280122 378120 280127 378176
rect 279068 378118 280127 378120
rect 279068 378116 279074 378118
rect 280061 378115 280127 378118
rect 409965 378180 410031 378181
rect 416957 378180 417023 378181
rect 418153 378180 418219 378181
rect 409965 378176 410012 378180
rect 410076 378178 410082 378180
rect 409965 378120 409970 378176
rect 409965 378116 410012 378120
rect 410076 378118 410122 378178
rect 416957 378176 417004 378180
rect 417068 378178 417074 378180
rect 418102 378178 418108 378180
rect 416957 378120 416962 378176
rect 410076 378116 410082 378118
rect 416957 378116 417004 378120
rect 417068 378118 417114 378178
rect 418062 378118 418108 378178
rect 418172 378176 418219 378180
rect 418214 378120 418219 378176
rect 417068 378116 417074 378118
rect 418102 378116 418108 378118
rect 418172 378116 418219 378120
rect 409965 378115 410031 378116
rect 416957 378115 417023 378116
rect 418153 378115 418219 378116
rect 423949 378180 424015 378181
rect 423949 378176 423996 378180
rect 424060 378178 424066 378180
rect 425145 378178 425211 378181
rect 426433 378180 426499 378181
rect 425278 378178 425284 378180
rect 423949 378120 423954 378176
rect 423949 378116 423996 378120
rect 424060 378118 424106 378178
rect 425145 378176 425284 378178
rect 425145 378120 425150 378176
rect 425206 378120 425284 378176
rect 425145 378118 425284 378120
rect 424060 378116 424066 378118
rect 423949 378115 424015 378116
rect 425145 378115 425211 378118
rect 425278 378116 425284 378118
rect 425348 378116 425354 378180
rect 426382 378178 426388 378180
rect 426342 378118 426388 378178
rect 426452 378176 426499 378180
rect 426494 378120 426499 378176
rect 426382 378116 426388 378118
rect 426452 378116 426499 378120
rect 426433 378115 426499 378116
rect 428273 378178 428339 378181
rect 432229 378180 432295 378181
rect 428590 378178 428596 378180
rect 428273 378176 428596 378178
rect 428273 378120 428278 378176
rect 428334 378120 428596 378176
rect 428273 378118 428596 378120
rect 428273 378115 428339 378118
rect 428590 378116 428596 378118
rect 428660 378116 428666 378180
rect 432229 378176 432276 378180
rect 432340 378178 432346 378180
rect 435173 378178 435239 378181
rect 435766 378178 435772 378180
rect 432229 378120 432234 378176
rect 432229 378116 432276 378120
rect 432340 378118 432386 378178
rect 435173 378176 435772 378178
rect 435173 378120 435178 378176
rect 435234 378120 435772 378176
rect 435173 378118 435772 378120
rect 432340 378116 432346 378118
rect 432229 378115 432295 378116
rect 435173 378115 435239 378118
rect 435766 378116 435772 378118
rect 435836 378116 435842 378180
rect 438117 378178 438183 378181
rect 439078 378178 439084 378180
rect 438117 378176 439084 378178
rect 438117 378120 438122 378176
rect 438178 378120 439084 378176
rect 438117 378118 439084 378120
rect 438117 378115 438183 378118
rect 439078 378116 439084 378118
rect 439148 378116 439154 378180
rect 458398 378116 458404 378180
rect 458468 378116 458474 378180
rect 54477 378042 54543 378045
rect 57094 378042 57100 378044
rect 54477 378040 57100 378042
rect 54477 377984 54482 378040
rect 54538 377984 57100 378040
rect 54477 377982 57100 377984
rect 54477 377979 54543 377982
rect 57094 377980 57100 377982
rect 57164 377980 57170 378044
rect 105302 377980 105308 378044
rect 105372 378042 105378 378044
rect 105372 377982 209790 378042
rect 105372 377980 105378 377982
rect 106406 377844 106412 377908
rect 106476 377906 106482 377908
rect 205357 377906 205423 377909
rect 106476 377904 205423 377906
rect 106476 377848 205362 377904
rect 205418 377848 205423 377904
rect 106476 377846 205423 377848
rect 209730 377906 209790 377982
rect 211838 377980 211844 378044
rect 211908 378042 211914 378044
rect 212441 378042 212507 378045
rect 211908 378040 212507 378042
rect 211908 377984 212446 378040
rect 212502 377984 212507 378040
rect 211908 377982 212507 377984
rect 211908 377980 211914 377982
rect 212441 377979 212507 377982
rect 213310 377980 213316 378044
rect 213380 378042 213386 378044
rect 213821 378042 213887 378045
rect 213380 378040 213887 378042
rect 213380 377984 213826 378040
rect 213882 377984 213887 378040
rect 213380 377982 213887 377984
rect 213380 377980 213386 377982
rect 213821 377979 213887 377982
rect 215334 377980 215340 378044
rect 215404 378042 215410 378044
rect 216581 378042 216647 378045
rect 215404 378040 216647 378042
rect 215404 377984 216586 378040
rect 216642 377984 216647 378040
rect 215404 377982 216647 377984
rect 215404 377980 215410 377982
rect 216581 377979 216647 377982
rect 359774 377980 359780 378044
rect 359844 378042 359850 378044
rect 458406 378042 458466 378116
rect 359844 377982 458466 378042
rect 359844 377980 359850 377982
rect 215385 377906 215451 377909
rect 219249 377906 219315 377909
rect 209730 377904 219315 377906
rect 209730 377848 215390 377904
rect 215446 377848 219254 377904
rect 219310 377848 219315 377904
rect 209730 377846 219315 377848
rect 106476 377844 106482 377846
rect 205357 377843 205423 377846
rect 215385 377843 215451 377846
rect 219249 377843 219315 377846
rect 372654 377844 372660 377908
rect 372724 377906 372730 377908
rect 373901 377906 373967 377909
rect 438117 377906 438183 377909
rect 372724 377904 373967 377906
rect 372724 377848 373906 377904
rect 373962 377848 373967 377904
rect 372724 377846 373967 377848
rect 372724 377844 372730 377846
rect 373901 377843 373967 377846
rect 383610 377904 438183 377906
rect 383610 377848 438122 377904
rect 438178 377848 438183 377904
rect 383610 377846 438183 377848
rect 108849 377770 108915 377773
rect 205449 377770 205515 377773
rect 108849 377768 205515 377770
rect 108849 377712 108854 377768
rect 108910 377712 205454 377768
rect 205510 377712 205515 377768
rect 108849 377710 205515 377712
rect 108849 377707 108915 377710
rect 205449 377707 205515 377710
rect 373073 377770 373139 377773
rect 383610 377770 383670 377846
rect 438117 377843 438183 377846
rect 373073 377768 383670 377770
rect 373073 377712 373078 377768
rect 373134 377712 383670 377768
rect 373073 377710 383670 377712
rect 373073 377707 373139 377710
rect 369577 376954 369643 376957
rect 369761 376954 369827 376957
rect 369577 376952 369827 376954
rect 369577 376896 369582 376952
rect 369638 376896 369766 376952
rect 369822 376896 369827 376952
rect 369577 376894 369827 376896
rect 369577 376891 369643 376894
rect 369761 376891 369827 376894
rect 214230 376620 214236 376684
rect 214300 376682 214306 376684
rect 215109 376682 215175 376685
rect 214300 376680 215175 376682
rect 214300 376624 215114 376680
rect 215170 376624 215175 376680
rect 214300 376622 215175 376624
rect 214300 376620 214306 376622
rect 215109 376619 215175 376622
rect 214046 376484 214052 376548
rect 214116 376546 214122 376548
rect 215017 376546 215083 376549
rect 214116 376544 215083 376546
rect 214116 376488 215022 376544
rect 215078 376488 215083 376544
rect 214116 376486 215083 376488
rect 214116 376484 214122 376486
rect 215017 376483 215083 376486
rect 359958 375940 359964 376004
rect 360028 376002 360034 376004
rect 375189 376002 375255 376005
rect 421741 376002 421807 376005
rect 360028 376000 421807 376002
rect 360028 375944 375194 376000
rect 375250 375944 421746 376000
rect 421802 375944 421807 376000
rect 360028 375942 421807 375944
rect 360028 375940 360034 375942
rect 375189 375939 375255 375942
rect 421741 375939 421807 375942
rect 217409 375730 217475 375733
rect 217542 375730 217548 375732
rect 217409 375728 217548 375730
rect 217409 375672 217414 375728
rect 217470 375672 217548 375728
rect 217409 375670 217548 375672
rect 217409 375667 217475 375670
rect 217542 375668 217548 375670
rect 217612 375668 217618 375732
rect 376753 375324 376819 375325
rect 376702 375322 376708 375324
rect 376662 375262 376708 375322
rect 376772 375320 376819 375324
rect 376814 375264 376819 375320
rect 376702 375260 376708 375262
rect 376772 375260 376819 375264
rect 377806 375260 377812 375324
rect 377876 375322 377882 375324
rect 381261 375322 381327 375325
rect 377876 375320 381327 375322
rect 377876 375264 381266 375320
rect 381322 375264 381327 375320
rect 377876 375262 381327 375264
rect 377876 375260 377882 375262
rect 376753 375259 376819 375260
rect 381261 375259 381327 375262
rect 207289 374642 207355 374645
rect 216673 374644 216739 374645
rect 216622 374642 216628 374644
rect 207289 374640 216628 374642
rect 216692 374640 216739 374644
rect 207289 374584 207294 374640
rect 207350 374584 216628 374640
rect 216734 374584 216739 374640
rect 207289 374582 216628 374584
rect 207289 374579 207355 374582
rect 216622 374580 216628 374582
rect 216692 374580 216739 374584
rect 216673 374579 216739 374580
rect 381261 374642 381327 374645
rect 435173 374642 435239 374645
rect 381261 374640 435239 374642
rect 381261 374584 381266 374640
rect 381322 374584 435178 374640
rect 435234 374584 435239 374640
rect 381261 374582 435239 374584
rect 381261 374579 381327 374582
rect 435173 374579 435239 374582
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect 178585 358868 178651 358869
rect 179689 358868 179755 358869
rect 190913 358868 190979 358869
rect 338481 358868 338547 358869
rect 339769 358868 339835 358869
rect 178534 358866 178540 358868
rect 178494 358806 178540 358866
rect 178604 358864 178651 358868
rect 179638 358866 179644 358868
rect 178646 358808 178651 358864
rect 178534 358804 178540 358806
rect 178604 358804 178651 358808
rect 179598 358806 179644 358866
rect 179708 358864 179755 358868
rect 190862 358866 190868 358868
rect 179750 358808 179755 358864
rect 179638 358804 179644 358806
rect 179708 358804 179755 358808
rect 190822 358806 190868 358866
rect 190932 358864 190979 358868
rect 338430 358866 338436 358868
rect 190974 358808 190979 358864
rect 190862 358804 190868 358806
rect 190932 358804 190979 358808
rect 338390 358806 338436 358866
rect 338500 358864 338547 358868
rect 339718 358866 339724 358868
rect 338542 358808 338547 358864
rect 338430 358804 338436 358806
rect 338500 358804 338547 358808
rect 339678 358806 339724 358866
rect 339788 358864 339835 358868
rect 339830 358808 339835 358864
rect 339718 358804 339724 358806
rect 339788 358804 339835 358808
rect 350942 358804 350948 358868
rect 351012 358866 351018 358868
rect 351729 358866 351795 358869
rect 351012 358864 351795 358866
rect 351012 358808 351734 358864
rect 351790 358808 351795 358864
rect 351012 358806 351795 358808
rect 351012 358804 351018 358806
rect 178585 358803 178651 358804
rect 179689 358803 179755 358804
rect 190913 358803 190979 358804
rect 338481 358803 338547 358804
rect 339769 358803 339835 358804
rect 351729 358803 351795 358806
rect 498510 358804 498516 358868
rect 498580 358866 498586 358868
rect 498837 358866 498903 358869
rect 498580 358864 498903 358866
rect 498580 358808 498842 358864
rect 498898 358808 498903 358864
rect 498580 358806 498903 358808
rect 498580 358804 498586 358806
rect 498837 358803 498903 358806
rect 499798 358804 499804 358868
rect 499868 358866 499874 358868
rect 500769 358866 500835 358869
rect 510889 358868 510955 358869
rect 510838 358866 510844 358868
rect 499868 358864 500835 358866
rect 499868 358808 500774 358864
rect 500830 358808 500835 358864
rect 499868 358806 500835 358808
rect 510798 358806 510844 358866
rect 510908 358864 510955 358868
rect 510950 358808 510955 358864
rect 499868 358804 499874 358806
rect 500769 358803 500835 358806
rect 510838 358804 510844 358806
rect 510908 358804 510955 358808
rect 510889 358803 510955 358804
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 57462 357308 57468 357372
rect 57532 357370 57538 357372
rect 59353 357370 59419 357373
rect 57532 357368 59419 357370
rect 57532 357312 59358 357368
rect 59414 357312 59419 357368
rect 57532 357310 59419 357312
rect 57532 357308 57538 357310
rect 59353 357307 59419 357310
rect 196558 353154 196618 353190
rect 198825 353154 198891 353157
rect 196558 353152 198891 353154
rect 196558 353096 198830 353152
rect 198886 353096 198891 353152
rect 196558 353094 198891 353096
rect 356562 353154 356622 353190
rect 359457 353154 359523 353157
rect 356562 353152 359523 353154
rect 356562 353096 359462 353152
rect 359518 353096 359523 353152
rect 356562 353094 359523 353096
rect 198825 353091 198891 353094
rect 359457 353091 359523 353094
rect 516558 352882 516618 353190
rect 519261 352882 519327 352885
rect 519445 352882 519511 352885
rect 516558 352880 519511 352882
rect 516558 352824 519266 352880
rect 519322 352824 519450 352880
rect 519506 352824 519511 352880
rect 516558 352822 519511 352824
rect 519261 352819 519327 352822
rect 519445 352819 519511 352822
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580257 325274 580323 325277
rect 583520 325274 584960 325364
rect 580257 325272 584960 325274
rect 580257 325216 580262 325272
rect 580318 325216 584960 325272
rect 580257 325214 584960 325216
rect 580257 325211 580323 325214
rect 583520 325124 584960 325214
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect 56685 311130 56751 311133
rect 57881 311130 57947 311133
rect 56685 311128 60062 311130
rect 56685 311072 56690 311128
rect 56746 311072 57886 311128
rect 57942 311072 60062 311128
rect 56685 311070 60062 311072
rect 56685 311067 56751 311070
rect 57881 311067 57947 311070
rect 60002 310894 60062 311070
rect 219390 310864 220064 310924
rect 379838 310864 380052 310924
rect 217501 310858 217567 310861
rect 217777 310858 217843 310861
rect 219390 310858 219450 310864
rect 217501 310856 219450 310858
rect 217501 310800 217506 310856
rect 217562 310800 217782 310856
rect 217838 310800 219450 310856
rect 217501 310798 219450 310800
rect 376937 310858 377003 310861
rect 377581 310858 377647 310861
rect 379838 310858 379898 310864
rect 376937 310856 379898 310858
rect 376937 310800 376942 310856
rect 376998 310800 377586 310856
rect 377642 310800 379898 310856
rect 376937 310798 379898 310800
rect 217501 310795 217567 310798
rect 217777 310795 217843 310798
rect 376937 310795 377003 310798
rect 377581 310795 377647 310798
rect 57145 310450 57211 310453
rect 57697 310450 57763 310453
rect 57145 310448 60062 310450
rect 57145 310392 57150 310448
rect 57206 310392 57702 310448
rect 57758 310392 60062 310448
rect 57145 310390 60062 310392
rect 57145 310387 57211 310390
rect 57697 310387 57763 310390
rect 60002 309942 60062 310390
rect 217409 310042 217475 310045
rect 217869 310042 217935 310045
rect 378041 310042 378107 310045
rect 217409 310040 219450 310042
rect 217409 309984 217414 310040
rect 217470 309984 217874 310040
rect 217930 309984 219450 310040
rect 217409 309982 219450 309984
rect 217409 309979 217475 309982
rect 217869 309979 217935 309982
rect 219390 309972 219450 309982
rect 378041 310040 379898 310042
rect 378041 309984 378046 310040
rect 378102 309984 379898 310040
rect 378041 309982 379898 309984
rect 378041 309979 378107 309982
rect 379838 309972 379898 309982
rect 219390 309912 220064 309972
rect 379838 309912 380052 309972
rect 57605 307866 57671 307869
rect 217593 307866 217659 307869
rect 377765 307866 377831 307869
rect 57605 307864 59922 307866
rect 57605 307808 57610 307864
rect 57666 307808 59922 307864
rect 57605 307806 59922 307808
rect 57605 307803 57671 307806
rect 59862 307796 59922 307806
rect 217593 307864 219450 307866
rect 217593 307808 217598 307864
rect 217654 307808 219450 307864
rect 217593 307806 219450 307808
rect 217593 307803 217659 307806
rect 219390 307796 219450 307806
rect 377765 307864 379898 307866
rect 377765 307808 377770 307864
rect 377826 307808 379898 307864
rect 377765 307806 379898 307808
rect 377765 307803 377831 307806
rect 379838 307796 379898 307806
rect 59862 307736 60032 307796
rect 219390 307736 220064 307796
rect 379838 307736 380052 307796
rect 216949 307730 217015 307733
rect 217685 307730 217751 307733
rect 216949 307728 217751 307730
rect 216949 307672 216954 307728
rect 217010 307672 217690 307728
rect 217746 307672 217751 307728
rect 216949 307670 217751 307672
rect 216949 307667 217015 307670
rect 217685 307667 217751 307670
rect 57329 306778 57395 306781
rect 60002 306778 60062 306814
rect 219390 306784 220064 306844
rect 379838 306784 380052 306844
rect 57329 306776 60062 306778
rect 57329 306720 57334 306776
rect 57390 306720 60062 306776
rect 57329 306718 60062 306720
rect 217685 306778 217751 306781
rect 219390 306778 219450 306784
rect 217685 306776 219450 306778
rect 217685 306720 217690 306776
rect 217746 306720 219450 306776
rect 217685 306718 219450 306720
rect 377673 306778 377739 306781
rect 379838 306778 379898 306784
rect 377673 306776 379898 306778
rect 377673 306720 377678 306776
rect 377734 306720 379898 306776
rect 377673 306718 379898 306720
rect 57329 306715 57395 306718
rect 217685 306715 217751 306718
rect 377673 306715 377739 306718
rect -960 306234 480 306324
rect -960 306174 674 306234
rect -960 306098 480 306174
rect 614 306098 674 306174
rect -960 306084 674 306098
rect 246 306038 674 306084
rect 246 305554 306 306038
rect 246 305494 6930 305554
rect 6870 305010 6930 305494
rect 53046 305010 53052 305012
rect 6870 304950 53052 305010
rect 53046 304948 53052 304950
rect 53116 304948 53122 305012
rect 57513 305010 57579 305013
rect 60002 305010 60062 305046
rect 219390 305016 220064 305076
rect 379838 305016 380052 305076
rect 57513 305008 60062 305010
rect 57513 304952 57518 305008
rect 57574 304952 60062 305008
rect 57513 304950 60062 304952
rect 217041 305010 217107 305013
rect 217869 305010 217935 305013
rect 219390 305010 219450 305016
rect 217041 305008 219450 305010
rect 217041 304952 217046 305008
rect 217102 304952 217874 305008
rect 217930 304952 219450 305008
rect 217041 304950 219450 304952
rect 377489 305010 377555 305013
rect 379838 305010 379898 305016
rect 377489 305008 379898 305010
rect 377489 304952 377494 305008
rect 377550 304952 379898 305008
rect 377489 304950 379898 304952
rect 57513 304947 57579 304950
rect 217041 304947 217107 304950
rect 217869 304947 217935 304950
rect 377489 304947 377555 304950
rect 57421 303922 57487 303925
rect 60002 303922 60062 303958
rect 219390 303928 220064 303988
rect 379838 303928 380052 303988
rect 57421 303920 60062 303922
rect 57421 303864 57426 303920
rect 57482 303864 60062 303920
rect 57421 303862 60062 303864
rect 217133 303922 217199 303925
rect 217777 303922 217843 303925
rect 219390 303922 219450 303928
rect 217133 303920 219450 303922
rect 217133 303864 217138 303920
rect 217194 303864 217782 303920
rect 217838 303864 219450 303920
rect 217133 303862 219450 303864
rect 377857 303922 377923 303925
rect 379838 303922 379898 303928
rect 377857 303920 379898 303922
rect 377857 303864 377862 303920
rect 377918 303864 379898 303920
rect 377857 303862 379898 303864
rect 57421 303859 57487 303862
rect 217133 303859 217199 303862
rect 217777 303859 217843 303862
rect 377857 303859 377923 303862
rect 377673 303650 377739 303653
rect 377857 303650 377923 303653
rect 377673 303648 377923 303650
rect 377673 303592 377678 303648
rect 377734 303592 377862 303648
rect 377918 303592 377923 303648
rect 377673 303590 377923 303592
rect 377673 303587 377739 303590
rect 377857 303587 377923 303590
rect 56961 301610 57027 301613
rect 60002 301610 60062 302190
rect 219390 302160 220064 302220
rect 379838 302160 380052 302220
rect 217041 302154 217107 302157
rect 217317 302154 217383 302157
rect 219390 302154 219450 302160
rect 217041 302152 219450 302154
rect 217041 302096 217046 302152
rect 217102 302096 217322 302152
rect 217378 302096 219450 302152
rect 217041 302094 219450 302096
rect 377305 302154 377371 302157
rect 377949 302154 378015 302157
rect 379838 302154 379898 302160
rect 377305 302152 379898 302154
rect 377305 302096 377310 302152
rect 377366 302096 377954 302152
rect 378010 302096 379898 302152
rect 377305 302094 379898 302096
rect 217041 302091 217107 302094
rect 217317 302091 217383 302094
rect 377305 302091 377371 302094
rect 377949 302091 378015 302094
rect 56961 301608 60062 301610
rect 56961 301552 56966 301608
rect 57022 301552 60062 301608
rect 56961 301550 60062 301552
rect 56961 301547 57027 301550
rect 583520 298604 584960 298844
rect 519353 293858 519419 293861
rect 516558 293856 519419 293858
rect 516558 293800 519358 293856
rect 519414 293800 519419 293856
rect 516558 293798 519419 293800
rect 516558 293350 516618 293798
rect 519353 293795 519419 293798
rect -960 293028 480 293268
rect 196558 292770 196618 293350
rect 199193 292770 199259 292773
rect 199561 292770 199627 292773
rect 196558 292768 199627 292770
rect 196558 292712 199198 292768
rect 199254 292712 199566 292768
rect 199622 292712 199627 292768
rect 196558 292710 199627 292712
rect 356562 292770 356622 293350
rect 359365 292770 359431 292773
rect 359549 292770 359615 292773
rect 356562 292768 359615 292770
rect 356562 292712 359370 292768
rect 359426 292712 359554 292768
rect 359610 292712 359615 292768
rect 356562 292710 359615 292712
rect 199193 292707 199259 292710
rect 199561 292707 199627 292710
rect 359365 292707 359431 292710
rect 359549 292707 359615 292710
rect 359641 291818 359707 291821
rect 356562 291816 359707 291818
rect 356562 291760 359646 291816
rect 359702 291760 359707 291816
rect 356562 291758 359707 291760
rect 356562 291718 356622 291758
rect 359641 291755 359707 291758
rect 196558 291682 196618 291718
rect 198733 291682 198799 291685
rect 199377 291682 199443 291685
rect 196558 291680 199443 291682
rect 196558 291624 198738 291680
rect 198794 291624 199382 291680
rect 199438 291624 199443 291680
rect 196558 291622 199443 291624
rect 516558 291682 516618 291718
rect 518893 291682 518959 291685
rect 516558 291680 518959 291682
rect 516558 291624 518898 291680
rect 518954 291624 518959 291680
rect 516558 291622 518959 291624
rect 198733 291619 198799 291622
rect 199377 291619 199443 291622
rect 518893 291619 518959 291622
rect 198917 291002 198983 291005
rect 199469 291002 199535 291005
rect 358905 291002 358971 291005
rect 196558 291000 199535 291002
rect 196558 290944 198922 291000
rect 198978 290944 199474 291000
rect 199530 290944 199535 291000
rect 196558 290942 199535 290944
rect 196558 290358 196618 290942
rect 198917 290939 198983 290942
rect 199469 290939 199535 290942
rect 356562 291000 358971 291002
rect 356562 290944 358910 291000
rect 358966 290944 358971 291000
rect 356562 290942 358971 290944
rect 356562 290358 356622 290942
rect 358905 290939 358971 290942
rect 516558 290322 516618 290358
rect 519537 290322 519603 290325
rect 516558 290320 519603 290322
rect 516558 290264 519542 290320
rect 519598 290264 519603 290320
rect 516558 290262 519603 290264
rect 519537 290259 519603 290262
rect 199101 289778 199167 289781
rect 199653 289778 199719 289781
rect 199101 289776 199719 289778
rect 199101 289720 199106 289776
rect 199162 289720 199658 289776
rect 199714 289720 199719 289776
rect 199101 289718 199719 289720
rect 199101 289715 199167 289718
rect 199653 289715 199719 289718
rect 196558 288826 196618 288862
rect 199101 288826 199167 288829
rect 196558 288824 199167 288826
rect 196558 288768 199106 288824
rect 199162 288768 199167 288824
rect 196558 288766 199167 288768
rect 356562 288826 356622 288862
rect 359181 288826 359247 288829
rect 356562 288824 359247 288826
rect 356562 288768 359186 288824
rect 359242 288768 359247 288824
rect 356562 288766 359247 288768
rect 516558 288826 516618 288862
rect 519077 288826 519143 288829
rect 520181 288826 520247 288829
rect 516558 288824 520247 288826
rect 516558 288768 519082 288824
rect 519138 288768 520186 288824
rect 520242 288768 520247 288824
rect 516558 288766 520247 288768
rect 199101 288763 199167 288766
rect 359181 288763 359247 288766
rect 519077 288763 519143 288766
rect 520181 288763 520247 288766
rect 199009 288418 199075 288421
rect 199745 288418 199811 288421
rect 199009 288416 199811 288418
rect 199009 288360 199014 288416
rect 199070 288360 199750 288416
rect 199806 288360 199811 288416
rect 199009 288358 199811 288360
rect 199009 288355 199075 288358
rect 199745 288355 199811 288358
rect 359273 288418 359339 288421
rect 359549 288418 359615 288421
rect 359273 288416 359615 288418
rect 359273 288360 359278 288416
rect 359334 288360 359554 288416
rect 359610 288360 359615 288416
rect 359273 288358 359615 288360
rect 359273 288355 359339 288358
rect 359549 288355 359615 288358
rect 196558 287602 196618 287638
rect 199009 287602 199075 287605
rect 196558 287600 199075 287602
rect 196558 287544 199014 287600
rect 199070 287544 199075 287600
rect 196558 287542 199075 287544
rect 356562 287602 356622 287638
rect 359549 287602 359615 287605
rect 356562 287600 359615 287602
rect 356562 287544 359554 287600
rect 359610 287544 359615 287600
rect 356562 287542 359615 287544
rect 516558 287602 516618 287638
rect 519169 287602 519235 287605
rect 516558 287600 519235 287602
rect 516558 287544 519174 287600
rect 519230 287544 519235 287600
rect 516558 287542 519235 287544
rect 199009 287539 199075 287542
rect 359549 287539 359615 287542
rect 519169 287539 519235 287542
rect 583520 285276 584960 285516
rect 58801 284202 58867 284205
rect 58801 284200 60062 284202
rect 58801 284144 58806 284200
rect 58862 284144 60062 284200
rect 58801 284142 60062 284144
rect 58801 284139 58867 284142
rect 60002 283966 60062 284142
rect 216673 284066 216739 284069
rect 376937 284066 377003 284069
rect 216673 284064 219450 284066
rect 216673 284008 216678 284064
rect 216734 284008 219450 284064
rect 216673 284006 219450 284008
rect 216673 284003 216739 284006
rect 219390 283996 219450 284006
rect 376937 284064 379530 284066
rect 376937 284008 376942 284064
rect 376998 284008 379530 284064
rect 376937 284006 379530 284008
rect 376937 284003 377003 284006
rect 379470 283996 379530 284006
rect 219390 283936 220064 283996
rect 379470 283936 380052 283996
rect 216673 282434 216739 282437
rect 216673 282432 219450 282434
rect 216673 282376 216678 282432
rect 216734 282376 219450 282432
rect 216673 282374 219450 282376
rect 216673 282371 216739 282374
rect 219390 282364 219450 282374
rect 59494 282304 60032 282364
rect 219390 282304 220064 282364
rect 379470 282304 380052 282364
rect 57513 282298 57579 282301
rect 59494 282298 59554 282304
rect 57513 282296 59554 282298
rect 57513 282240 57518 282296
rect 57574 282240 59554 282296
rect 57513 282238 59554 282240
rect 376937 282298 377003 282301
rect 379470 282298 379530 282304
rect 376937 282296 379530 282298
rect 376937 282240 376942 282296
rect 376998 282240 379530 282296
rect 376937 282238 379530 282240
rect 57513 282235 57579 282238
rect 376937 282235 377003 282238
rect 216765 282162 216831 282165
rect 376753 282162 376819 282165
rect 216765 282160 219450 282162
rect 216765 282104 216770 282160
rect 216826 282104 219450 282160
rect 216765 282102 219450 282104
rect 216765 282099 216831 282102
rect 219390 282092 219450 282102
rect 376753 282160 379530 282162
rect 376753 282104 376758 282160
rect 376814 282104 379530 282160
rect 376753 282102 379530 282104
rect 376753 282099 376819 282102
rect 379470 282092 379530 282102
rect 58709 282026 58775 282029
rect 60002 282026 60062 282062
rect 219390 282032 220064 282092
rect 379470 282032 380052 282092
rect 58709 282024 60062 282026
rect 58709 281968 58714 282024
rect 58770 281968 60062 282024
rect 58709 281966 60062 281968
rect 58709 281963 58775 281966
rect -960 279972 480 280212
rect 95969 273868 96035 273869
rect 95904 273804 95910 273868
rect 95974 273866 96035 273868
rect 95974 273864 96066 273866
rect 96030 273808 96066 273864
rect 95974 273806 96066 273808
rect 95974 273804 96035 273806
rect 95969 273803 96035 273804
rect 131021 273732 131087 273733
rect 130992 273668 130998 273732
rect 131062 273730 131087 273732
rect 145925 273732 145991 273733
rect 440877 273732 440943 273733
rect 145925 273730 145958 273732
rect 131062 273728 131154 273730
rect 131082 273672 131154 273728
rect 131062 273670 131154 273672
rect 145866 273728 145958 273730
rect 145866 273672 145930 273728
rect 145866 273670 145958 273672
rect 131062 273668 131087 273670
rect 131021 273667 131087 273668
rect 145925 273668 145958 273670
rect 146022 273668 146028 273732
rect 440877 273730 440934 273732
rect 440842 273728 440934 273730
rect 440842 273672 440882 273728
rect 440842 273670 440934 273672
rect 440877 273668 440934 273670
rect 440998 273668 441004 273732
rect 145925 273667 145991 273668
rect 440877 273667 440943 273668
rect 133413 273596 133479 273597
rect 135897 273596 135963 273597
rect 138473 273596 138539 273597
rect 140865 273596 140931 273597
rect 250713 273596 250779 273597
rect 272241 273596 272307 273597
rect 133413 273594 133446 273596
rect 133354 273592 133446 273594
rect 133354 273536 133418 273592
rect 133354 273534 133446 273536
rect 133413 273532 133446 273534
rect 133510 273532 133516 273596
rect 135888 273532 135894 273596
rect 135958 273594 135964 273596
rect 138472 273594 138478 273596
rect 135958 273534 136050 273594
rect 138386 273534 138478 273594
rect 135958 273532 135964 273534
rect 138472 273532 138478 273534
rect 138542 273532 138548 273596
rect 140865 273594 140926 273596
rect 140834 273592 140926 273594
rect 140834 273536 140870 273592
rect 140834 273534 140926 273536
rect 140865 273532 140926 273534
rect 140990 273532 140996 273596
rect 250713 273594 250742 273596
rect 250650 273592 250742 273594
rect 250650 273536 250718 273592
rect 250650 273534 250742 273536
rect 250713 273532 250742 273534
rect 250806 273532 250812 273596
rect 272224 273532 272230 273596
rect 272294 273594 272307 273596
rect 280889 273596 280955 273597
rect 416037 273596 416103 273597
rect 427629 273596 427695 273597
rect 433333 273596 433399 273597
rect 280889 273594 280934 273596
rect 272294 273592 272386 273594
rect 272302 273536 272386 273592
rect 272294 273534 272386 273536
rect 280842 273592 280934 273594
rect 280842 273536 280894 273592
rect 280842 273534 280934 273536
rect 272294 273532 272307 273534
rect 133413 273531 133479 273532
rect 135897 273531 135963 273532
rect 138473 273531 138539 273532
rect 140865 273531 140931 273532
rect 250713 273531 250779 273532
rect 272241 273531 272307 273532
rect 280889 273532 280934 273534
rect 280998 273532 281004 273596
rect 416037 273594 416046 273596
rect 415954 273592 416046 273594
rect 415954 273536 416042 273592
rect 415954 273534 416046 273536
rect 416037 273532 416046 273534
rect 416110 273532 416116 273596
rect 427600 273532 427606 273596
rect 427670 273594 427695 273596
rect 427670 273592 427762 273594
rect 427690 273536 427762 273592
rect 427670 273534 427762 273536
rect 427670 273532 427695 273534
rect 433312 273532 433318 273596
rect 433382 273594 433399 273596
rect 433382 273592 433474 273594
rect 433394 273536 433474 273592
rect 433382 273534 433474 273536
rect 433382 273532 433399 273534
rect 280889 273531 280955 273532
rect 416037 273531 416103 273532
rect 427629 273531 427695 273532
rect 433333 273531 433399 273532
rect 273253 273460 273319 273461
rect 273253 273458 273300 273460
rect 273208 273456 273300 273458
rect 273208 273400 273258 273456
rect 273208 273398 273300 273400
rect 273253 273396 273300 273398
rect 273364 273396 273370 273460
rect 273253 273395 273319 273396
rect 371785 273322 371851 273325
rect 376886 273322 376892 273324
rect 371785 273320 376892 273322
rect 371785 273264 371790 273320
rect 371846 273264 376892 273320
rect 371785 273262 376892 273264
rect 371785 273259 371851 273262
rect 376886 273260 376892 273262
rect 376956 273322 376962 273324
rect 377990 273322 377996 273324
rect 376956 273262 377996 273322
rect 376956 273260 376962 273262
rect 377990 273260 377996 273262
rect 378060 273260 378066 273324
rect 378358 273260 378364 273324
rect 378428 273322 378434 273324
rect 379421 273322 379487 273325
rect 430941 273324 431007 273325
rect 430941 273322 430988 273324
rect 378428 273320 379487 273322
rect 378428 273264 379426 273320
rect 379482 273264 379487 273320
rect 378428 273262 379487 273264
rect 430896 273320 430988 273322
rect 430896 273264 430946 273320
rect 430896 273262 430988 273264
rect 378428 273260 378434 273262
rect 379421 273259 379487 273262
rect 430941 273260 430988 273262
rect 431052 273260 431058 273324
rect 430941 273259 431007 273260
rect 77109 273188 77175 273189
rect 88333 273188 88399 273189
rect 90725 273188 90791 273189
rect 93669 273188 93735 273189
rect 98085 273188 98151 273189
rect 77109 273186 77156 273188
rect 77064 273184 77156 273186
rect 77064 273128 77114 273184
rect 77064 273126 77156 273128
rect 77109 273124 77156 273126
rect 77220 273124 77226 273188
rect 88333 273186 88380 273188
rect 88288 273184 88380 273186
rect 88288 273128 88338 273184
rect 88288 273126 88380 273128
rect 88333 273124 88380 273126
rect 88444 273124 88450 273188
rect 90725 273186 90772 273188
rect 90680 273184 90772 273186
rect 90680 273128 90730 273184
rect 90680 273126 90772 273128
rect 90725 273124 90772 273126
rect 90836 273124 90842 273188
rect 93669 273186 93716 273188
rect 93624 273184 93716 273186
rect 93624 273128 93674 273184
rect 93624 273126 93716 273128
rect 93669 273124 93716 273126
rect 93780 273124 93786 273188
rect 98085 273186 98132 273188
rect 98040 273184 98132 273186
rect 98040 273128 98090 273184
rect 98040 273126 98132 273128
rect 98085 273124 98132 273126
rect 98196 273124 98202 273188
rect 101806 273124 101812 273188
rect 101876 273186 101882 273188
rect 196750 273186 196756 273188
rect 101876 273126 196756 273186
rect 101876 273124 101882 273126
rect 196750 273124 196756 273126
rect 196820 273124 196826 273188
rect 198038 273124 198044 273188
rect 198108 273186 198114 273188
rect 318374 273186 318380 273188
rect 198108 273126 318380 273186
rect 198108 273124 198114 273126
rect 318374 273124 318380 273126
rect 318444 273124 318450 273188
rect 358537 273186 358603 273189
rect 485998 273186 486004 273188
rect 358537 273184 486004 273186
rect 358537 273128 358542 273184
rect 358598 273128 486004 273184
rect 358537 273126 486004 273128
rect 77109 273123 77175 273124
rect 88333 273123 88399 273124
rect 90725 273123 90791 273124
rect 93669 273123 93735 273124
rect 98085 273123 98151 273124
rect 358537 273123 358603 273126
rect 485998 273124 486004 273126
rect 486068 273124 486074 273188
rect 50337 273050 50403 273053
rect 112110 273050 112116 273052
rect 50337 273048 112116 273050
rect 50337 272992 50342 273048
rect 50398 272992 112116 273048
rect 50337 272990 112116 272992
rect 50337 272987 50403 272990
rect 112110 272988 112116 272990
rect 112180 272988 112186 273052
rect 198222 272988 198228 273052
rect 198292 273050 198298 273052
rect 311014 273050 311020 273052
rect 198292 272990 311020 273050
rect 198292 272988 198298 272990
rect 311014 272988 311020 272990
rect 311084 272988 311090 273052
rect 365529 273050 365595 273053
rect 483238 273050 483244 273052
rect 365529 273048 483244 273050
rect 365529 272992 365534 273048
rect 365590 272992 483244 273048
rect 365529 272990 483244 272992
rect 365529 272987 365595 272990
rect 483238 272988 483244 272990
rect 483308 272988 483314 273052
rect 50521 272914 50587 272917
rect 54569 272914 54635 272917
rect 98453 272916 98519 272917
rect 99373 272916 99439 272917
rect 423397 272916 423463 272917
rect 423765 272916 423831 272917
rect 426433 272916 426499 272917
rect 98453 272914 98500 272916
rect 50521 272912 97274 272914
rect 50521 272856 50526 272912
rect 50582 272856 54574 272912
rect 54630 272856 97274 272912
rect 50521 272854 97274 272856
rect 98408 272912 98500 272914
rect 98408 272856 98458 272912
rect 98408 272854 98500 272856
rect 50521 272851 50587 272854
rect 54569 272851 54635 272854
rect 51625 272778 51691 272781
rect 95693 272778 95759 272781
rect 95877 272780 95943 272781
rect 95877 272778 95924 272780
rect 51625 272776 95759 272778
rect 51625 272720 51630 272776
rect 51686 272720 95698 272776
rect 95754 272720 95759 272776
rect 51625 272718 95759 272720
rect 95832 272776 95924 272778
rect 95832 272720 95882 272776
rect 95832 272718 95924 272720
rect 51625 272715 51691 272718
rect 95693 272715 95759 272718
rect 95877 272716 95924 272718
rect 95988 272716 95994 272780
rect 97214 272778 97274 272854
rect 98453 272852 98500 272854
rect 98564 272852 98570 272916
rect 99373 272914 99420 272916
rect 99328 272912 99420 272914
rect 99328 272856 99378 272912
rect 99328 272854 99420 272856
rect 99373 272852 99420 272854
rect 99484 272852 99490 272916
rect 199326 272852 199332 272916
rect 199396 272914 199402 272916
rect 305862 272914 305868 272916
rect 199396 272854 305868 272914
rect 199396 272852 199402 272854
rect 305862 272852 305868 272854
rect 305932 272852 305938 272916
rect 359406 272852 359412 272916
rect 359476 272914 359482 272916
rect 423397 272914 423444 272916
rect 359476 272854 423138 272914
rect 423352 272912 423444 272914
rect 423352 272856 423402 272912
rect 423352 272854 423444 272856
rect 359476 272852 359482 272854
rect 98453 272851 98519 272852
rect 99373 272851 99439 272852
rect 283373 272780 283439 272781
rect 288157 272780 288223 272781
rect 290917 272780 290983 272781
rect 295885 272780 295951 272781
rect 100702 272778 100708 272780
rect 97214 272718 100708 272778
rect 100702 272716 100708 272718
rect 100772 272716 100778 272780
rect 199510 272716 199516 272780
rect 199580 272778 199586 272780
rect 283373 272778 283420 272780
rect 199580 272718 281642 272778
rect 283328 272776 283420 272778
rect 283328 272720 283378 272776
rect 283328 272718 283420 272720
rect 199580 272716 199586 272718
rect 95877 272715 95943 272716
rect 59629 272642 59695 272645
rect 117998 272642 118004 272644
rect 59629 272640 118004 272642
rect 59629 272584 59634 272640
rect 59690 272584 118004 272640
rect 59629 272582 118004 272584
rect 59629 272579 59695 272582
rect 117998 272580 118004 272582
rect 118068 272580 118074 272644
rect 196566 272580 196572 272644
rect 196636 272642 196642 272644
rect 278446 272642 278452 272644
rect 196636 272582 278452 272642
rect 196636 272580 196642 272582
rect 278446 272580 278452 272582
rect 278516 272580 278522 272644
rect 281582 272642 281642 272718
rect 283373 272716 283420 272718
rect 283484 272716 283490 272780
rect 288157 272778 288204 272780
rect 288112 272776 288204 272778
rect 288112 272720 288162 272776
rect 288112 272718 288204 272720
rect 288157 272716 288204 272718
rect 288268 272716 288274 272780
rect 290917 272778 290964 272780
rect 290872 272776 290964 272778
rect 290872 272720 290922 272776
rect 290872 272718 290964 272720
rect 290917 272716 290964 272718
rect 291028 272716 291034 272780
rect 295885 272778 295932 272780
rect 295840 272776 295932 272778
rect 295840 272720 295890 272776
rect 295840 272718 295932 272720
rect 295885 272716 295932 272718
rect 295996 272716 296002 272780
rect 377990 272716 377996 272780
rect 378060 272778 378066 272780
rect 422886 272778 422892 272780
rect 378060 272718 422892 272778
rect 378060 272716 378066 272718
rect 422886 272716 422892 272718
rect 422956 272716 422962 272780
rect 423078 272778 423138 272854
rect 423397 272852 423444 272854
rect 423508 272852 423514 272916
rect 423765 272914 423812 272916
rect 423720 272912 423812 272914
rect 423720 272856 423770 272912
rect 423720 272854 423812 272856
rect 423765 272852 423812 272854
rect 423876 272852 423882 272916
rect 426382 272852 426388 272916
rect 426452 272914 426499 272916
rect 428181 272916 428247 272917
rect 468477 272916 468543 272917
rect 470869 272916 470935 272917
rect 428181 272914 428228 272916
rect 426452 272912 426544 272914
rect 426494 272856 426544 272912
rect 426452 272854 426544 272856
rect 428136 272912 428228 272914
rect 428136 272856 428186 272912
rect 428136 272854 428228 272856
rect 426452 272852 426499 272854
rect 423397 272851 423463 272852
rect 423765 272851 423831 272852
rect 426433 272851 426499 272852
rect 428181 272852 428228 272854
rect 428292 272852 428298 272916
rect 468477 272914 468524 272916
rect 468432 272912 468524 272914
rect 468432 272856 468482 272912
rect 468432 272854 468524 272856
rect 468477 272852 468524 272854
rect 468588 272852 468594 272916
rect 470869 272914 470916 272916
rect 470824 272912 470916 272914
rect 470824 272856 470874 272912
rect 470824 272854 470916 272856
rect 470869 272852 470916 272854
rect 470980 272852 470986 272916
rect 428181 272851 428247 272852
rect 468477 272851 468543 272852
rect 470869 272851 470935 272852
rect 478413 272780 478479 272781
rect 480805 272780 480871 272781
rect 426014 272778 426020 272780
rect 423078 272718 426020 272778
rect 426014 272716 426020 272718
rect 426084 272716 426090 272780
rect 478413 272778 478460 272780
rect 478368 272776 478460 272778
rect 478368 272720 478418 272776
rect 478368 272718 478460 272720
rect 478413 272716 478460 272718
rect 478524 272716 478530 272780
rect 480805 272778 480852 272780
rect 480760 272776 480852 272778
rect 480760 272720 480810 272776
rect 480760 272718 480852 272720
rect 480805 272716 480852 272718
rect 480916 272716 480922 272780
rect 283373 272715 283439 272716
rect 288157 272715 288223 272716
rect 290917 272715 290983 272716
rect 295885 272715 295951 272716
rect 478413 272715 478479 272716
rect 480805 272715 480871 272716
rect 298461 272644 298527 272645
rect 300853 272644 300919 272645
rect 473445 272644 473511 272645
rect 475837 272644 475903 272645
rect 285990 272642 285996 272644
rect 281582 272582 285996 272642
rect 285990 272580 285996 272582
rect 286060 272580 286066 272644
rect 298461 272642 298508 272644
rect 298416 272640 298508 272642
rect 298416 272584 298466 272640
rect 298416 272582 298508 272584
rect 298461 272580 298508 272582
rect 298572 272580 298578 272644
rect 300853 272642 300900 272644
rect 300808 272640 300900 272642
rect 300808 272584 300858 272640
rect 300808 272582 300900 272584
rect 300853 272580 300900 272582
rect 300964 272580 300970 272644
rect 473445 272642 473492 272644
rect 473400 272640 473492 272642
rect 473400 272584 473450 272640
rect 473400 272582 473492 272584
rect 473445 272580 473492 272582
rect 473556 272580 473562 272644
rect 475837 272642 475884 272644
rect 475792 272640 475884 272642
rect 475792 272584 475842 272640
rect 475792 272582 475884 272584
rect 475837 272580 475884 272582
rect 475948 272580 475954 272644
rect 298461 272579 298527 272580
rect 300853 272579 300919 272580
rect 473445 272579 473511 272580
rect 475837 272579 475903 272580
rect 57462 272444 57468 272508
rect 57532 272506 57538 272508
rect 60917 272506 60983 272509
rect 119102 272506 119108 272508
rect 57532 272504 119108 272506
rect 57532 272448 60922 272504
rect 60978 272448 119108 272504
rect 57532 272446 119108 272448
rect 57532 272444 57538 272446
rect 60917 272443 60983 272446
rect 119102 272444 119108 272446
rect 119172 272444 119178 272508
rect 217174 272444 217180 272508
rect 217244 272506 217250 272508
rect 293350 272506 293356 272508
rect 217244 272446 293356 272506
rect 217244 272444 217250 272446
rect 293350 272444 293356 272446
rect 293420 272444 293426 272508
rect 82997 272372 83063 272373
rect 82997 272370 83044 272372
rect 82952 272368 83044 272370
rect 82952 272312 83002 272368
rect 82952 272310 83044 272312
rect 82997 272308 83044 272310
rect 83108 272308 83114 272372
rect 95693 272370 95759 272373
rect 101806 272370 101812 272372
rect 95693 272368 101812 272370
rect 95693 272312 95698 272368
rect 95754 272312 101812 272368
rect 95693 272310 101812 272312
rect 82997 272307 83063 272308
rect 95693 272307 95759 272310
rect 101806 272308 101812 272310
rect 101876 272308 101882 272372
rect 85389 272236 85455 272237
rect 113541 272236 113607 272237
rect 235993 272236 236059 272237
rect 85389 272234 85436 272236
rect 85344 272232 85436 272234
rect 85344 272176 85394 272232
rect 85344 272174 85436 272176
rect 85389 272172 85436 272174
rect 85500 272172 85506 272236
rect 113541 272234 113588 272236
rect 113496 272232 113588 272234
rect 113496 272176 113546 272232
rect 113496 272174 113588 272176
rect 113541 272172 113588 272174
rect 113652 272172 113658 272236
rect 235942 272172 235948 272236
rect 236012 272234 236059 272236
rect 401685 272236 401751 272237
rect 455781 272236 455847 272237
rect 401685 272234 401732 272236
rect 236012 272232 236104 272234
rect 236054 272176 236104 272232
rect 236012 272174 236104 272176
rect 401640 272232 401732 272234
rect 401640 272176 401690 272232
rect 401640 272174 401732 272176
rect 236012 272172 236059 272174
rect 85389 272171 85455 272172
rect 113541 272171 113607 272172
rect 235993 272171 236059 272172
rect 401685 272172 401732 272174
rect 401796 272172 401802 272236
rect 455781 272234 455828 272236
rect 455736 272232 455828 272234
rect 455736 272176 455786 272232
rect 455736 272174 455828 272176
rect 455781 272172 455828 272174
rect 455892 272172 455898 272236
rect 580349 272234 580415 272237
rect 583520 272234 584960 272324
rect 580349 272232 584960 272234
rect 580349 272176 580354 272232
rect 580410 272176 584960 272232
rect 580349 272174 584960 272176
rect 401685 272171 401751 272172
rect 455781 272171 455847 272172
rect 580349 272171 580415 272174
rect 583520 272084 584960 272174
rect 47485 271826 47551 271829
rect 49049 271826 49115 271829
rect 47485 271824 49115 271826
rect 47485 271768 47490 271824
rect 47546 271768 49054 271824
rect 49110 271768 49115 271824
rect 47485 271766 49115 271768
rect 47485 271763 47551 271766
rect 49049 271763 49115 271766
rect 75913 271826 75979 271829
rect 76046 271826 76052 271828
rect 75913 271824 76052 271826
rect 75913 271768 75918 271824
rect 75974 271768 76052 271824
rect 75913 271766 76052 271768
rect 75913 271763 75979 271766
rect 76046 271764 76052 271766
rect 76116 271764 76122 271828
rect 83958 271764 83964 271828
rect 84028 271826 84034 271828
rect 84193 271826 84259 271829
rect 84028 271824 84259 271826
rect 84028 271768 84198 271824
rect 84254 271768 84259 271824
rect 84028 271766 84259 271768
rect 84028 271764 84034 271766
rect 84193 271763 84259 271766
rect 88333 271826 88399 271829
rect 88742 271826 88748 271828
rect 88333 271824 88748 271826
rect 88333 271768 88338 271824
rect 88394 271768 88748 271824
rect 88333 271766 88748 271768
rect 88333 271763 88399 271766
rect 88742 271764 88748 271766
rect 88812 271764 88818 271828
rect 94221 271826 94287 271829
rect 94446 271826 94452 271828
rect 94221 271824 94452 271826
rect 94221 271768 94226 271824
rect 94282 271768 94452 271824
rect 94221 271766 94452 271768
rect 94221 271763 94287 271766
rect 94446 271764 94452 271766
rect 94516 271764 94522 271828
rect 102133 271826 102199 271829
rect 102726 271826 102732 271828
rect 102133 271824 102732 271826
rect 102133 271768 102138 271824
rect 102194 271768 102732 271824
rect 102133 271766 102732 271768
rect 102133 271763 102199 271766
rect 102726 271764 102732 271766
rect 102796 271764 102802 271828
rect 107653 271826 107719 271829
rect 108246 271826 108252 271828
rect 107653 271824 108252 271826
rect 107653 271768 107658 271824
rect 107714 271768 108252 271824
rect 107653 271766 108252 271768
rect 107653 271763 107719 271766
rect 108246 271764 108252 271766
rect 108316 271764 108322 271828
rect 125593 271826 125659 271829
rect 143533 271828 143599 271829
rect 125910 271826 125916 271828
rect 125593 271824 125916 271826
rect 125593 271768 125598 271824
rect 125654 271768 125916 271824
rect 125593 271766 125916 271768
rect 125593 271763 125659 271766
rect 125910 271764 125916 271766
rect 125980 271764 125986 271828
rect 143533 271826 143580 271828
rect 143488 271824 143580 271826
rect 143488 271768 143538 271824
rect 143488 271766 143580 271768
rect 143533 271764 143580 271766
rect 143644 271764 143650 271828
rect 154062 271764 154068 271828
rect 154132 271826 154138 271828
rect 154481 271826 154547 271829
rect 154132 271824 154547 271826
rect 154132 271768 154486 271824
rect 154542 271768 154547 271824
rect 154132 271766 154547 271768
rect 154132 271764 154138 271766
rect 143533 271763 143599 271764
rect 154481 271763 154547 271766
rect 155902 271764 155908 271828
rect 155972 271826 155978 271828
rect 157241 271826 157307 271829
rect 155972 271824 157307 271826
rect 155972 271768 157246 271824
rect 157302 271768 157307 271824
rect 155972 271766 157307 271768
rect 155972 271764 155978 271766
rect 157241 271763 157307 271766
rect 158478 271764 158484 271828
rect 158548 271826 158554 271828
rect 158621 271826 158687 271829
rect 158548 271824 158687 271826
rect 158548 271768 158626 271824
rect 158682 271768 158687 271824
rect 158548 271766 158687 271768
rect 158548 271764 158554 271766
rect 158621 271763 158687 271766
rect 213862 271764 213868 271828
rect 213932 271826 213938 271828
rect 214097 271826 214163 271829
rect 213932 271824 214163 271826
rect 213932 271768 214102 271824
rect 214158 271768 214163 271824
rect 213932 271766 214163 271768
rect 213932 271764 213938 271766
rect 214097 271763 214163 271766
rect 255313 271826 255379 271829
rect 263593 271828 263659 271829
rect 256182 271826 256188 271828
rect 255313 271824 256188 271826
rect 255313 271768 255318 271824
rect 255374 271768 256188 271824
rect 255313 271766 256188 271768
rect 255313 271763 255379 271766
rect 256182 271764 256188 271766
rect 256252 271764 256258 271828
rect 263542 271764 263548 271828
rect 263612 271826 263659 271828
rect 264973 271826 265039 271829
rect 265934 271826 265940 271828
rect 263612 271824 263704 271826
rect 263654 271768 263704 271824
rect 263612 271766 263704 271768
rect 264973 271824 265940 271826
rect 264973 271768 264978 271824
rect 265034 271768 265940 271824
rect 264973 271766 265940 271768
rect 263612 271764 263659 271766
rect 263593 271763 263659 271764
rect 264973 271763 265039 271766
rect 265934 271764 265940 271766
rect 266004 271764 266010 271828
rect 268009 271826 268075 271829
rect 268326 271826 268332 271828
rect 268009 271824 268332 271826
rect 268009 271768 268014 271824
rect 268070 271768 268332 271824
rect 268009 271766 268332 271768
rect 268009 271763 268075 271766
rect 268326 271764 268332 271766
rect 268396 271764 268402 271828
rect 270493 271826 270559 271829
rect 270902 271826 270908 271828
rect 270493 271824 270908 271826
rect 270493 271768 270498 271824
rect 270554 271768 270908 271824
rect 270493 271766 270908 271768
rect 270493 271763 270559 271766
rect 270902 271764 270908 271766
rect 270972 271764 270978 271828
rect 273253 271826 273319 271829
rect 273478 271826 273484 271828
rect 273253 271824 273484 271826
rect 273253 271768 273258 271824
rect 273314 271768 273484 271824
rect 273253 271766 273484 271768
rect 273253 271763 273319 271766
rect 273478 271764 273484 271766
rect 273548 271764 273554 271828
rect 275318 271764 275324 271828
rect 275388 271826 275394 271828
rect 275921 271826 275987 271829
rect 275388 271824 275987 271826
rect 275388 271768 275926 271824
rect 275982 271768 275987 271824
rect 275388 271766 275987 271768
rect 275388 271764 275394 271766
rect 275921 271763 275987 271766
rect 276105 271826 276171 271829
rect 276238 271826 276244 271828
rect 276105 271824 276244 271826
rect 276105 271768 276110 271824
rect 276166 271768 276244 271824
rect 276105 271766 276244 271768
rect 276105 271763 276171 271766
rect 276238 271764 276244 271766
rect 276308 271764 276314 271828
rect 276974 271764 276980 271828
rect 277044 271826 277050 271828
rect 277209 271826 277275 271829
rect 277044 271824 277275 271826
rect 277044 271768 277214 271824
rect 277270 271768 277275 271824
rect 277044 271766 277275 271768
rect 277044 271764 277050 271766
rect 277209 271763 277275 271766
rect 278078 271764 278084 271828
rect 278148 271826 278154 271828
rect 278681 271826 278747 271829
rect 278148 271824 278747 271826
rect 278148 271768 278686 271824
rect 278742 271768 278747 271824
rect 278148 271766 278747 271768
rect 278148 271764 278154 271766
rect 278681 271763 278747 271766
rect 302233 271826 302299 271829
rect 303470 271826 303476 271828
rect 302233 271824 303476 271826
rect 302233 271768 302238 271824
rect 302294 271768 303476 271824
rect 302233 271766 303476 271768
rect 302233 271763 302299 271766
rect 303470 271764 303476 271766
rect 303540 271764 303546 271828
rect 307753 271826 307819 271829
rect 308622 271826 308628 271828
rect 307753 271824 308628 271826
rect 307753 271768 307758 271824
rect 307814 271768 308628 271824
rect 307753 271766 308628 271768
rect 307753 271763 307819 271766
rect 308622 271764 308628 271766
rect 308692 271764 308698 271828
rect 403525 271826 403591 271829
rect 404118 271826 404124 271828
rect 403525 271824 404124 271826
rect 403525 271768 403530 271824
rect 403586 271768 404124 271824
rect 403525 271766 404124 271768
rect 403525 271763 403591 271766
rect 404118 271764 404124 271766
rect 404188 271764 404194 271828
rect 425053 271826 425119 271829
rect 425278 271826 425284 271828
rect 425053 271824 425284 271826
rect 425053 271768 425058 271824
rect 425114 271768 425284 271824
rect 425053 271766 425284 271768
rect 425053 271763 425119 271766
rect 425278 271764 425284 271766
rect 425348 271764 425354 271828
rect 427997 271826 428063 271829
rect 428590 271826 428596 271828
rect 427997 271824 428596 271826
rect 427997 271768 428002 271824
rect 428058 271768 428596 271824
rect 427997 271766 428596 271768
rect 427997 271763 428063 271766
rect 428590 271764 428596 271766
rect 428660 271764 428666 271828
rect 439262 271764 439268 271828
rect 439332 271826 439338 271828
rect 440141 271826 440207 271829
rect 439332 271824 440207 271826
rect 439332 271768 440146 271824
rect 440202 271768 440207 271824
rect 439332 271766 440207 271768
rect 439332 271764 439338 271766
rect 440141 271763 440207 271766
rect 447133 271826 447199 271829
rect 448278 271826 448284 271828
rect 447133 271824 448284 271826
rect 447133 271768 447138 271824
rect 447194 271768 448284 271824
rect 447133 271766 448284 271768
rect 447133 271763 447199 271766
rect 448278 271764 448284 271766
rect 448348 271764 448354 271828
rect 449893 271826 449959 271829
rect 451038 271826 451044 271828
rect 449893 271824 451044 271826
rect 449893 271768 449898 271824
rect 449954 271768 451044 271824
rect 449893 271766 451044 271768
rect 449893 271763 449959 271766
rect 451038 271764 451044 271766
rect 451108 271764 451114 271828
rect 452653 271826 452719 271829
rect 453430 271826 453436 271828
rect 452653 271824 453436 271826
rect 452653 271768 452658 271824
rect 452714 271768 453436 271824
rect 452653 271766 453436 271768
rect 452653 271763 452719 271766
rect 453430 271764 453436 271766
rect 453500 271764 453506 271828
rect 458173 271826 458239 271829
rect 460933 271828 460999 271829
rect 458398 271826 458404 271828
rect 458173 271824 458404 271826
rect 458173 271768 458178 271824
rect 458234 271768 458404 271824
rect 458173 271766 458404 271768
rect 458173 271763 458239 271766
rect 458398 271764 458404 271766
rect 458468 271764 458474 271828
rect 460933 271824 460980 271828
rect 461044 271826 461050 271828
rect 460933 271768 460938 271824
rect 460933 271764 460980 271768
rect 461044 271766 461090 271826
rect 461044 271764 461050 271766
rect 460933 271763 460999 271764
rect 47853 271690 47919 271693
rect 80462 271690 80468 271692
rect 47853 271688 80468 271690
rect 47853 271632 47858 271688
rect 47914 271632 80468 271688
rect 47853 271630 80468 271632
rect 47853 271627 47919 271630
rect 80462 271628 80468 271630
rect 80532 271628 80538 271692
rect 103513 271690 103579 271693
rect 103830 271690 103836 271692
rect 103513 271688 103836 271690
rect 103513 271632 103518 271688
rect 103574 271632 103836 271688
rect 103513 271630 103836 271632
rect 103513 271627 103579 271630
rect 103830 271628 103836 271630
rect 103900 271628 103906 271692
rect 110413 271690 110479 271693
rect 111006 271690 111012 271692
rect 110413 271688 111012 271690
rect 110413 271632 110418 271688
rect 110474 271632 111012 271688
rect 110413 271630 111012 271632
rect 110413 271627 110479 271630
rect 111006 271628 111012 271630
rect 111076 271628 111082 271692
rect 120073 271690 120139 271693
rect 120758 271690 120764 271692
rect 120073 271688 120764 271690
rect 120073 271632 120078 271688
rect 120134 271632 120764 271688
rect 120073 271630 120764 271632
rect 120073 271627 120139 271630
rect 120758 271628 120764 271630
rect 120828 271628 120834 271692
rect 123109 271690 123175 271693
rect 123518 271690 123524 271692
rect 123109 271688 123524 271690
rect 123109 271632 123114 271688
rect 123170 271632 123524 271688
rect 123109 271630 123524 271632
rect 123109 271627 123175 271630
rect 123518 271628 123524 271630
rect 123588 271628 123594 271692
rect 160870 271628 160876 271692
rect 160940 271690 160946 271692
rect 161381 271690 161447 271693
rect 160940 271688 161447 271690
rect 160940 271632 161386 271688
rect 161442 271632 161447 271688
rect 160940 271630 161447 271632
rect 160940 271628 160946 271630
rect 161381 271627 161447 271630
rect 163446 271628 163452 271692
rect 163516 271690 163522 271692
rect 164141 271690 164207 271693
rect 163516 271688 164207 271690
rect 163516 271632 164146 271688
rect 164202 271632 164207 271688
rect 163516 271630 164207 271632
rect 163516 271628 163522 271630
rect 164141 271627 164207 271630
rect 166022 271628 166028 271692
rect 166092 271690 166098 271692
rect 198958 271690 198964 271692
rect 166092 271630 198964 271690
rect 166092 271628 166098 271630
rect 198958 271628 198964 271630
rect 199028 271628 199034 271692
rect 216213 271690 216279 271693
rect 325550 271690 325556 271692
rect 216213 271688 325556 271690
rect 216213 271632 216218 271688
rect 216274 271632 325556 271688
rect 216213 271630 325556 271632
rect 216213 271627 216279 271630
rect 325550 271628 325556 271630
rect 325620 271628 325626 271692
rect 343214 271628 343220 271692
rect 343284 271690 343290 271692
rect 343541 271690 343607 271693
rect 343284 271688 343607 271690
rect 343284 271632 343546 271688
rect 343602 271632 343607 271688
rect 343284 271630 343607 271632
rect 343284 271628 343290 271630
rect 343541 271627 343607 271630
rect 379053 271690 379119 271693
rect 465942 271690 465948 271692
rect 379053 271688 465948 271690
rect 379053 271632 379058 271688
rect 379114 271632 465948 271688
rect 379053 271630 465948 271632
rect 379053 271627 379119 271630
rect 465942 271628 465948 271630
rect 466012 271628 466018 271692
rect 52453 271554 52519 271557
rect 52729 271554 52795 271557
rect 67541 271554 67607 271557
rect 52453 271552 67607 271554
rect 52453 271496 52458 271552
rect 52514 271496 52734 271552
rect 52790 271496 67546 271552
rect 67602 271496 67607 271552
rect 52453 271494 67607 271496
rect 52453 271491 52519 271494
rect 52729 271491 52795 271494
rect 67541 271491 67607 271494
rect 100753 271554 100819 271557
rect 115933 271556 115999 271557
rect 101070 271554 101076 271556
rect 100753 271552 101076 271554
rect 100753 271496 100758 271552
rect 100814 271496 101076 271552
rect 100753 271494 101076 271496
rect 100753 271491 100819 271494
rect 101070 271492 101076 271494
rect 101140 271492 101146 271556
rect 115933 271554 115980 271556
rect 115888 271552 115980 271554
rect 115888 271496 115938 271552
rect 115888 271494 115980 271496
rect 115933 271492 115980 271494
rect 116044 271492 116050 271556
rect 117313 271554 117379 271557
rect 118366 271554 118372 271556
rect 117313 271552 118372 271554
rect 117313 271496 117318 271552
rect 117374 271496 118372 271552
rect 117313 271494 118372 271496
rect 115933 271491 115999 271492
rect 117313 271491 117379 271494
rect 118366 271492 118372 271494
rect 118436 271492 118442 271556
rect 150934 271492 150940 271556
rect 151004 271554 151010 271556
rect 198774 271554 198780 271556
rect 151004 271494 198780 271554
rect 151004 271492 151010 271494
rect 198774 271492 198780 271494
rect 198844 271492 198850 271556
rect 206461 271554 206527 271557
rect 343449 271556 343515 271557
rect 315062 271554 315068 271556
rect 206461 271552 315068 271554
rect 206461 271496 206466 271552
rect 206522 271496 315068 271552
rect 206461 271494 315068 271496
rect 206461 271491 206527 271494
rect 315062 271492 315068 271494
rect 315132 271492 315138 271556
rect 343398 271492 343404 271556
rect 343468 271554 343515 271556
rect 343468 271552 343560 271554
rect 343510 271496 343560 271552
rect 343468 271494 343560 271496
rect 343468 271492 343515 271494
rect 379462 271492 379468 271556
rect 379532 271554 379538 271556
rect 413686 271554 413692 271556
rect 379532 271494 413692 271554
rect 379532 271492 379538 271494
rect 413686 271492 413692 271494
rect 413756 271492 413762 271556
rect 442993 271554 443059 271557
rect 443494 271554 443500 271556
rect 442993 271552 443500 271554
rect 442993 271496 442998 271552
rect 443054 271496 443500 271552
rect 442993 271494 443500 271496
rect 343449 271491 343515 271492
rect 442993 271491 443059 271494
rect 443494 271492 443500 271494
rect 443564 271492 443570 271556
rect 503478 271492 503484 271556
rect 503548 271554 503554 271556
rect 503621 271554 503687 271557
rect 503548 271552 503687 271554
rect 503548 271496 503626 271552
rect 503682 271496 503687 271552
rect 503548 271494 503687 271496
rect 503548 271492 503554 271494
rect 503621 271491 503687 271494
rect 77293 271418 77359 271421
rect 78254 271418 78260 271420
rect 77293 271416 78260 271418
rect 77293 271360 77298 271416
rect 77354 271360 78260 271416
rect 77293 271358 78260 271360
rect 77293 271355 77359 271358
rect 78254 271356 78260 271358
rect 78324 271356 78330 271420
rect 91185 271418 91251 271421
rect 91502 271418 91508 271420
rect 91185 271416 91508 271418
rect 91185 271360 91190 271416
rect 91246 271360 91508 271416
rect 91185 271358 91508 271360
rect 91185 271355 91251 271358
rect 91502 271356 91508 271358
rect 91572 271356 91578 271420
rect 104893 271418 104959 271421
rect 105854 271418 105860 271420
rect 104893 271416 105860 271418
rect 104893 271360 104898 271416
rect 104954 271360 105860 271416
rect 104893 271358 105860 271360
rect 104893 271355 104959 271358
rect 105854 271356 105860 271358
rect 105924 271356 105930 271420
rect 183134 271356 183140 271420
rect 183204 271418 183210 271420
rect 183461 271418 183527 271421
rect 183204 271416 183527 271418
rect 183204 271360 183466 271416
rect 183522 271360 183527 271416
rect 183204 271358 183527 271360
rect 183204 271356 183210 271358
rect 183461 271355 183527 271358
rect 213545 271418 213611 271421
rect 313406 271418 313412 271420
rect 213545 271416 313412 271418
rect 213545 271360 213550 271416
rect 213606 271360 313412 271416
rect 213545 271358 313412 271360
rect 213545 271355 213611 271358
rect 313406 271356 313412 271358
rect 313476 271356 313482 271420
rect 377254 271356 377260 271420
rect 377324 271418 377330 271420
rect 408166 271418 408172 271420
rect 377324 271358 408172 271418
rect 377324 271356 377330 271358
rect 408166 271356 408172 271358
rect 408236 271356 408242 271420
rect 418337 271418 418403 271421
rect 418470 271418 418476 271420
rect 418337 271416 418476 271418
rect 418337 271360 418342 271416
rect 418398 271360 418476 271416
rect 418337 271358 418476 271360
rect 418337 271355 418403 271358
rect 418470 271356 418476 271358
rect 418540 271356 418546 271420
rect 434713 271418 434779 271421
rect 435950 271418 435956 271420
rect 434713 271416 435956 271418
rect 434713 271360 434718 271416
rect 434774 271360 435956 271416
rect 434713 271358 435956 271360
rect 434713 271355 434779 271358
rect 435950 271356 435956 271358
rect 436020 271356 436026 271420
rect 445753 271418 445819 271421
rect 445886 271418 445892 271420
rect 445753 271416 445892 271418
rect 445753 271360 445758 271416
rect 445814 271360 445892 271416
rect 445753 271358 445892 271360
rect 445753 271355 445819 271358
rect 445886 271356 445892 271358
rect 445956 271356 445962 271420
rect 503110 271356 503116 271420
rect 503180 271418 503186 271420
rect 503529 271418 503595 271421
rect 503180 271416 503595 271418
rect 503180 271360 503534 271416
rect 503590 271360 503595 271416
rect 503180 271358 503595 271360
rect 503180 271356 503186 271358
rect 503529 271355 503595 271358
rect 49049 271282 49115 271285
rect 81934 271282 81940 271284
rect 49049 271280 81940 271282
rect 49049 271224 49054 271280
rect 49110 271224 81940 271280
rect 49049 271222 81940 271224
rect 49049 271219 49115 271222
rect 81934 271220 81940 271222
rect 82004 271220 82010 271284
rect 106273 271282 106339 271285
rect 107510 271282 107516 271284
rect 106273 271280 107516 271282
rect 106273 271224 106278 271280
rect 106334 271224 107516 271280
rect 106273 271222 107516 271224
rect 106273 271219 106339 271222
rect 107510 271220 107516 271222
rect 107580 271220 107586 271284
rect 258257 271282 258323 271285
rect 258390 271282 258396 271284
rect 258257 271280 258396 271282
rect 258257 271224 258262 271280
rect 258318 271224 258396 271280
rect 258257 271222 258396 271224
rect 258257 271219 258323 271222
rect 258390 271220 258396 271222
rect 258460 271220 258466 271284
rect 260833 271282 260899 271285
rect 260966 271282 260972 271284
rect 260833 271280 260972 271282
rect 260833 271224 260838 271280
rect 260894 271224 260972 271280
rect 260833 271222 260972 271224
rect 260833 271219 260899 271222
rect 260966 271220 260972 271222
rect 261036 271220 261042 271284
rect 278998 271220 279004 271284
rect 279068 271282 279074 271284
rect 280061 271282 280127 271285
rect 279068 271280 280127 271282
rect 279068 271224 280066 271280
rect 280122 271224 280127 271280
rect 279068 271222 280127 271224
rect 279068 271220 279074 271222
rect 280061 271219 280127 271222
rect 374361 271282 374427 271285
rect 397126 271282 397132 271284
rect 374361 271280 397132 271282
rect 374361 271224 374366 271280
rect 374422 271224 397132 271280
rect 374361 271222 397132 271224
rect 374361 271219 374427 271222
rect 397126 271220 397132 271222
rect 397196 271220 397202 271284
rect 416998 271282 417004 271284
rect 402930 271222 417004 271282
rect 47710 271084 47716 271148
rect 47780 271146 47786 271148
rect 53005 271146 53071 271149
rect 109534 271146 109540 271148
rect 47780 271144 109540 271146
rect 47780 271088 53010 271144
rect 53066 271088 109540 271144
rect 47780 271086 109540 271088
rect 47780 271084 47786 271086
rect 53005 271083 53071 271086
rect 109534 271084 109540 271086
rect 109604 271084 109610 271148
rect 128353 271146 128419 271149
rect 183461 271148 183527 271149
rect 128670 271146 128676 271148
rect 128353 271144 128676 271146
rect 128353 271088 128358 271144
rect 128414 271088 128676 271144
rect 128353 271086 128676 271088
rect 128353 271083 128419 271086
rect 128670 271084 128676 271086
rect 128740 271084 128746 271148
rect 183461 271146 183508 271148
rect 183416 271144 183508 271146
rect 183416 271088 183466 271144
rect 183416 271086 183508 271088
rect 183461 271084 183508 271086
rect 183572 271084 183578 271148
rect 239121 271146 239187 271149
rect 239254 271146 239260 271148
rect 239121 271144 239260 271146
rect 239121 271088 239126 271144
rect 239182 271088 239260 271144
rect 239121 271086 239260 271088
rect 183461 271083 183527 271084
rect 239121 271083 239187 271086
rect 239254 271084 239260 271086
rect 239324 271084 239330 271148
rect 247033 271146 247099 271149
rect 248270 271146 248276 271148
rect 247033 271144 248276 271146
rect 247033 271088 247038 271144
rect 247094 271088 248276 271144
rect 247033 271086 248276 271088
rect 247033 271083 247099 271086
rect 248270 271084 248276 271086
rect 248340 271084 248346 271148
rect 252553 271146 252619 271149
rect 253606 271146 253612 271148
rect 252553 271144 253612 271146
rect 252553 271088 252558 271144
rect 252614 271088 253612 271144
rect 252553 271086 253612 271088
rect 252553 271083 252619 271086
rect 253606 271084 253612 271086
rect 253676 271084 253682 271148
rect 260833 271146 260899 271149
rect 266353 271148 266419 271149
rect 262070 271146 262076 271148
rect 260833 271144 262076 271146
rect 260833 271088 260838 271144
rect 260894 271088 262076 271144
rect 260833 271086 262076 271088
rect 260833 271083 260899 271086
rect 262070 271084 262076 271086
rect 262140 271084 262146 271148
rect 266302 271084 266308 271148
rect 266372 271146 266419 271148
rect 268101 271146 268167 271149
rect 268694 271146 268700 271148
rect 266372 271144 266464 271146
rect 266414 271088 266464 271144
rect 266372 271086 266464 271088
rect 268101 271144 268700 271146
rect 268101 271088 268106 271144
rect 268162 271088 268700 271144
rect 268101 271086 268700 271088
rect 266372 271084 266419 271086
rect 266353 271083 266419 271084
rect 268101 271083 268167 271086
rect 268694 271084 268700 271086
rect 268764 271084 268770 271148
rect 270493 271146 270559 271149
rect 271270 271146 271276 271148
rect 270493 271144 271276 271146
rect 270493 271088 270498 271144
rect 270554 271088 271276 271144
rect 270493 271086 271276 271088
rect 270493 271083 270559 271086
rect 271270 271084 271276 271086
rect 271340 271084 271346 271148
rect 396717 271146 396783 271149
rect 402930 271146 402990 271222
rect 416998 271220 417004 271222
rect 417068 271220 417074 271284
rect 433333 271282 433399 271285
rect 433558 271282 433564 271284
rect 433333 271280 433564 271282
rect 433333 271224 433338 271280
rect 433394 271224 433564 271280
rect 433333 271222 433564 271224
rect 433333 271219 433399 271222
rect 433558 271220 433564 271222
rect 433628 271220 433634 271284
rect 437473 271282 437539 271285
rect 438526 271282 438532 271284
rect 437473 271280 438532 271282
rect 437473 271224 437478 271280
rect 437534 271224 438532 271280
rect 437473 271222 438532 271224
rect 437473 271219 437539 271222
rect 438526 271220 438532 271222
rect 438596 271220 438602 271284
rect 396717 271144 402990 271146
rect 396717 271088 396722 271144
rect 396778 271088 402990 271144
rect 396717 271086 402990 271088
rect 420913 271146 420979 271149
rect 421046 271146 421052 271148
rect 420913 271144 421052 271146
rect 420913 271088 420918 271144
rect 420974 271088 421052 271144
rect 420913 271086 421052 271088
rect 396717 271083 396783 271086
rect 420913 271083 420979 271086
rect 421046 271084 421052 271086
rect 421116 271084 421122 271148
rect 78673 271010 78739 271013
rect 79542 271010 79548 271012
rect 78673 271008 79548 271010
rect 78673 270952 78678 271008
rect 78734 270952 79548 271008
rect 78673 270950 79548 270952
rect 78673 270947 78739 270950
rect 79542 270948 79548 270950
rect 79612 270948 79618 271012
rect 104893 271010 104959 271013
rect 105302 271010 105308 271012
rect 104893 271008 105308 271010
rect 104893 270952 104898 271008
rect 104954 270952 105308 271008
rect 104893 270950 105308 270952
rect 104893 270947 104959 270950
rect 105302 270948 105308 270950
rect 105372 270948 105378 271012
rect 207749 271010 207815 271013
rect 320950 271010 320956 271012
rect 207749 271008 320956 271010
rect 207749 270952 207754 271008
rect 207810 270952 320956 271008
rect 207749 270950 320956 270952
rect 207749 270947 207815 270950
rect 320950 270948 320956 270950
rect 321020 270948 321026 271012
rect 409873 271010 409939 271013
rect 410742 271010 410748 271012
rect 409873 271008 410748 271010
rect 409873 270952 409878 271008
rect 409934 270952 410748 271008
rect 409873 270950 410748 270952
rect 409873 270947 409939 270950
rect 410742 270948 410748 270950
rect 410812 270948 410818 271012
rect 429193 271010 429259 271013
rect 429694 271010 429700 271012
rect 429193 271008 429700 271010
rect 429193 270952 429198 271008
rect 429254 270952 429700 271008
rect 429193 270950 429700 270952
rect 429193 270947 429259 270950
rect 429694 270948 429700 270950
rect 429764 270948 429770 271012
rect 437473 271010 437539 271013
rect 438342 271010 438348 271012
rect 437473 271008 438348 271010
rect 437473 270952 437478 271008
rect 437534 270952 438348 271008
rect 437473 270950 438348 270952
rect 437473 270947 437539 270950
rect 438342 270948 438348 270950
rect 438412 270948 438418 271012
rect 96613 270874 96679 270877
rect 97022 270874 97028 270876
rect 96613 270872 97028 270874
rect 96613 270816 96618 270872
rect 96674 270816 97028 270872
rect 96613 270814 97028 270816
rect 96613 270811 96679 270814
rect 97022 270812 97028 270814
rect 97092 270812 97098 270876
rect 115933 270874 115999 270877
rect 116894 270874 116900 270876
rect 115933 270872 116900 270874
rect 115933 270816 115938 270872
rect 115994 270816 116900 270872
rect 115933 270814 116900 270816
rect 115933 270811 115999 270814
rect 116894 270812 116900 270814
rect 116964 270812 116970 270876
rect 147673 270874 147739 270877
rect 148542 270874 148548 270876
rect 147673 270872 148548 270874
rect 147673 270816 147678 270872
rect 147734 270816 148548 270872
rect 147673 270814 148548 270816
rect 147673 270811 147739 270814
rect 148542 270812 148548 270814
rect 148612 270812 148618 270876
rect 252553 270874 252619 270877
rect 253422 270874 253428 270876
rect 252553 270872 253428 270874
rect 252553 270816 252558 270872
rect 252614 270816 253428 270872
rect 252553 270814 253428 270816
rect 252553 270811 252619 270814
rect 253422 270812 253428 270814
rect 253492 270812 253498 270876
rect 264973 270874 265039 270877
rect 265750 270874 265756 270876
rect 264973 270872 265756 270874
rect 264973 270816 264978 270872
rect 265034 270816 265756 270872
rect 264973 270814 265756 270816
rect 264973 270811 265039 270814
rect 265750 270812 265756 270814
rect 265820 270812 265826 270876
rect 364057 270874 364123 270877
rect 462630 270874 462636 270876
rect 364057 270872 462636 270874
rect 364057 270816 364062 270872
rect 364118 270816 462636 270872
rect 364057 270814 462636 270816
rect 364057 270811 364123 270814
rect 462630 270812 462636 270814
rect 462700 270812 462706 270876
rect 85573 270738 85639 270741
rect 86534 270738 86540 270740
rect 85573 270736 86540 270738
rect 85573 270680 85578 270736
rect 85634 270680 86540 270736
rect 85573 270678 86540 270680
rect 85573 270675 85639 270678
rect 86534 270676 86540 270678
rect 86604 270676 86610 270740
rect 89713 270738 89779 270741
rect 90030 270738 90036 270740
rect 89713 270736 90036 270738
rect 89713 270680 89718 270736
rect 89774 270680 90036 270736
rect 89713 270678 90036 270680
rect 89713 270675 89779 270678
rect 90030 270676 90036 270678
rect 90100 270676 90106 270740
rect 92473 270738 92539 270741
rect 93342 270738 93348 270740
rect 92473 270736 93348 270738
rect 92473 270680 92478 270736
rect 92534 270680 93348 270736
rect 92473 270678 93348 270680
rect 92473 270675 92539 270678
rect 93342 270676 93348 270678
rect 93412 270676 93418 270740
rect 244273 270738 244339 270741
rect 245326 270738 245332 270740
rect 244273 270736 245332 270738
rect 244273 270680 244278 270736
rect 244334 270680 245332 270736
rect 244273 270678 245332 270680
rect 244273 270675 244339 270678
rect 245326 270676 245332 270678
rect 245396 270676 245402 270740
rect 251265 270738 251331 270741
rect 252318 270738 252324 270740
rect 251265 270736 252324 270738
rect 251265 270680 251270 270736
rect 251326 270680 252324 270736
rect 251265 270678 252324 270680
rect 251265 270675 251331 270678
rect 252318 270676 252324 270678
rect 252388 270676 252394 270740
rect 259545 270738 259611 270741
rect 260598 270738 260604 270740
rect 259545 270736 260604 270738
rect 259545 270680 259550 270736
rect 259606 270680 260604 270736
rect 259545 270678 260604 270680
rect 259545 270675 259611 270678
rect 260598 270676 260604 270678
rect 260668 270676 260674 270740
rect 265617 270738 265683 270741
rect 411345 270740 411411 270741
rect 267590 270738 267596 270740
rect 265617 270736 267596 270738
rect 265617 270680 265622 270736
rect 265678 270680 267596 270736
rect 265617 270678 267596 270680
rect 265617 270675 265683 270678
rect 267590 270676 267596 270678
rect 267660 270676 267666 270740
rect 411294 270676 411300 270740
rect 411364 270738 411411 270740
rect 431953 270738 432019 270741
rect 432270 270738 432276 270740
rect 411364 270736 411456 270738
rect 411406 270680 411456 270736
rect 411364 270678 411456 270680
rect 431953 270736 432276 270738
rect 431953 270680 431958 270736
rect 432014 270680 432276 270736
rect 431953 270678 432276 270680
rect 411364 270676 411411 270678
rect 411345 270675 411411 270676
rect 431953 270675 432019 270678
rect 432270 270676 432276 270678
rect 432340 270676 432346 270740
rect 54569 270602 54635 270605
rect 58709 270602 58775 270605
rect 54569 270600 58775 270602
rect 54569 270544 54574 270600
rect 54630 270544 58714 270600
rect 58770 270544 58775 270600
rect 54569 270542 58775 270544
rect 54569 270539 54635 270542
rect 58709 270539 58775 270542
rect 86953 270602 87019 270605
rect 87638 270602 87644 270604
rect 86953 270600 87644 270602
rect 86953 270544 86958 270600
rect 87014 270544 87644 270600
rect 86953 270542 87644 270544
rect 86953 270539 87019 270542
rect 87638 270540 87644 270542
rect 87708 270540 87714 270604
rect 91093 270602 91159 270605
rect 91318 270602 91324 270604
rect 91093 270600 91324 270602
rect 91093 270544 91098 270600
rect 91154 270544 91324 270600
rect 91093 270542 91324 270544
rect 91093 270539 91159 270542
rect 91318 270540 91324 270542
rect 91388 270540 91394 270604
rect 103697 270602 103763 270605
rect 106365 270604 106431 270605
rect 104014 270602 104020 270604
rect 103697 270600 104020 270602
rect 103697 270544 103702 270600
rect 103758 270544 104020 270600
rect 103697 270542 104020 270544
rect 103697 270539 103763 270542
rect 104014 270540 104020 270542
rect 104084 270540 104090 270604
rect 106365 270602 106412 270604
rect 106320 270600 106412 270602
rect 106320 270544 106370 270600
rect 106320 270542 106412 270544
rect 106365 270540 106412 270542
rect 106476 270540 106482 270604
rect 107653 270602 107719 270605
rect 108614 270602 108620 270604
rect 107653 270600 108620 270602
rect 107653 270544 107658 270600
rect 107714 270544 108620 270600
rect 107653 270542 108620 270544
rect 106365 270539 106431 270540
rect 107653 270539 107719 270542
rect 108614 270540 108620 270542
rect 108684 270540 108690 270604
rect 110413 270602 110479 270605
rect 113173 270604 113239 270605
rect 114461 270604 114527 270605
rect 115841 270604 115907 270605
rect 111190 270602 111196 270604
rect 110413 270600 111196 270602
rect 110413 270544 110418 270600
rect 110474 270544 111196 270600
rect 110413 270542 111196 270544
rect 110413 270539 110479 270542
rect 111190 270540 111196 270542
rect 111260 270540 111266 270604
rect 113173 270600 113220 270604
rect 113284 270602 113290 270604
rect 114461 270602 114508 270604
rect 113173 270544 113178 270600
rect 113173 270540 113220 270544
rect 113284 270542 113330 270602
rect 114416 270600 114508 270602
rect 114416 270544 114466 270600
rect 114416 270542 114508 270544
rect 113284 270540 113290 270542
rect 114461 270540 114508 270542
rect 114572 270540 114578 270604
rect 115790 270540 115796 270604
rect 115860 270602 115907 270604
rect 235993 270602 236059 270605
rect 237046 270602 237052 270604
rect 115860 270600 115952 270602
rect 115902 270544 115952 270600
rect 115860 270542 115952 270544
rect 235993 270600 237052 270602
rect 235993 270544 235998 270600
rect 236054 270544 237052 270600
rect 235993 270542 237052 270544
rect 115860 270540 115907 270542
rect 113173 270539 113239 270540
rect 114461 270539 114527 270540
rect 115841 270539 115907 270540
rect 235993 270539 236059 270542
rect 237046 270540 237052 270542
rect 237116 270540 237122 270604
rect 237373 270602 237439 270605
rect 242893 270604 242959 270605
rect 238150 270602 238156 270604
rect 237373 270600 238156 270602
rect 237373 270544 237378 270600
rect 237434 270544 238156 270600
rect 237373 270542 238156 270544
rect 237373 270539 237439 270542
rect 238150 270540 238156 270542
rect 238220 270540 238226 270604
rect 242893 270602 242940 270604
rect 242848 270600 242940 270602
rect 242848 270544 242898 270600
rect 242848 270542 242940 270544
rect 242893 270540 242940 270542
rect 243004 270540 243010 270604
rect 244222 270540 244228 270604
rect 244292 270602 244298 270604
rect 244365 270602 244431 270605
rect 244292 270600 244431 270602
rect 244292 270544 244370 270600
rect 244426 270544 244431 270600
rect 244292 270542 244431 270544
rect 244292 270540 244298 270542
rect 242893 270539 242959 270540
rect 244365 270539 244431 270542
rect 245653 270602 245719 270605
rect 246430 270602 246436 270604
rect 245653 270600 246436 270602
rect 245653 270544 245658 270600
rect 245714 270544 246436 270600
rect 245653 270542 246436 270544
rect 245653 270539 245719 270542
rect 246430 270540 246436 270542
rect 246500 270540 246506 270604
rect 247033 270602 247099 270605
rect 247718 270602 247724 270604
rect 247033 270600 247724 270602
rect 247033 270544 247038 270600
rect 247094 270544 247724 270600
rect 247033 270542 247724 270544
rect 247033 270539 247099 270542
rect 247718 270540 247724 270542
rect 247788 270540 247794 270604
rect 248505 270602 248571 270605
rect 248638 270602 248644 270604
rect 248505 270600 248644 270602
rect 248505 270544 248510 270600
rect 248566 270544 248644 270600
rect 248505 270542 248644 270544
rect 248505 270539 248571 270542
rect 248638 270540 248644 270542
rect 248708 270540 248714 270604
rect 249793 270602 249859 270605
rect 251173 270604 251239 270605
rect 250110 270602 250116 270604
rect 249793 270600 250116 270602
rect 249793 270544 249798 270600
rect 249854 270544 250116 270600
rect 249793 270542 250116 270544
rect 249793 270539 249859 270542
rect 250110 270540 250116 270542
rect 250180 270540 250186 270604
rect 251173 270602 251220 270604
rect 251128 270600 251220 270602
rect 251128 270544 251178 270600
rect 251128 270542 251220 270544
rect 251173 270540 251220 270542
rect 251284 270540 251290 270604
rect 253933 270602 253999 270605
rect 254526 270602 254532 270604
rect 253933 270600 254532 270602
rect 253933 270544 253938 270600
rect 253994 270544 254532 270600
rect 253933 270542 254532 270544
rect 251173 270539 251239 270540
rect 253933 270539 253999 270542
rect 254526 270540 254532 270542
rect 254596 270540 254602 270604
rect 255313 270602 255379 270605
rect 255814 270602 255820 270604
rect 255313 270600 255820 270602
rect 255313 270544 255318 270600
rect 255374 270544 255820 270600
rect 255313 270542 255820 270544
rect 255313 270539 255379 270542
rect 255814 270540 255820 270542
rect 255884 270540 255890 270604
rect 256693 270602 256759 270605
rect 256918 270602 256924 270604
rect 256693 270600 256924 270602
rect 256693 270544 256698 270600
rect 256754 270544 256924 270600
rect 256693 270542 256924 270544
rect 256693 270539 256759 270542
rect 256918 270540 256924 270542
rect 256988 270540 256994 270604
rect 258073 270602 258139 270605
rect 259453 270604 259519 270605
rect 258390 270602 258396 270604
rect 258073 270600 258396 270602
rect 258073 270544 258078 270600
rect 258134 270544 258396 270600
rect 258073 270542 258396 270544
rect 258073 270539 258139 270542
rect 258390 270540 258396 270542
rect 258460 270540 258466 270604
rect 259453 270602 259500 270604
rect 259408 270600 259500 270602
rect 259408 270544 259458 270600
rect 259408 270542 259500 270544
rect 259453 270540 259500 270542
rect 259564 270540 259570 270604
rect 262213 270602 262279 270605
rect 262806 270602 262812 270604
rect 262213 270600 262812 270602
rect 262213 270544 262218 270600
rect 262274 270544 262812 270600
rect 262213 270542 262812 270544
rect 259453 270539 259519 270540
rect 262213 270539 262279 270542
rect 262806 270540 262812 270542
rect 262876 270540 262882 270604
rect 263593 270602 263659 270605
rect 263910 270602 263916 270604
rect 263593 270600 263916 270602
rect 263593 270544 263598 270600
rect 263654 270544 263916 270600
rect 263593 270542 263916 270544
rect 263593 270539 263659 270542
rect 263910 270540 263916 270542
rect 263980 270540 263986 270604
rect 269113 270602 269179 270605
rect 269798 270602 269804 270604
rect 269113 270600 269804 270602
rect 269113 270544 269118 270600
rect 269174 270544 269804 270600
rect 269113 270542 269804 270544
rect 269113 270539 269179 270542
rect 269798 270540 269804 270542
rect 269868 270540 269874 270604
rect 273253 270602 273319 270605
rect 396073 270604 396139 270605
rect 274398 270602 274404 270604
rect 273253 270600 274404 270602
rect 273253 270544 273258 270600
rect 273314 270544 274404 270600
rect 273253 270542 274404 270544
rect 273253 270539 273319 270542
rect 274398 270540 274404 270542
rect 274468 270540 274474 270604
rect 396022 270540 396028 270604
rect 396092 270602 396139 270604
rect 397453 270604 397519 270605
rect 397453 270602 397500 270604
rect 396092 270600 396184 270602
rect 396134 270544 396184 270600
rect 396092 270542 396184 270544
rect 397408 270600 397500 270602
rect 397408 270544 397458 270600
rect 397408 270542 397500 270544
rect 396092 270540 396139 270542
rect 396073 270539 396139 270540
rect 397453 270540 397500 270542
rect 397564 270540 397570 270604
rect 398833 270602 398899 270605
rect 399518 270602 399524 270604
rect 398833 270600 399524 270602
rect 398833 270544 398838 270600
rect 398894 270544 399524 270600
rect 398833 270542 399524 270544
rect 397453 270539 397519 270540
rect 398833 270539 398899 270542
rect 399518 270540 399524 270542
rect 399588 270540 399594 270604
rect 400213 270602 400279 270605
rect 402973 270604 403039 270605
rect 400438 270602 400444 270604
rect 400213 270600 400444 270602
rect 400213 270544 400218 270600
rect 400274 270544 400444 270600
rect 400213 270542 400444 270544
rect 400213 270539 400279 270542
rect 400438 270540 400444 270542
rect 400508 270540 400514 270604
rect 402973 270600 403020 270604
rect 403084 270602 403090 270604
rect 404353 270602 404419 270605
rect 405038 270602 405044 270604
rect 402973 270544 402978 270600
rect 402973 270540 403020 270544
rect 403084 270542 403130 270602
rect 404353 270600 405044 270602
rect 404353 270544 404358 270600
rect 404414 270544 405044 270600
rect 404353 270542 405044 270544
rect 403084 270540 403090 270542
rect 402973 270539 403039 270540
rect 404353 270539 404419 270542
rect 405038 270540 405044 270542
rect 405108 270540 405114 270604
rect 405733 270602 405799 270605
rect 406510 270602 406516 270604
rect 405733 270600 406516 270602
rect 405733 270544 405738 270600
rect 405794 270544 406516 270600
rect 405733 270542 406516 270544
rect 405733 270539 405799 270542
rect 406510 270540 406516 270542
rect 406580 270540 406586 270604
rect 407113 270602 407179 270605
rect 407614 270602 407620 270604
rect 407113 270600 407620 270602
rect 407113 270544 407118 270600
rect 407174 270544 407620 270600
rect 407113 270542 407620 270544
rect 407113 270539 407179 270542
rect 407614 270540 407620 270542
rect 407684 270540 407690 270604
rect 408493 270602 408559 270605
rect 408718 270602 408724 270604
rect 408493 270600 408724 270602
rect 408493 270544 408498 270600
rect 408554 270544 408724 270600
rect 408493 270542 408724 270544
rect 408493 270539 408559 270542
rect 408718 270540 408724 270542
rect 408788 270540 408794 270604
rect 409873 270602 409939 270605
rect 410006 270602 410012 270604
rect 409873 270600 410012 270602
rect 409873 270544 409878 270600
rect 409934 270544 410012 270600
rect 409873 270542 410012 270544
rect 409873 270539 409939 270542
rect 410006 270540 410012 270542
rect 410076 270540 410082 270604
rect 411253 270602 411319 270605
rect 412398 270602 412404 270604
rect 411253 270600 412404 270602
rect 411253 270544 411258 270600
rect 411314 270544 412404 270600
rect 411253 270542 412404 270544
rect 411253 270539 411319 270542
rect 412398 270540 412404 270542
rect 412468 270540 412474 270604
rect 413001 270602 413067 270605
rect 413318 270602 413324 270604
rect 413001 270600 413324 270602
rect 413001 270544 413006 270600
rect 413062 270544 413324 270600
rect 413001 270542 413324 270544
rect 413001 270539 413067 270542
rect 413318 270540 413324 270542
rect 413388 270540 413394 270604
rect 414013 270602 414079 270605
rect 414422 270602 414428 270604
rect 414013 270600 414428 270602
rect 414013 270544 414018 270600
rect 414074 270544 414428 270600
rect 414013 270542 414428 270544
rect 414013 270539 414079 270542
rect 414422 270540 414428 270542
rect 414492 270540 414498 270604
rect 415393 270602 415459 270605
rect 415526 270602 415532 270604
rect 415393 270600 415532 270602
rect 415393 270544 415398 270600
rect 415454 270544 415532 270600
rect 415393 270542 415532 270544
rect 415393 270539 415459 270542
rect 415526 270540 415532 270542
rect 415596 270540 415602 270604
rect 418153 270602 418219 270605
rect 418286 270602 418292 270604
rect 418153 270600 418292 270602
rect 418153 270544 418158 270600
rect 418214 270544 418292 270600
rect 418153 270542 418292 270544
rect 418153 270539 418219 270542
rect 418286 270540 418292 270542
rect 418356 270540 418362 270604
rect 418521 270602 418587 270605
rect 419206 270602 419212 270604
rect 418521 270600 419212 270602
rect 418521 270544 418526 270600
rect 418582 270544 419212 270600
rect 418521 270542 419212 270544
rect 418521 270539 418587 270542
rect 419206 270540 419212 270542
rect 419276 270540 419282 270604
rect 419533 270602 419599 270605
rect 420678 270602 420684 270604
rect 419533 270600 420684 270602
rect 419533 270544 419538 270600
rect 419594 270544 420684 270600
rect 419533 270542 420684 270544
rect 419533 270539 419599 270542
rect 420678 270540 420684 270542
rect 420748 270540 420754 270604
rect 420913 270602 420979 270605
rect 421782 270602 421788 270604
rect 420913 270600 421788 270602
rect 420913 270544 420918 270600
rect 420974 270544 421788 270600
rect 420913 270542 421788 270544
rect 420913 270539 420979 270542
rect 421782 270540 421788 270542
rect 421852 270540 421858 270604
rect 436093 270602 436159 270605
rect 436870 270602 436876 270604
rect 436093 270600 436876 270602
rect 436093 270544 436098 270600
rect 436154 270544 436876 270600
rect 436093 270542 436876 270544
rect 436093 270539 436159 270542
rect 436870 270540 436876 270542
rect 436940 270540 436946 270604
rect 202505 270466 202571 270469
rect 323342 270466 323348 270468
rect 202505 270464 323348 270466
rect 202505 270408 202510 270464
rect 202566 270408 323348 270464
rect 202505 270406 323348 270408
rect 202505 270403 202571 270406
rect 323342 270404 323348 270406
rect 323412 270404 323418 270468
rect 369577 270466 369643 270469
rect 372153 270466 372219 270469
rect 369577 270464 372219 270466
rect 369577 270408 369582 270464
rect 369638 270408 372158 270464
rect 372214 270408 372219 270464
rect 369577 270406 372219 270408
rect 369577 270403 369643 270406
rect 372153 270403 372219 270406
rect 375005 270466 375071 270469
rect 375925 270466 375991 270469
rect 435766 270466 435772 270468
rect 375005 270464 435772 270466
rect 375005 270408 375010 270464
rect 375066 270408 375930 270464
rect 375986 270408 435772 270464
rect 375005 270406 435772 270408
rect 375005 270403 375071 270406
rect 375925 270403 375991 270406
rect 435766 270404 435772 270406
rect 435836 270404 435842 270468
rect 208117 270330 208183 270333
rect 241646 270330 241652 270332
rect 208117 270328 241652 270330
rect 208117 270272 208122 270328
rect 208178 270272 241652 270328
rect 208117 270270 241652 270272
rect 208117 270267 208183 270270
rect 241646 270268 241652 270270
rect 241716 270268 241722 270332
rect 212901 270194 212967 270197
rect 214465 270194 214531 270197
rect 240542 270194 240548 270196
rect 212901 270192 240548 270194
rect 212901 270136 212906 270192
rect 212962 270136 214470 270192
rect 214526 270136 240548 270192
rect 212901 270134 240548 270136
rect 212901 270131 212967 270134
rect 214465 270131 214531 270134
rect 240542 270132 240548 270134
rect 240612 270132 240618 270196
rect 217317 270060 217383 270061
rect 217317 270058 217364 270060
rect 217272 270056 217364 270058
rect 217272 270000 217322 270056
rect 217272 269998 217364 270000
rect 217317 269996 217364 269998
rect 217428 269996 217434 270060
rect 217317 269995 217383 269996
rect 371601 269922 371667 269925
rect 376385 269922 376451 269925
rect 434662 269922 434668 269924
rect 371601 269920 434668 269922
rect 371601 269864 371606 269920
rect 371662 269864 376390 269920
rect 376446 269864 434668 269920
rect 371601 269862 434668 269864
rect 371601 269859 371667 269862
rect 376385 269859 376451 269862
rect 434662 269860 434668 269862
rect 434732 269860 434738 269924
rect 372153 269786 372219 269789
rect 431166 269786 431172 269788
rect 372153 269784 431172 269786
rect 372153 269728 372158 269784
rect 372214 269728 431172 269784
rect 372153 269726 431172 269728
rect 372153 269723 372219 269726
rect 431166 269724 431172 269726
rect 431236 269724 431242 269788
rect 217542 268364 217548 268428
rect 217612 268426 217618 268428
rect 229093 268426 229159 268429
rect 230381 268426 230447 268429
rect 217612 268424 230447 268426
rect 217612 268368 229098 268424
rect 229154 268368 230386 268424
rect 230442 268368 230447 268424
rect 217612 268366 230447 268368
rect 217612 268364 217618 268366
rect 229093 268363 229159 268366
rect 230381 268363 230447 268366
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 254146 480 254236
rect -960 254086 6930 254146
rect -960 253996 480 254086
rect 6870 254010 6930 254086
rect 54334 254010 54340 254012
rect 6870 253950 54340 254010
rect 54334 253948 54340 253950
rect 54404 253948 54410 254012
rect 339718 253404 339724 253468
rect 339788 253466 339794 253468
rect 340781 253466 340847 253469
rect 339788 253464 340847 253466
rect 339788 253408 340786 253464
rect 340842 253408 340847 253464
rect 339788 253406 340847 253408
rect 339788 253404 339794 253406
rect 340781 253403 340847 253406
rect 179638 253268 179644 253332
rect 179708 253330 179714 253332
rect 180149 253330 180215 253333
rect 179708 253328 180215 253330
rect 179708 253272 180154 253328
rect 180210 253272 180215 253328
rect 179708 253270 180215 253272
rect 179708 253268 179714 253270
rect 180149 253267 180215 253270
rect 499798 253268 499804 253332
rect 499868 253330 499874 253332
rect 500861 253330 500927 253333
rect 499868 253328 500927 253330
rect 499868 253272 500866 253328
rect 500922 253272 500927 253328
rect 499868 253270 500927 253272
rect 499868 253268 499874 253270
rect 500861 253267 500927 253270
rect 178534 253132 178540 253196
rect 178604 253194 178610 253196
rect 179321 253194 179387 253197
rect 178604 253192 179387 253194
rect 178604 253136 179326 253192
rect 179382 253136 179387 253192
rect 178604 253134 179387 253136
rect 178604 253132 178610 253134
rect 179321 253131 179387 253134
rect 350942 253132 350948 253196
rect 351012 253194 351018 253196
rect 351821 253194 351887 253197
rect 351012 253192 351887 253194
rect 351012 253136 351826 253192
rect 351882 253136 351887 253192
rect 351012 253134 351887 253136
rect 351012 253132 351018 253134
rect 351821 253131 351887 253134
rect 338430 252996 338436 253060
rect 338500 253058 338506 253060
rect 339401 253058 339467 253061
rect 338500 253056 339467 253058
rect 338500 253000 339406 253056
rect 339462 253000 339467 253056
rect 338500 252998 339467 253000
rect 338500 252996 338506 252998
rect 339401 252995 339467 252998
rect 498510 252724 498516 252788
rect 498580 252786 498586 252788
rect 499205 252786 499271 252789
rect 498580 252784 499271 252786
rect 498580 252728 499210 252784
rect 499266 252728 499271 252784
rect 498580 252726 499271 252728
rect 498580 252724 498586 252726
rect 499205 252723 499271 252726
rect 190862 252588 190868 252652
rect 190932 252650 190938 252652
rect 191741 252650 191807 252653
rect 510889 252652 510955 252653
rect 510838 252650 510844 252652
rect 190932 252648 191807 252650
rect 190932 252592 191746 252648
rect 191802 252592 191807 252648
rect 190932 252590 191807 252592
rect 510798 252590 510844 252650
rect 510908 252648 510955 252652
rect 510950 252592 510955 252648
rect 190932 252588 190938 252590
rect 191741 252587 191807 252590
rect 510838 252588 510844 252590
rect 510908 252588 510955 252592
rect 510889 252587 510955 252588
rect 57462 252452 57468 252516
rect 57532 252514 57538 252516
rect 60733 252514 60799 252517
rect 57532 252512 60799 252514
rect 57532 252456 60738 252512
rect 60794 252456 60799 252512
rect 57532 252454 60799 252456
rect 57532 252452 57538 252454
rect 60733 252451 60799 252454
rect 216622 252452 216628 252516
rect 216692 252514 216698 252516
rect 217358 252514 217364 252516
rect 216692 252454 217364 252514
rect 216692 252452 216698 252454
rect 217358 252452 217364 252454
rect 217428 252514 217434 252516
rect 217961 252514 218027 252517
rect 217428 252512 218027 252514
rect 217428 252456 217966 252512
rect 218022 252456 218027 252512
rect 217428 252454 218027 252456
rect 217428 252452 217434 252454
rect 217961 252451 218027 252454
rect 217542 251772 217548 251836
rect 217612 251834 217618 251836
rect 231853 251834 231919 251837
rect 217612 251832 231919 251834
rect 217612 251776 231858 251832
rect 231914 251776 231919 251832
rect 217612 251774 231919 251776
rect 217612 251772 217618 251774
rect 231853 251771 231919 251774
rect 377990 251772 377996 251836
rect 378060 251834 378066 251836
rect 389173 251834 389239 251837
rect 378060 251832 389239 251834
rect 378060 251776 389178 251832
rect 389234 251776 389239 251832
rect 378060 251774 389239 251776
rect 378060 251772 378066 251774
rect 389173 251771 389239 251774
rect 44950 251092 44956 251156
rect 45020 251154 45026 251156
rect 58525 251154 58591 251157
rect 45020 251152 58591 251154
rect 45020 251096 58530 251152
rect 58586 251096 58591 251152
rect 45020 251094 58591 251096
rect 45020 251092 45026 251094
rect 58525 251091 58591 251094
rect 44030 250956 44036 251020
rect 44100 251018 44106 251020
rect 53833 251018 53899 251021
rect 54385 251018 54451 251021
rect 44100 251016 54451 251018
rect 44100 250960 53838 251016
rect 53894 250960 54390 251016
rect 54446 250960 54451 251016
rect 44100 250958 54451 250960
rect 44100 250956 44106 250958
rect 53833 250955 53899 250958
rect 54385 250955 54451 250958
rect 198825 246258 198891 246261
rect 519261 246258 519327 246261
rect 196558 246256 198891 246258
rect 196558 246200 198830 246256
rect 198886 246200 198891 246256
rect 196558 246198 198891 246200
rect 196558 246190 196618 246198
rect 198825 246195 198891 246198
rect 516558 246256 519327 246258
rect 516558 246200 519266 246256
rect 519322 246200 519327 246256
rect 516558 246198 519327 246200
rect 516558 246190 516618 246198
rect 519261 246195 519327 246198
rect 356562 245714 356622 246190
rect 358997 245714 359063 245717
rect 359457 245714 359523 245717
rect 356562 245712 359523 245714
rect 356562 245656 359002 245712
rect 359058 245656 359462 245712
rect 359518 245656 359523 245712
rect 356562 245654 359523 245656
rect 358997 245651 359063 245654
rect 359457 245651 359523 245654
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 580257 232386 580323 232389
rect 583520 232386 584960 232476
rect 580257 232384 584960 232386
rect 580257 232328 580262 232384
rect 580318 232328 584960 232384
rect 580257 232326 584960 232328
rect 580257 232323 580323 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect 56685 204234 56751 204237
rect 57145 204234 57211 204237
rect 56685 204232 57211 204234
rect 56685 204176 56690 204232
rect 56746 204176 57150 204232
rect 57206 204176 57211 204232
rect 56685 204174 57211 204176
rect 56685 204171 56751 204174
rect 57145 204171 57211 204174
rect 57053 203962 57119 203965
rect 57881 203962 57947 203965
rect 217501 203962 217567 203965
rect 376937 203962 377003 203965
rect 57053 203960 60062 203962
rect 57053 203904 57058 203960
rect 57114 203904 57886 203960
rect 57942 203904 60062 203960
rect 57053 203902 60062 203904
rect 57053 203899 57119 203902
rect 57881 203899 57947 203902
rect 60002 203894 60062 203902
rect 217501 203960 219450 203962
rect 217501 203904 217506 203960
rect 217562 203924 219450 203960
rect 376937 203960 379530 203962
rect 217562 203904 220064 203924
rect 217501 203902 220064 203904
rect 217501 203899 217567 203902
rect 219390 203864 220064 203902
rect 376937 203904 376942 203960
rect 376998 203924 379530 203960
rect 376998 203904 380052 203924
rect 376937 203902 380052 203904
rect 376937 203899 377003 203902
rect 379470 203864 380052 203902
rect 56685 203010 56751 203013
rect 216857 203010 216923 203013
rect 217409 203010 217475 203013
rect 377857 203010 377923 203013
rect 378041 203010 378107 203013
rect 56685 203008 60062 203010
rect 56685 202952 56690 203008
rect 56746 202952 60062 203008
rect 56685 202950 60062 202952
rect 56685 202947 56751 202950
rect 60002 202942 60062 202950
rect 216857 203008 219450 203010
rect 216857 202952 216862 203008
rect 216918 202952 217414 203008
rect 217470 202972 219450 203008
rect 377857 203008 379530 203010
rect 217470 202952 220064 202972
rect 216857 202950 220064 202952
rect 216857 202947 216923 202950
rect 217409 202947 217475 202950
rect 219390 202912 220064 202950
rect 377857 202952 377862 203008
rect 377918 202952 378046 203008
rect 378102 202972 379530 203008
rect 378102 202952 380052 202972
rect 377857 202950 380052 202952
rect 377857 202947 377923 202950
rect 378041 202947 378107 202950
rect 379470 202912 380052 202950
rect -960 201922 480 202012
rect -960 201862 6930 201922
rect -960 201772 480 201862
rect 6870 201514 6930 201862
rect 51574 201514 51580 201516
rect 6870 201454 51580 201514
rect 51574 201452 51580 201454
rect 51644 201452 51650 201516
rect 57605 200834 57671 200837
rect 217593 200834 217659 200837
rect 377765 200834 377831 200837
rect 57605 200832 60062 200834
rect 57605 200776 57610 200832
rect 57666 200776 60062 200832
rect 57605 200774 60062 200776
rect 57605 200771 57671 200774
rect 60002 200766 60062 200774
rect 217593 200832 219450 200834
rect 217593 200776 217598 200832
rect 217654 200796 219450 200832
rect 377765 200832 379530 200834
rect 217654 200776 220064 200796
rect 217593 200774 220064 200776
rect 217593 200771 217659 200774
rect 219390 200736 220064 200774
rect 377765 200776 377770 200832
rect 377826 200796 379530 200832
rect 377826 200776 380052 200796
rect 377765 200774 380052 200776
rect 377765 200771 377831 200774
rect 379470 200736 380052 200774
rect 57329 199882 57395 199885
rect 217685 199882 217751 199885
rect 377581 199882 377647 199885
rect 57329 199880 60062 199882
rect 57329 199824 57334 199880
rect 57390 199824 60062 199880
rect 57329 199822 60062 199824
rect 57329 199819 57395 199822
rect 60002 199814 60062 199822
rect 217685 199880 219450 199882
rect 217685 199824 217690 199880
rect 217746 199844 219450 199880
rect 377581 199880 379530 199882
rect 217746 199824 220064 199844
rect 217685 199822 220064 199824
rect 217685 199819 217751 199822
rect 219390 199784 220064 199822
rect 377581 199824 377586 199880
rect 377642 199844 379530 199880
rect 377642 199824 380052 199844
rect 377581 199822 380052 199824
rect 377581 199819 377647 199822
rect 379470 199784 380052 199822
rect 57145 198794 57211 198797
rect 57329 198794 57395 198797
rect 57145 198792 57395 198794
rect 57145 198736 57150 198792
rect 57206 198736 57334 198792
rect 57390 198736 57395 198792
rect 57145 198734 57395 198736
rect 57145 198731 57211 198734
rect 57329 198731 57395 198734
rect 217409 198794 217475 198797
rect 217685 198794 217751 198797
rect 217409 198792 217751 198794
rect 217409 198736 217414 198792
rect 217470 198736 217690 198792
rect 217746 198736 217751 198792
rect 217409 198734 217751 198736
rect 217409 198731 217475 198734
rect 217685 198731 217751 198734
rect 376845 198794 376911 198797
rect 377581 198794 377647 198797
rect 376845 198792 377647 198794
rect 376845 198736 376850 198792
rect 376906 198736 377586 198792
rect 377642 198736 377647 198792
rect 376845 198734 377647 198736
rect 376845 198731 376911 198734
rect 377581 198731 377647 198734
rect 217869 198114 217935 198117
rect 377489 198114 377555 198117
rect 217869 198112 219450 198114
rect 217869 198056 217874 198112
rect 217930 198076 219450 198112
rect 377489 198112 379530 198114
rect 217930 198056 220064 198076
rect 217869 198054 220064 198056
rect 217869 198051 217935 198054
rect 57513 197434 57579 197437
rect 57697 197434 57763 197437
rect 60002 197434 60062 198046
rect 219390 198016 220064 198054
rect 377489 198056 377494 198112
rect 377550 198076 379530 198112
rect 377550 198056 380052 198076
rect 377489 198054 380052 198056
rect 377489 198051 377555 198054
rect 379470 198016 380052 198054
rect 57513 197432 60062 197434
rect 57513 197376 57518 197432
rect 57574 197376 57702 197432
rect 57758 197376 60062 197432
rect 57513 197374 60062 197376
rect 57513 197371 57579 197374
rect 57697 197371 57763 197374
rect 217777 197026 217843 197029
rect 377673 197026 377739 197029
rect 217777 197024 219450 197026
rect 217777 196968 217782 197024
rect 217838 196988 219450 197024
rect 377673 197024 379530 197026
rect 217838 196968 220064 196988
rect 217777 196966 220064 196968
rect 217777 196963 217843 196966
rect 57421 196346 57487 196349
rect 60002 196346 60062 196958
rect 219390 196928 220064 196966
rect 377673 196968 377678 197024
rect 377734 196988 379530 197024
rect 377734 196968 380052 196988
rect 377673 196966 380052 196968
rect 377673 196963 377739 196966
rect 379470 196928 380052 196966
rect 57421 196344 60062 196346
rect 57421 196288 57426 196344
rect 57482 196288 60062 196344
rect 57421 196286 60062 196288
rect 57421 196283 57487 196286
rect 56961 195258 57027 195261
rect 57789 195258 57855 195261
rect 217041 195258 217107 195261
rect 217685 195258 217751 195261
rect 377305 195258 377371 195261
rect 377581 195258 377647 195261
rect 56961 195256 60062 195258
rect 56961 195200 56966 195256
rect 57022 195200 57794 195256
rect 57850 195200 60062 195256
rect 56961 195198 60062 195200
rect 56961 195195 57027 195198
rect 57789 195195 57855 195198
rect 60002 195190 60062 195198
rect 217041 195256 219450 195258
rect 217041 195200 217046 195256
rect 217102 195200 217690 195256
rect 217746 195220 219450 195256
rect 377305 195256 379530 195258
rect 217746 195200 220064 195220
rect 217041 195198 220064 195200
rect 217041 195195 217107 195198
rect 217685 195195 217751 195198
rect 219390 195160 220064 195198
rect 377305 195200 377310 195256
rect 377366 195200 377586 195256
rect 377642 195220 379530 195256
rect 377642 195200 380052 195220
rect 377305 195198 380052 195200
rect 377305 195195 377371 195198
rect 377581 195195 377647 195198
rect 379470 195160 380052 195198
rect 580349 192538 580415 192541
rect 583520 192538 584960 192628
rect 580349 192536 584960 192538
rect 580349 192480 580354 192536
rect 580410 192480 584960 192536
rect 580349 192478 584960 192480
rect 580349 192475 580415 192478
rect 583520 192388 584960 192478
rect -960 188716 480 188956
rect 199285 186418 199351 186421
rect 359457 186418 359523 186421
rect 518893 186418 518959 186421
rect 519353 186418 519419 186421
rect 196558 186416 199351 186418
rect 196558 186360 199290 186416
rect 199346 186360 199351 186416
rect 196558 186358 199351 186360
rect 196558 186350 196618 186358
rect 199285 186355 199351 186358
rect 356562 186416 359523 186418
rect 356562 186360 359462 186416
rect 359518 186360 359523 186416
rect 356562 186358 359523 186360
rect 356562 186350 356622 186358
rect 359457 186355 359523 186358
rect 516558 186416 519419 186418
rect 516558 186360 518898 186416
rect 518954 186360 519358 186416
rect 519414 186360 519419 186416
rect 516558 186358 519419 186360
rect 516558 186350 516618 186358
rect 518893 186355 518959 186358
rect 519353 186355 519419 186358
rect 198733 184922 198799 184925
rect 199193 184922 199259 184925
rect 359273 184922 359339 184925
rect 359641 184922 359707 184925
rect 196558 184920 199259 184922
rect 196558 184864 198738 184920
rect 198794 184864 199198 184920
rect 199254 184864 199259 184920
rect 196558 184862 199259 184864
rect 196558 184718 196618 184862
rect 198733 184859 198799 184862
rect 199193 184859 199259 184862
rect 356562 184920 359707 184922
rect 356562 184864 359278 184920
rect 359334 184864 359646 184920
rect 359702 184864 359707 184920
rect 356562 184862 359707 184864
rect 356562 184718 356622 184862
rect 359273 184859 359339 184862
rect 359641 184859 359707 184862
rect 518985 184786 519051 184789
rect 520181 184786 520247 184789
rect 516558 184784 520247 184786
rect 516558 184728 518990 184784
rect 519046 184728 520186 184784
rect 520242 184728 520247 184784
rect 516558 184726 520247 184728
rect 516558 184718 516618 184726
rect 518985 184723 519051 184726
rect 520181 184723 520247 184726
rect 198733 183562 198799 183565
rect 198917 183562 198983 183565
rect 358905 183562 358971 183565
rect 359365 183562 359431 183565
rect 196558 183560 198983 183562
rect 196558 183504 198738 183560
rect 198794 183504 198922 183560
rect 198978 183504 198983 183560
rect 196558 183502 198983 183504
rect 196558 183358 196618 183502
rect 198733 183499 198799 183502
rect 198917 183499 198983 183502
rect 356562 183560 359431 183562
rect 356562 183504 358910 183560
rect 358966 183504 359370 183560
rect 359426 183504 359431 183560
rect 356562 183502 359431 183504
rect 356562 183358 356622 183502
rect 358905 183499 358971 183502
rect 359365 183499 359431 183502
rect 519445 183426 519511 183429
rect 520089 183426 520155 183429
rect 516558 183424 520155 183426
rect 516558 183368 519450 183424
rect 519506 183368 520094 183424
rect 520150 183368 520155 183424
rect 516558 183366 520155 183368
rect 516558 183358 516618 183366
rect 519445 183363 519511 183366
rect 520089 183363 520155 183366
rect 198917 182066 198983 182069
rect 199101 182066 199167 182069
rect 196558 182064 199167 182066
rect 196558 182008 198922 182064
rect 198978 182008 199106 182064
rect 199162 182008 199167 182064
rect 196558 182006 199167 182008
rect 196558 181862 196618 182006
rect 198917 182003 198983 182006
rect 199101 182003 199167 182006
rect 359181 181930 359247 181933
rect 519077 181930 519143 181933
rect 356562 181928 359247 181930
rect 356562 181872 359186 181928
rect 359242 181872 359247 181928
rect 356562 181870 359247 181872
rect 356562 181862 356622 181870
rect 359181 181867 359247 181870
rect 516558 181928 519143 181930
rect 516558 181872 519082 181928
rect 519138 181872 519143 181928
rect 516558 181870 519143 181872
rect 516558 181862 516618 181870
rect 519077 181867 519143 181870
rect 199009 180706 199075 180709
rect 359549 180706 359615 180709
rect 519169 180706 519235 180709
rect 196558 180704 199075 180706
rect 196558 180648 199014 180704
rect 199070 180648 199075 180704
rect 196558 180646 199075 180648
rect 196558 180638 196618 180646
rect 199009 180643 199075 180646
rect 356562 180704 359615 180706
rect 356562 180648 359554 180704
rect 359610 180648 359615 180704
rect 356562 180646 359615 180648
rect 356562 180638 356622 180646
rect 359549 180643 359615 180646
rect 516558 180704 519235 180706
rect 516558 180648 519174 180704
rect 519230 180648 519235 180704
rect 516558 180646 519235 180648
rect 516558 180638 516618 180646
rect 519169 180643 519235 180646
rect 359089 179482 359155 179485
rect 359549 179482 359615 179485
rect 359089 179480 359615 179482
rect 359089 179424 359094 179480
rect 359150 179424 359554 179480
rect 359610 179424 359615 179480
rect 359089 179422 359615 179424
rect 359089 179419 359155 179422
rect 359549 179419 359615 179422
rect 583520 179060 584960 179300
rect 58893 177578 58959 177581
rect 58893 177576 60062 177578
rect 58893 177520 58898 177576
rect 58954 177520 60062 177576
rect 58893 177518 60062 177520
rect 58893 177515 58959 177518
rect 60002 176966 60062 177518
rect 216673 177034 216739 177037
rect 377029 177034 377095 177037
rect 216673 177032 219450 177034
rect 216673 176976 216678 177032
rect 216734 176996 219450 177032
rect 377029 177032 379530 177034
rect 216734 176976 220064 176996
rect 216673 176974 220064 176976
rect 216673 176971 216739 176974
rect 219390 176936 220064 176974
rect 377029 176976 377034 177032
rect 377090 176996 379530 177032
rect 377090 176976 380052 176996
rect 377029 176974 380052 176976
rect 377029 176971 377095 176974
rect 379470 176936 380052 176974
rect -960 175796 480 176036
rect 57237 175402 57303 175405
rect 57881 175402 57947 175405
rect 216673 175402 216739 175405
rect 376937 175402 377003 175405
rect 57237 175400 60062 175402
rect 57237 175344 57242 175400
rect 57298 175344 57886 175400
rect 57942 175344 60062 175400
rect 57237 175342 60062 175344
rect 57237 175339 57303 175342
rect 57881 175339 57947 175342
rect 60002 175334 60062 175342
rect 216673 175400 219450 175402
rect 216673 175344 216678 175400
rect 216734 175364 219450 175400
rect 376937 175400 379530 175402
rect 216734 175344 220064 175364
rect 216673 175342 220064 175344
rect 216673 175339 216739 175342
rect 219390 175304 220064 175342
rect 376937 175344 376942 175400
rect 376998 175364 379530 175400
rect 376998 175344 380052 175364
rect 376937 175342 380052 175344
rect 376937 175339 377003 175342
rect 379470 175304 380052 175342
rect 56777 175130 56843 175133
rect 216673 175130 216739 175133
rect 377213 175130 377279 175133
rect 56777 175128 59554 175130
rect 56777 175072 56782 175128
rect 56838 175092 59554 175128
rect 216673 175128 219450 175130
rect 56838 175072 60032 175092
rect 56777 175070 60032 175072
rect 56777 175067 56843 175070
rect 59494 175032 60032 175070
rect 216673 175072 216678 175128
rect 216734 175092 219450 175128
rect 377213 175128 379530 175130
rect 216734 175072 220064 175092
rect 216673 175070 220064 175072
rect 216673 175067 216739 175070
rect 219390 175032 220064 175070
rect 377213 175072 377218 175128
rect 377274 175092 379530 175128
rect 377274 175072 380052 175092
rect 377213 175070 380052 175072
rect 377213 175067 377279 175070
rect 379470 175032 380052 175070
rect 219617 167106 219683 167109
rect 219934 167106 219940 167108
rect 219617 167104 219940 167106
rect 219617 167048 219622 167104
rect 219678 167048 219940 167104
rect 219617 167046 219940 167048
rect 219617 167043 219683 167046
rect 219934 167044 219940 167046
rect 220004 167044 220010 167108
rect 57646 166908 57652 166972
rect 57716 166970 57722 166972
rect 148358 166970 148364 166972
rect 57716 166910 148364 166970
rect 57716 166908 57722 166910
rect 148358 166908 148364 166910
rect 148428 166908 148434 166972
rect 206318 166908 206324 166972
rect 206388 166970 206394 166972
rect 206388 166910 313500 166970
rect 206388 166908 206394 166910
rect 138473 166836 138539 166837
rect 143533 166836 143599 166837
rect 57830 166772 57836 166836
rect 57900 166834 57906 166836
rect 57900 166774 122850 166834
rect 57900 166772 57906 166774
rect 98453 166700 98519 166701
rect 101029 166700 101095 166701
rect 105813 166700 105879 166701
rect 108205 166700 108271 166701
rect 98453 166698 98500 166700
rect 98408 166696 98500 166698
rect 98408 166640 98458 166696
rect 98408 166638 98500 166640
rect 98453 166636 98500 166638
rect 98564 166636 98570 166700
rect 101029 166698 101076 166700
rect 100984 166696 101076 166698
rect 100984 166640 101034 166696
rect 100984 166638 101076 166640
rect 101029 166636 101076 166638
rect 101140 166636 101146 166700
rect 105813 166698 105860 166700
rect 105768 166696 105860 166698
rect 105768 166640 105818 166696
rect 105768 166638 105860 166640
rect 105813 166636 105860 166638
rect 105924 166636 105930 166700
rect 108205 166698 108252 166700
rect 108160 166696 108252 166698
rect 108160 166640 108210 166696
rect 108160 166638 108252 166640
rect 108205 166636 108252 166638
rect 108316 166636 108322 166700
rect 122790 166698 122850 166774
rect 138472 166772 138478 166836
rect 138542 166834 138548 166836
rect 143504 166834 143510 166836
rect 138542 166774 138630 166834
rect 143442 166774 143510 166834
rect 143574 166832 143599 166836
rect 143594 166776 143599 166832
rect 138542 166772 138548 166774
rect 143504 166772 143510 166774
rect 143574 166772 143599 166776
rect 138473 166771 138539 166772
rect 143533 166771 143599 166772
rect 145925 166836 145991 166837
rect 298461 166836 298527 166837
rect 303521 166836 303587 166837
rect 313440 166836 313500 166910
rect 416037 166836 416103 166837
rect 418429 166836 418495 166837
rect 423397 166836 423463 166837
rect 425973 166836 426039 166837
rect 470961 166836 471027 166837
rect 473445 166836 473511 166837
rect 145925 166832 145958 166836
rect 146022 166834 146028 166836
rect 145925 166776 145930 166832
rect 145925 166772 145958 166776
rect 146022 166774 146082 166834
rect 146022 166772 146028 166774
rect 210550 166772 210556 166836
rect 210620 166834 210626 166836
rect 210620 166774 296730 166834
rect 210620 166772 210626 166774
rect 145925 166771 145991 166772
rect 163313 166700 163379 166701
rect 165889 166700 165955 166701
rect 288249 166700 288315 166701
rect 295885 166700 295951 166701
rect 140920 166698 140926 166700
rect 122790 166638 140926 166698
rect 140920 166636 140926 166638
rect 140990 166636 140996 166700
rect 163313 166696 163366 166700
rect 163430 166698 163436 166700
rect 163313 166640 163318 166696
rect 163313 166636 163366 166640
rect 163430 166638 163470 166698
rect 165889 166696 165950 166700
rect 165889 166640 165894 166696
rect 163430 166636 163436 166638
rect 165889 166636 165950 166640
rect 166014 166698 166020 166700
rect 166014 166638 166046 166698
rect 166014 166636 166020 166638
rect 208158 166636 208164 166700
rect 208228 166698 208234 166700
rect 208228 166638 277410 166698
rect 208228 166636 208234 166638
rect 98453 166635 98519 166636
rect 101029 166635 101095 166636
rect 105813 166635 105879 166636
rect 108205 166635 108271 166636
rect 163313 166635 163379 166636
rect 165889 166635 165955 166636
rect 113265 166564 113331 166565
rect 150893 166564 150959 166565
rect 153285 166564 153351 166565
rect 253565 166564 253631 166565
rect 265893 166564 265959 166565
rect 270861 166564 270927 166565
rect 113265 166560 113318 166564
rect 113382 166562 113388 166564
rect 150893 166562 150940 166564
rect 113265 166504 113270 166560
rect 113265 166500 113318 166504
rect 113382 166502 113422 166562
rect 150848 166560 150940 166562
rect 150848 166504 150898 166560
rect 150848 166502 150940 166504
rect 113382 166500 113388 166502
rect 150893 166500 150940 166502
rect 151004 166500 151010 166564
rect 153285 166562 153332 166564
rect 153240 166560 153332 166562
rect 153240 166504 153290 166560
rect 153240 166502 153332 166504
rect 153285 166500 153332 166502
rect 153396 166500 153402 166564
rect 253565 166562 253612 166564
rect 253520 166560 253612 166562
rect 253520 166504 253570 166560
rect 253520 166502 253612 166504
rect 253565 166500 253612 166502
rect 253676 166500 253682 166564
rect 265893 166562 265940 166564
rect 265848 166560 265940 166562
rect 265848 166504 265898 166560
rect 265848 166502 265940 166504
rect 265893 166500 265940 166502
rect 266004 166500 266010 166564
rect 270861 166562 270908 166564
rect 270816 166560 270908 166562
rect 270816 166504 270866 166560
rect 270816 166502 270908 166504
rect 270861 166500 270908 166502
rect 270972 166500 270978 166564
rect 277350 166562 277410 166638
rect 288249 166696 288278 166700
rect 288342 166698 288348 166700
rect 288249 166640 288254 166696
rect 288249 166636 288278 166640
rect 288342 166638 288406 166698
rect 295885 166696 295894 166700
rect 295958 166698 295964 166700
rect 296670 166698 296730 166774
rect 298461 166832 298478 166836
rect 298542 166834 298548 166836
rect 303504 166834 303510 166836
rect 298461 166776 298466 166832
rect 298461 166772 298478 166776
rect 298542 166774 298618 166834
rect 303430 166774 303510 166834
rect 303574 166832 303587 166836
rect 303582 166776 303587 166832
rect 298542 166772 298548 166774
rect 303504 166772 303510 166774
rect 303574 166772 303587 166776
rect 313432 166772 313438 166836
rect 313502 166772 313508 166836
rect 416037 166832 416046 166836
rect 416110 166834 416116 166836
rect 418429 166834 418476 166836
rect 416037 166776 416042 166832
rect 416037 166772 416046 166776
rect 416110 166774 416194 166834
rect 418384 166832 418476 166834
rect 418384 166776 418434 166832
rect 418384 166774 418476 166776
rect 416110 166772 416116 166774
rect 418429 166772 418476 166774
rect 418540 166772 418546 166836
rect 423397 166834 423444 166836
rect 423352 166832 423444 166834
rect 423352 166776 423402 166832
rect 423352 166774 423444 166776
rect 423397 166772 423444 166774
rect 423508 166772 423514 166836
rect 425973 166834 426020 166836
rect 425928 166832 426020 166834
rect 425928 166776 425978 166832
rect 425928 166774 426020 166776
rect 425973 166772 426020 166774
rect 426084 166772 426090 166836
rect 470961 166832 470990 166836
rect 471054 166834 471060 166836
rect 473432 166834 473438 166836
rect 470961 166776 470966 166832
rect 470961 166772 470990 166776
rect 471054 166774 471118 166834
rect 473354 166774 473438 166834
rect 473502 166832 473511 166836
rect 473506 166776 473511 166832
rect 471054 166772 471060 166774
rect 473432 166772 473438 166774
rect 473502 166772 473511 166776
rect 298461 166771 298527 166772
rect 303521 166771 303587 166772
rect 416037 166771 416103 166772
rect 418429 166771 418495 166772
rect 423397 166771 423463 166772
rect 425973 166771 426039 166772
rect 470961 166771 471027 166772
rect 473445 166771 473511 166772
rect 475837 166836 475903 166837
rect 478413 166836 478479 166837
rect 480897 166836 480963 166837
rect 475837 166832 475886 166836
rect 475950 166834 475956 166836
rect 475837 166776 475842 166832
rect 475837 166772 475886 166776
rect 475950 166774 475994 166834
rect 478413 166832 478470 166836
rect 478534 166834 478540 166836
rect 478413 166776 478418 166832
rect 475950 166772 475956 166774
rect 478413 166772 478470 166776
rect 478534 166774 478570 166834
rect 480897 166832 480918 166836
rect 480982 166834 480988 166836
rect 480897 166776 480902 166832
rect 478534 166772 478540 166774
rect 480897 166772 480918 166776
rect 480982 166774 481054 166834
rect 480982 166772 480988 166774
rect 475837 166771 475903 166772
rect 478413 166771 478479 166772
rect 480897 166771 480963 166772
rect 308489 166700 308555 166701
rect 315849 166700 315915 166701
rect 483381 166700 483447 166701
rect 485957 166700 486023 166701
rect 305952 166698 305958 166700
rect 295885 166640 295890 166696
rect 288342 166636 288348 166638
rect 295885 166636 295894 166640
rect 295958 166638 296042 166698
rect 296670 166638 305958 166698
rect 295958 166636 295964 166638
rect 305952 166636 305958 166638
rect 306022 166636 306028 166700
rect 308489 166696 308542 166700
rect 308606 166698 308612 166700
rect 308489 166640 308494 166696
rect 308489 166636 308542 166640
rect 308606 166638 308646 166698
rect 315849 166696 315886 166700
rect 315950 166698 315956 166700
rect 483360 166698 483366 166700
rect 315849 166640 315854 166696
rect 308606 166636 308612 166638
rect 315849 166636 315886 166640
rect 315950 166638 316006 166698
rect 483290 166638 483366 166698
rect 483430 166696 483447 166700
rect 485944 166698 485950 166700
rect 483442 166640 483447 166696
rect 315950 166636 315956 166638
rect 483360 166636 483366 166638
rect 483430 166636 483447 166640
rect 485866 166638 485950 166698
rect 486014 166696 486023 166700
rect 486018 166640 486023 166696
rect 485944 166636 485950 166638
rect 486014 166636 486023 166640
rect 288249 166635 288315 166636
rect 295885 166635 295951 166636
rect 308489 166635 308555 166636
rect 315849 166635 315915 166636
rect 483381 166635 483447 166636
rect 485957 166635 486023 166636
rect 413553 166564 413619 166565
rect 503253 166564 503319 166565
rect 290992 166562 290998 166564
rect 277350 166502 290998 166562
rect 290992 166500 290998 166502
rect 291062 166500 291068 166564
rect 413553 166560 413598 166564
rect 413662 166562 413668 166564
rect 503216 166562 503222 166564
rect 413553 166504 413558 166560
rect 413553 166500 413598 166504
rect 413662 166502 413710 166562
rect 503162 166502 503222 166562
rect 503286 166560 503319 166564
rect 503314 166504 503319 166560
rect 413662 166500 413668 166502
rect 503216 166500 503222 166502
rect 503286 166500 503319 166504
rect 113265 166499 113331 166500
rect 150893 166499 150959 166500
rect 153285 166499 153351 166500
rect 253565 166499 253631 166500
rect 265893 166499 265959 166500
rect 270861 166499 270927 166500
rect 413553 166499 413619 166500
rect 503253 166499 503319 166500
rect 96061 166292 96127 166293
rect 408125 166292 408191 166293
rect 428181 166292 428247 166293
rect 96061 166290 96108 166292
rect 96016 166288 96108 166290
rect 96016 166232 96066 166288
rect 96016 166230 96108 166232
rect 96061 166228 96108 166230
rect 96172 166228 96178 166292
rect 408125 166290 408172 166292
rect 408080 166288 408172 166290
rect 408080 166232 408130 166288
rect 408080 166230 408172 166232
rect 408125 166228 408172 166230
rect 408236 166228 408242 166292
rect 428181 166290 428228 166292
rect 428136 166288 428228 166290
rect 428136 166232 428186 166288
rect 428136 166230 428228 166232
rect 428181 166228 428228 166230
rect 428292 166228 428298 166292
rect 96061 166227 96127 166228
rect 408125 166227 408191 166228
rect 428181 166227 428247 166228
rect 583520 165732 584960 165972
rect 81433 165610 81499 165613
rect 81750 165610 81756 165612
rect 81433 165608 81756 165610
rect 81433 165552 81438 165608
rect 81494 165552 81756 165608
rect 81433 165550 81756 165552
rect 81433 165547 81499 165550
rect 81750 165548 81756 165550
rect 81820 165548 81826 165612
rect 84285 165610 84351 165613
rect 85430 165610 85436 165612
rect 84285 165608 85436 165610
rect 84285 165552 84290 165608
rect 84346 165552 85436 165608
rect 84285 165550 85436 165552
rect 84285 165547 84351 165550
rect 85430 165548 85436 165550
rect 85500 165548 85506 165612
rect 89897 165610 89963 165613
rect 90766 165610 90772 165612
rect 89897 165608 90772 165610
rect 89897 165552 89902 165608
rect 89958 165552 90772 165608
rect 89897 165550 90772 165552
rect 89897 165547 89963 165550
rect 90766 165548 90772 165550
rect 90836 165548 90842 165612
rect 91093 165610 91159 165613
rect 92422 165610 92428 165612
rect 91093 165608 92428 165610
rect 91093 165552 91098 165608
rect 91154 165552 92428 165608
rect 91093 165550 92428 165552
rect 91093 165547 91159 165550
rect 92422 165548 92428 165550
rect 92492 165548 92498 165612
rect 95233 165610 95299 165613
rect 99373 165612 99439 165613
rect 103513 165612 103579 165613
rect 95734 165610 95740 165612
rect 95233 165608 95740 165610
rect 95233 165552 95238 165608
rect 95294 165552 95740 165608
rect 95233 165550 95740 165552
rect 95233 165547 95299 165550
rect 95734 165548 95740 165550
rect 95804 165548 95810 165612
rect 99373 165608 99420 165612
rect 99484 165610 99490 165612
rect 99373 165552 99378 165608
rect 99373 165548 99420 165552
rect 99484 165550 99530 165610
rect 99484 165548 99490 165550
rect 103462 165548 103468 165612
rect 103532 165610 103579 165612
rect 109677 165612 109743 165613
rect 103532 165608 103624 165610
rect 103574 165552 103624 165608
rect 103532 165550 103624 165552
rect 109677 165608 109724 165612
rect 109788 165610 109794 165612
rect 110873 165610 110939 165613
rect 111149 165612 111215 165613
rect 111006 165610 111012 165612
rect 109677 165552 109682 165608
rect 103532 165548 103579 165550
rect 99373 165547 99439 165548
rect 103513 165547 103579 165548
rect 109677 165548 109724 165552
rect 109788 165550 109834 165610
rect 110873 165608 111012 165610
rect 110873 165552 110878 165608
rect 110934 165552 111012 165608
rect 110873 165550 111012 165552
rect 109788 165548 109794 165550
rect 109677 165547 109743 165548
rect 110873 165547 110939 165550
rect 111006 165548 111012 165550
rect 111076 165548 111082 165612
rect 111149 165608 111196 165612
rect 111260 165610 111266 165612
rect 111885 165610 111951 165613
rect 113541 165612 113607 165613
rect 115933 165612 115999 165613
rect 112110 165610 112116 165612
rect 111149 165552 111154 165608
rect 111149 165548 111196 165552
rect 111260 165550 111306 165610
rect 111885 165608 112116 165610
rect 111885 165552 111890 165608
rect 111946 165552 112116 165608
rect 111885 165550 112116 165552
rect 111260 165548 111266 165550
rect 111149 165547 111215 165548
rect 111885 165547 111951 165550
rect 112110 165548 112116 165550
rect 112180 165548 112186 165612
rect 113541 165608 113588 165612
rect 113652 165610 113658 165612
rect 113541 165552 113546 165608
rect 113541 165548 113588 165552
rect 113652 165550 113698 165610
rect 115933 165608 115980 165612
rect 116044 165610 116050 165612
rect 116393 165610 116459 165613
rect 116894 165610 116900 165612
rect 115933 165552 115938 165608
rect 113652 165548 113658 165550
rect 115933 165548 115980 165552
rect 116044 165550 116090 165610
rect 116393 165608 116900 165610
rect 116393 165552 116398 165608
rect 116454 165552 116900 165608
rect 116393 165550 116900 165552
rect 116044 165548 116050 165550
rect 113541 165547 113607 165548
rect 115933 165547 115999 165548
rect 116393 165547 116459 165550
rect 116894 165548 116900 165550
rect 116964 165548 116970 165612
rect 117865 165610 117931 165613
rect 118325 165612 118391 165613
rect 120901 165612 120967 165613
rect 123477 165612 123543 165613
rect 125869 165612 125935 165613
rect 117998 165610 118004 165612
rect 117865 165608 118004 165610
rect 117865 165552 117870 165608
rect 117926 165552 118004 165608
rect 117865 165550 118004 165552
rect 117865 165547 117931 165550
rect 117998 165548 118004 165550
rect 118068 165548 118074 165612
rect 118325 165608 118372 165612
rect 118436 165610 118442 165612
rect 118325 165552 118330 165608
rect 118325 165548 118372 165552
rect 118436 165550 118482 165610
rect 120901 165608 120948 165612
rect 121012 165610 121018 165612
rect 120901 165552 120906 165608
rect 118436 165548 118442 165550
rect 120901 165548 120948 165552
rect 121012 165550 121058 165610
rect 123477 165608 123524 165612
rect 123588 165610 123594 165612
rect 123477 165552 123482 165608
rect 121012 165548 121018 165550
rect 123477 165548 123524 165552
rect 123588 165550 123634 165610
rect 125869 165608 125916 165612
rect 125980 165610 125986 165612
rect 128353 165610 128419 165613
rect 128486 165610 128492 165612
rect 125869 165552 125874 165608
rect 123588 165548 123594 165550
rect 125869 165548 125916 165552
rect 125980 165550 126026 165610
rect 128353 165608 128492 165610
rect 128353 165552 128358 165608
rect 128414 165552 128492 165608
rect 128353 165550 128492 165552
rect 125980 165548 125986 165550
rect 118325 165547 118391 165548
rect 120901 165547 120967 165548
rect 123477 165547 123543 165548
rect 125869 165547 125935 165548
rect 128353 165547 128419 165550
rect 128486 165548 128492 165550
rect 128556 165548 128562 165612
rect 129733 165610 129799 165613
rect 130878 165610 130884 165612
rect 129733 165608 130884 165610
rect 129733 165552 129738 165608
rect 129794 165552 130884 165608
rect 129733 165550 130884 165552
rect 129733 165547 129799 165550
rect 130878 165548 130884 165550
rect 130948 165548 130954 165612
rect 132493 165610 132559 165613
rect 183185 165612 183251 165613
rect 133454 165610 133460 165612
rect 132493 165608 133460 165610
rect 132493 165552 132498 165608
rect 132554 165552 133460 165608
rect 132493 165550 133460 165552
rect 132493 165547 132559 165550
rect 133454 165548 133460 165550
rect 133524 165548 133530 165612
rect 183134 165610 183140 165612
rect 183094 165550 183140 165610
rect 183204 165608 183251 165612
rect 183246 165552 183251 165608
rect 183134 165548 183140 165550
rect 183204 165548 183251 165552
rect 183185 165547 183251 165548
rect 236085 165612 236151 165613
rect 236085 165608 236132 165612
rect 236196 165610 236202 165612
rect 238753 165610 238819 165613
rect 239622 165610 239628 165612
rect 236085 165552 236090 165608
rect 236085 165548 236132 165552
rect 236196 165550 236242 165610
rect 238753 165608 239628 165610
rect 238753 165552 238758 165608
rect 238814 165552 239628 165608
rect 238753 165550 239628 165552
rect 236196 165548 236202 165550
rect 236085 165547 236151 165548
rect 238753 165547 238819 165550
rect 239622 165548 239628 165550
rect 239692 165548 239698 165612
rect 242893 165610 242959 165613
rect 243118 165610 243124 165612
rect 242893 165608 243124 165610
rect 242893 165552 242898 165608
rect 242954 165552 243124 165608
rect 242893 165550 243124 165552
rect 242893 165547 242959 165550
rect 243118 165548 243124 165550
rect 243188 165548 243194 165612
rect 247125 165610 247191 165613
rect 247534 165610 247540 165612
rect 247125 165608 247540 165610
rect 247125 165552 247130 165608
rect 247186 165552 247540 165608
rect 247125 165550 247540 165552
rect 247125 165547 247191 165550
rect 247534 165548 247540 165550
rect 247604 165548 247610 165612
rect 258022 165548 258028 165612
rect 258092 165610 258098 165612
rect 258165 165610 258231 165613
rect 258092 165608 258231 165610
rect 258092 165552 258170 165608
rect 258226 165552 258231 165608
rect 258092 165550 258231 165552
rect 258092 165548 258098 165550
rect 258165 165547 258231 165550
rect 260833 165610 260899 165613
rect 273437 165612 273503 165613
rect 276013 165612 276079 165613
rect 278405 165612 278471 165613
rect 280797 165612 280863 165613
rect 285949 165612 286015 165613
rect 293309 165612 293375 165613
rect 300853 165612 300919 165613
rect 310973 165612 311039 165613
rect 325877 165612 325943 165613
rect 343265 165612 343331 165613
rect 261702 165610 261708 165612
rect 260833 165608 261708 165610
rect 260833 165552 260838 165608
rect 260894 165552 261708 165608
rect 260833 165550 261708 165552
rect 260833 165547 260899 165550
rect 261702 165548 261708 165550
rect 261772 165548 261778 165612
rect 273437 165608 273484 165612
rect 273548 165610 273554 165612
rect 273437 165552 273442 165608
rect 273437 165548 273484 165552
rect 273548 165550 273594 165610
rect 276013 165608 276060 165612
rect 276124 165610 276130 165612
rect 276013 165552 276018 165608
rect 273548 165548 273554 165550
rect 276013 165548 276060 165552
rect 276124 165550 276170 165610
rect 278405 165608 278452 165612
rect 278516 165610 278522 165612
rect 278405 165552 278410 165608
rect 276124 165548 276130 165550
rect 278405 165548 278452 165552
rect 278516 165550 278562 165610
rect 280797 165608 280844 165612
rect 280908 165610 280914 165612
rect 280797 165552 280802 165608
rect 278516 165548 278522 165550
rect 280797 165548 280844 165552
rect 280908 165550 280954 165610
rect 285949 165608 285996 165612
rect 286060 165610 286066 165612
rect 285949 165552 285954 165608
rect 280908 165548 280914 165550
rect 285949 165548 285996 165552
rect 286060 165550 286106 165610
rect 293309 165608 293356 165612
rect 293420 165610 293426 165612
rect 293309 165552 293314 165608
rect 286060 165548 286066 165550
rect 293309 165548 293356 165552
rect 293420 165550 293466 165610
rect 300853 165608 300900 165612
rect 300964 165610 300970 165612
rect 300853 165552 300858 165608
rect 293420 165548 293426 165550
rect 300853 165548 300900 165552
rect 300964 165550 301010 165610
rect 310973 165608 311020 165612
rect 311084 165610 311090 165612
rect 310973 165552 310978 165608
rect 300964 165548 300970 165550
rect 310973 165548 311020 165552
rect 311084 165550 311130 165610
rect 325877 165608 325924 165612
rect 325988 165610 325994 165612
rect 343214 165610 343220 165612
rect 325877 165552 325882 165608
rect 311084 165548 311090 165550
rect 325877 165548 325924 165552
rect 325988 165550 326034 165610
rect 343174 165550 343220 165610
rect 343284 165608 343331 165612
rect 343326 165552 343331 165608
rect 325988 165548 325994 165550
rect 343214 165548 343220 165550
rect 343284 165548 343331 165552
rect 273437 165547 273503 165548
rect 276013 165547 276079 165548
rect 278405 165547 278471 165548
rect 280797 165547 280863 165548
rect 285949 165547 286015 165548
rect 293309 165547 293375 165548
rect 300853 165547 300919 165548
rect 310973 165547 311039 165548
rect 325877 165547 325943 165548
rect 343265 165547 343331 165548
rect 397453 165610 397519 165613
rect 398230 165610 398236 165612
rect 397453 165608 398236 165610
rect 397453 165552 397458 165608
rect 397514 165552 398236 165608
rect 397453 165550 398236 165552
rect 397453 165547 397519 165550
rect 398230 165548 398236 165550
rect 398300 165548 398306 165612
rect 401593 165610 401659 165613
rect 401726 165610 401732 165612
rect 401593 165608 401732 165610
rect 401593 165552 401598 165608
rect 401654 165552 401732 165608
rect 401593 165550 401732 165552
rect 401593 165547 401659 165550
rect 401726 165548 401732 165550
rect 401796 165548 401802 165612
rect 404353 165610 404419 165613
rect 405406 165610 405412 165612
rect 404353 165608 405412 165610
rect 404353 165552 404358 165608
rect 404414 165552 405412 165608
rect 404353 165550 405412 165552
rect 404353 165547 404419 165550
rect 405406 165548 405412 165550
rect 405476 165548 405482 165612
rect 410425 165610 410491 165613
rect 410742 165610 410748 165612
rect 410425 165608 410748 165610
rect 410425 165552 410430 165608
rect 410486 165552 410748 165608
rect 410425 165550 410748 165552
rect 410425 165547 410491 165550
rect 410742 165548 410748 165550
rect 410812 165548 410818 165612
rect 415393 165610 415459 165613
rect 415894 165610 415900 165612
rect 415393 165608 415900 165610
rect 415393 165552 415398 165608
rect 415454 165552 415900 165608
rect 415393 165550 415900 165552
rect 415393 165547 415459 165550
rect 415894 165548 415900 165550
rect 415964 165548 415970 165612
rect 416865 165610 416931 165613
rect 416998 165610 417004 165612
rect 416865 165608 417004 165610
rect 416865 165552 416870 165608
rect 416926 165552 417004 165608
rect 416865 165550 417004 165552
rect 416865 165547 416931 165550
rect 416998 165548 417004 165550
rect 417068 165548 417074 165612
rect 418153 165610 418219 165613
rect 423765 165612 423831 165613
rect 419390 165610 419396 165612
rect 418153 165608 419396 165610
rect 418153 165552 418158 165608
rect 418214 165552 419396 165608
rect 418153 165550 419396 165552
rect 418153 165547 418219 165550
rect 419390 165548 419396 165550
rect 419460 165548 419466 165612
rect 423765 165610 423812 165612
rect 423720 165608 423812 165610
rect 423720 165552 423770 165608
rect 423720 165550 423812 165552
rect 423765 165548 423812 165550
rect 423876 165548 423882 165612
rect 426433 165610 426499 165613
rect 427486 165610 427492 165612
rect 426433 165608 427492 165610
rect 426433 165552 426438 165608
rect 426494 165552 427492 165608
rect 426433 165550 427492 165552
rect 423765 165547 423831 165548
rect 426433 165547 426499 165550
rect 427486 165548 427492 165550
rect 427556 165548 427562 165612
rect 433374 165548 433380 165612
rect 433444 165610 433450 165612
rect 434621 165610 434687 165613
rect 433444 165608 434687 165610
rect 433444 165552 434626 165608
rect 434682 165552 434687 165608
rect 433444 165550 434687 165552
rect 433444 165548 433450 165550
rect 434621 165547 434687 165550
rect 434805 165610 434871 165613
rect 435950 165610 435956 165612
rect 434805 165608 435956 165610
rect 434805 165552 434810 165608
rect 434866 165552 435956 165608
rect 434805 165550 435956 165552
rect 434805 165547 434871 165550
rect 435950 165548 435956 165550
rect 436020 165548 436026 165612
rect 437841 165610 437907 165613
rect 437974 165610 437980 165612
rect 437841 165608 437980 165610
rect 437841 165552 437846 165608
rect 437902 165552 437980 165608
rect 437841 165550 437980 165552
rect 437841 165547 437907 165550
rect 437974 165548 437980 165550
rect 438044 165548 438050 165612
rect 440233 165610 440299 165613
rect 440918 165610 440924 165612
rect 440233 165608 440924 165610
rect 440233 165552 440238 165608
rect 440294 165552 440924 165608
rect 440233 165550 440924 165552
rect 440233 165547 440299 165550
rect 440918 165548 440924 165550
rect 440988 165548 440994 165612
rect 442993 165610 443059 165613
rect 443494 165610 443500 165612
rect 442993 165608 443500 165610
rect 442993 165552 442998 165608
rect 443054 165552 443500 165608
rect 442993 165550 443500 165552
rect 442993 165547 443059 165550
rect 443494 165548 443500 165550
rect 443564 165548 443570 165612
rect 447317 165610 447383 165613
rect 448278 165610 448284 165612
rect 447317 165608 448284 165610
rect 447317 165552 447322 165608
rect 447378 165552 448284 165608
rect 447317 165550 448284 165552
rect 447317 165547 447383 165550
rect 448278 165548 448284 165550
rect 448348 165548 448354 165612
rect 449893 165610 449959 165613
rect 451038 165610 451044 165612
rect 449893 165608 451044 165610
rect 449893 165552 449898 165608
rect 449954 165552 451044 165608
rect 449893 165550 451044 165552
rect 449893 165547 449959 165550
rect 451038 165548 451044 165550
rect 451108 165548 451114 165612
rect 452653 165610 452719 165613
rect 453430 165610 453436 165612
rect 452653 165608 453436 165610
rect 452653 165552 452658 165608
rect 452714 165552 453436 165608
rect 452653 165550 453436 165552
rect 452653 165547 452719 165550
rect 453430 165548 453436 165550
rect 453500 165548 453506 165612
rect 455413 165610 455479 165613
rect 458357 165612 458423 165613
rect 455822 165610 455828 165612
rect 455413 165608 455828 165610
rect 455413 165552 455418 165608
rect 455474 165552 455828 165608
rect 455413 165550 455828 165552
rect 455413 165547 455479 165550
rect 455822 165548 455828 165550
rect 455892 165548 455898 165612
rect 458357 165608 458404 165612
rect 458468 165610 458474 165612
rect 458357 165552 458362 165608
rect 458357 165548 458404 165552
rect 458468 165550 458514 165610
rect 458468 165548 458474 165550
rect 458357 165547 458423 165548
rect 50613 165474 50679 165477
rect 155902 165474 155908 165476
rect 50613 165472 155908 165474
rect 50613 165416 50618 165472
rect 50674 165416 155908 165472
rect 50613 165414 155908 165416
rect 50613 165411 50679 165414
rect 155902 165412 155908 165414
rect 155972 165412 155978 165476
rect 203517 165474 203583 165477
rect 318374 165474 318380 165476
rect 203517 165472 318380 165474
rect 203517 165416 203522 165472
rect 203578 165416 318380 165472
rect 203517 165414 318380 165416
rect 203517 165411 203583 165414
rect 318374 165412 318380 165414
rect 318444 165412 318450 165476
rect 376201 165474 376267 165477
rect 468518 165474 468524 165476
rect 376201 165472 468524 165474
rect 376201 165416 376206 165472
rect 376262 165416 468524 165472
rect 376201 165414 468524 165416
rect 376201 165411 376267 165414
rect 468518 165412 468524 165414
rect 468588 165412 468594 165476
rect 53281 165338 53347 165341
rect 158478 165338 158484 165340
rect 53281 165336 158484 165338
rect 53281 165280 53286 165336
rect 53342 165280 158484 165336
rect 53281 165278 158484 165280
rect 53281 165275 53347 165278
rect 158478 165276 158484 165278
rect 158548 165276 158554 165340
rect 216254 165276 216260 165340
rect 216324 165338 216330 165340
rect 283414 165338 283420 165340
rect 216324 165278 283420 165338
rect 216324 165276 216330 165278
rect 283414 165276 283420 165278
rect 283484 165276 283490 165340
rect 374821 165338 374887 165341
rect 465942 165338 465948 165340
rect 374821 165336 465948 165338
rect 374821 165280 374826 165336
rect 374882 165280 465948 165336
rect 374821 165278 465948 165280
rect 374821 165275 374887 165278
rect 465942 165276 465948 165278
rect 466012 165276 466018 165340
rect 56317 165202 56383 165205
rect 135846 165202 135852 165204
rect 56317 165200 135852 165202
rect 56317 165144 56322 165200
rect 56378 165144 135852 165200
rect 56317 165142 135852 165144
rect 56317 165139 56383 165142
rect 135846 165140 135852 165142
rect 135916 165140 135922 165204
rect 200798 165140 200804 165204
rect 200868 165202 200874 165204
rect 260966 165202 260972 165204
rect 200868 165142 260972 165202
rect 200868 165140 200874 165142
rect 260966 165140 260972 165142
rect 261036 165140 261042 165204
rect 263593 165202 263659 165205
rect 263726 165202 263732 165204
rect 263593 165200 263732 165202
rect 263593 165144 263598 165200
rect 263654 165144 263732 165200
rect 263593 165142 263732 165144
rect 263593 165139 263659 165142
rect 263726 165140 263732 165142
rect 263796 165140 263802 165204
rect 265382 165140 265388 165204
rect 265452 165202 265458 165204
rect 266261 165202 266327 165205
rect 265452 165200 266327 165202
rect 265452 165144 266266 165200
rect 266322 165144 266327 165200
rect 265452 165142 266327 165144
rect 265452 165140 265458 165142
rect 266261 165139 266327 165142
rect 271873 165202 271939 165205
rect 272190 165202 272196 165204
rect 271873 165200 272196 165202
rect 271873 165144 271878 165200
rect 271934 165144 272196 165200
rect 271873 165142 272196 165144
rect 271873 165139 271939 165142
rect 272190 165140 272196 165142
rect 272260 165140 272266 165204
rect 275277 165202 275343 165205
rect 275686 165202 275692 165204
rect 275277 165200 275692 165202
rect 275277 165144 275282 165200
rect 275338 165144 275692 165200
rect 275277 165142 275692 165144
rect 275277 165139 275343 165142
rect 275686 165140 275692 165142
rect 275756 165140 275762 165204
rect 279182 165140 279188 165204
rect 279252 165202 279258 165204
rect 280061 165202 280127 165205
rect 279252 165200 280127 165202
rect 279252 165144 280066 165200
rect 280122 165144 280127 165200
rect 279252 165142 280127 165144
rect 279252 165140 279258 165142
rect 280061 165139 280127 165142
rect 378910 165140 378916 165204
rect 378980 165202 378986 165204
rect 463550 165202 463556 165204
rect 378980 165142 463556 165202
rect 378980 165140 378986 165142
rect 463550 165140 463556 165142
rect 463620 165140 463626 165204
rect 47894 165004 47900 165068
rect 47964 165066 47970 165068
rect 93710 165066 93716 165068
rect 47964 165006 93716 165066
rect 47964 165004 47970 165006
rect 93710 165004 93716 165006
rect 93780 165004 93786 165068
rect 118877 165066 118943 165069
rect 183461 165068 183527 165069
rect 119102 165066 119108 165068
rect 118877 165064 119108 165066
rect 118877 165008 118882 165064
rect 118938 165008 119108 165064
rect 118877 165006 119108 165008
rect 118877 165003 118943 165006
rect 119102 165004 119108 165006
rect 119172 165004 119178 165068
rect 183461 165064 183508 165068
rect 183572 165066 183578 165068
rect 267733 165066 267799 165069
rect 268326 165066 268332 165068
rect 183461 165008 183466 165064
rect 183461 165004 183508 165008
rect 183572 165006 183618 165066
rect 267733 165064 268332 165066
rect 267733 165008 267738 165064
rect 267794 165008 268332 165064
rect 267733 165006 268332 165008
rect 183572 165004 183578 165006
rect 183461 165003 183527 165004
rect 267733 165003 267799 165006
rect 268326 165004 268332 165006
rect 268396 165004 268402 165068
rect 437749 165066 437815 165069
rect 438526 165066 438532 165068
rect 437749 165064 438532 165066
rect 437749 165008 437754 165064
rect 437810 165008 438532 165064
rect 437749 165006 438532 165008
rect 437749 165003 437815 165006
rect 438526 165004 438532 165006
rect 438596 165004 438602 165068
rect 445753 165066 445819 165069
rect 445886 165066 445892 165068
rect 445753 165064 445892 165066
rect 445753 165008 445758 165064
rect 445814 165008 445892 165064
rect 445753 165006 445892 165008
rect 445753 165003 445819 165006
rect 445886 165004 445892 165006
rect 445956 165004 445962 165068
rect 104893 164930 104959 164933
rect 105302 164930 105308 164932
rect 104893 164928 105308 164930
rect 104893 164872 104898 164928
rect 104954 164872 105308 164928
rect 104893 164870 105308 164872
rect 104893 164867 104959 164870
rect 105302 164868 105308 164870
rect 105372 164868 105378 164932
rect 106406 164868 106412 164932
rect 106476 164930 106482 164932
rect 107561 164930 107627 164933
rect 106476 164928 107627 164930
rect 106476 164872 107566 164928
rect 107622 164872 107627 164928
rect 106476 164870 107627 164872
rect 106476 164868 106482 164870
rect 107561 164867 107627 164870
rect 114461 164932 114527 164933
rect 114461 164928 114508 164932
rect 114572 164930 114578 164932
rect 247033 164930 247099 164933
rect 248270 164930 248276 164932
rect 114461 164872 114466 164928
rect 114461 164868 114508 164872
rect 114572 164870 114618 164930
rect 247033 164928 248276 164930
rect 247033 164872 247038 164928
rect 247094 164872 248276 164928
rect 247033 164870 248276 164872
rect 114572 164868 114578 164870
rect 114461 164867 114527 164868
rect 247033 164867 247099 164870
rect 248270 164868 248276 164870
rect 248340 164868 248346 164932
rect 249793 164930 249859 164933
rect 250662 164930 250668 164932
rect 249793 164928 250668 164930
rect 249793 164872 249798 164928
rect 249854 164872 250668 164928
rect 249793 164870 250668 164872
rect 249793 164867 249859 164870
rect 250662 164868 250668 164870
rect 250732 164868 250738 164932
rect 255313 164930 255379 164933
rect 256182 164930 256188 164932
rect 255313 164928 256188 164930
rect 255313 164872 255318 164928
rect 255374 164872 256188 164928
rect 255313 164870 256188 164872
rect 255313 164867 255379 164870
rect 256182 164868 256188 164870
rect 256252 164868 256258 164932
rect 258073 164930 258139 164933
rect 258390 164930 258396 164932
rect 258073 164928 258396 164930
rect 258073 164872 258078 164928
rect 258134 164872 258396 164928
rect 258073 164870 258396 164872
rect 258073 164867 258139 164870
rect 258390 164868 258396 164870
rect 258460 164868 258466 164932
rect 343398 164868 343404 164932
rect 343468 164930 343474 164932
rect 343541 164930 343607 164933
rect 343468 164928 343607 164930
rect 343468 164872 343546 164928
rect 343602 164872 343607 164928
rect 343468 164870 343607 164872
rect 343468 164868 343474 164870
rect 343541 164867 343607 164870
rect 420913 164930 420979 164933
rect 421046 164930 421052 164932
rect 420913 164928 421052 164930
rect 420913 164872 420918 164928
rect 420974 164872 421052 164928
rect 420913 164870 421052 164872
rect 420913 164867 420979 164870
rect 421046 164868 421052 164870
rect 421116 164868 421122 164932
rect 433333 164930 433399 164933
rect 433558 164930 433564 164932
rect 433333 164928 433564 164930
rect 433333 164872 433338 164928
rect 433394 164872 433564 164928
rect 433333 164870 433564 164872
rect 433333 164867 433399 164870
rect 433558 164868 433564 164870
rect 433628 164868 433634 164932
rect 88333 164796 88399 164797
rect 88333 164794 88380 164796
rect 88288 164792 88380 164794
rect 88288 164736 88338 164792
rect 88288 164734 88380 164736
rect 88333 164732 88380 164734
rect 88444 164732 88450 164796
rect 106273 164794 106339 164797
rect 107510 164794 107516 164796
rect 106273 164792 107516 164794
rect 106273 164736 106278 164792
rect 106334 164736 107516 164792
rect 106273 164734 107516 164736
rect 88333 164731 88399 164732
rect 106273 164731 106339 164734
rect 107510 164732 107516 164734
rect 107580 164732 107586 164796
rect 202454 164732 202460 164796
rect 202524 164794 202530 164796
rect 323342 164794 323348 164796
rect 202524 164734 323348 164794
rect 202524 164732 202530 164734
rect 323342 164732 323348 164734
rect 323412 164732 323418 164796
rect 363781 164794 363847 164797
rect 460974 164794 460980 164796
rect 363781 164792 460980 164794
rect 363781 164736 363786 164792
rect 363842 164736 460980 164792
rect 363781 164734 460980 164736
rect 363781 164731 363847 164734
rect 460974 164732 460980 164734
rect 461044 164732 461050 164796
rect 49233 164658 49299 164661
rect 160870 164658 160876 164660
rect 49233 164656 160876 164658
rect 49233 164600 49238 164656
rect 49294 164600 160876 164656
rect 49233 164598 160876 164600
rect 49233 164595 49299 164598
rect 160870 164596 160876 164598
rect 160940 164596 160946 164660
rect 433333 164658 433399 164661
rect 434662 164658 434668 164660
rect 433333 164656 434668 164658
rect 433333 164600 433338 164656
rect 433394 164600 434668 164656
rect 433333 164598 434668 164600
rect 433333 164595 433399 164598
rect 434662 164596 434668 164598
rect 434732 164596 434738 164660
rect 503294 164596 503300 164660
rect 503364 164658 503370 164660
rect 503621 164658 503687 164661
rect 503364 164656 503687 164658
rect 503364 164600 503626 164656
rect 503682 164600 503687 164656
rect 503364 164598 503687 164600
rect 503364 164596 503370 164598
rect 503621 164595 503687 164598
rect 100753 164524 100819 164525
rect 100702 164460 100708 164524
rect 100772 164522 100819 164524
rect 107745 164522 107811 164525
rect 108614 164522 108620 164524
rect 100772 164520 100864 164522
rect 100814 164464 100864 164520
rect 100772 164462 100864 164464
rect 107745 164520 108620 164522
rect 107745 164464 107750 164520
rect 107806 164464 108620 164520
rect 107745 164462 108620 164464
rect 100772 164460 100819 164462
rect 100753 164459 100819 164460
rect 107745 164459 107811 164462
rect 108614 164460 108620 164462
rect 108684 164460 108690 164524
rect 115790 164460 115796 164524
rect 115860 164522 115866 164524
rect 116025 164522 116091 164525
rect 115860 164520 116091 164522
rect 115860 164464 116030 164520
rect 116086 164464 116091 164520
rect 115860 164462 116091 164464
rect 115860 164460 115866 164462
rect 116025 164459 116091 164462
rect 76005 164386 76071 164389
rect 244365 164388 244431 164389
rect 77150 164386 77156 164388
rect 76005 164384 77156 164386
rect 76005 164328 76010 164384
rect 76066 164328 77156 164384
rect 76005 164326 77156 164328
rect 76005 164323 76071 164326
rect 77150 164324 77156 164326
rect 77220 164324 77226 164388
rect 244365 164384 244412 164388
rect 244476 164386 244482 164388
rect 251265 164386 251331 164389
rect 252318 164386 252324 164388
rect 244365 164328 244370 164384
rect 244365 164324 244412 164328
rect 244476 164326 244522 164386
rect 251265 164384 252324 164386
rect 251265 164328 251270 164384
rect 251326 164328 252324 164384
rect 251265 164326 252324 164328
rect 244476 164324 244482 164326
rect 244365 164323 244431 164324
rect 251265 164323 251331 164326
rect 252318 164324 252324 164326
rect 252388 164324 252394 164388
rect 256693 164386 256759 164389
rect 256918 164386 256924 164388
rect 256693 164384 256924 164386
rect 256693 164328 256698 164384
rect 256754 164328 256924 164384
rect 256693 164326 256924 164328
rect 256693 164323 256759 164326
rect 256918 164324 256924 164326
rect 256988 164324 256994 164388
rect 259545 164386 259611 164389
rect 260598 164386 260604 164388
rect 259545 164384 260604 164386
rect 259545 164328 259550 164384
rect 259606 164328 260604 164384
rect 259545 164326 260604 164328
rect 259545 164323 259611 164326
rect 260598 164324 260604 164326
rect 260668 164324 260674 164388
rect 266537 164386 266603 164389
rect 267590 164386 267596 164388
rect 266537 164384 267596 164386
rect 266537 164328 266542 164384
rect 266598 164328 267596 164384
rect 266537 164326 267596 164328
rect 266537 164323 266603 164326
rect 267590 164324 267596 164326
rect 267660 164324 267666 164388
rect 273805 164386 273871 164389
rect 274398 164386 274404 164388
rect 273805 164384 274404 164386
rect 273805 164328 273810 164384
rect 273866 164328 274404 164384
rect 273805 164326 274404 164328
rect 273805 164323 273871 164326
rect 274398 164324 274404 164326
rect 274468 164324 274474 164388
rect 396165 164386 396231 164389
rect 397126 164386 397132 164388
rect 396165 164384 397132 164386
rect 396165 164328 396170 164384
rect 396226 164328 397132 164384
rect 396165 164326 397132 164328
rect 396165 164323 396231 164326
rect 397126 164324 397132 164326
rect 397196 164324 397202 164388
rect 402973 164386 403039 164389
rect 404118 164386 404124 164388
rect 402973 164384 404124 164386
rect 402973 164328 402978 164384
rect 403034 164328 404124 164384
rect 402973 164326 404124 164328
rect 402973 164323 403039 164326
rect 404118 164324 404124 164326
rect 404188 164324 404194 164388
rect 411345 164386 411411 164389
rect 412398 164386 412404 164388
rect 411345 164384 412404 164386
rect 411345 164328 411350 164384
rect 411406 164328 412404 164384
rect 411345 164326 412404 164328
rect 411345 164323 411411 164326
rect 412398 164324 412404 164326
rect 412468 164324 412474 164388
rect 429285 164386 429351 164389
rect 429694 164386 429700 164388
rect 429285 164384 429700 164386
rect 429285 164328 429290 164384
rect 429346 164328 429700 164384
rect 429285 164326 429700 164328
rect 429285 164323 429351 164326
rect 429694 164324 429700 164326
rect 429764 164324 429770 164388
rect 430665 164386 430731 164389
rect 431166 164386 431172 164388
rect 430665 164384 431172 164386
rect 430665 164328 430670 164384
rect 430726 164328 431172 164384
rect 430665 164326 431172 164328
rect 430665 164323 430731 164326
rect 431166 164324 431172 164326
rect 431236 164324 431242 164388
rect 57462 164188 57468 164252
rect 57532 164250 57538 164252
rect 59445 164250 59511 164253
rect 57532 164248 59511 164250
rect 57532 164192 59450 164248
rect 59506 164192 59511 164248
rect 57532 164190 59511 164192
rect 57532 164188 57538 164190
rect 59445 164187 59511 164190
rect 75913 164250 75979 164253
rect 76046 164250 76052 164252
rect 75913 164248 76052 164250
rect 75913 164192 75918 164248
rect 75974 164192 76052 164248
rect 75913 164190 76052 164192
rect 75913 164187 75979 164190
rect 76046 164188 76052 164190
rect 76116 164188 76122 164252
rect 77293 164250 77359 164253
rect 78254 164250 78260 164252
rect 77293 164248 78260 164250
rect 77293 164192 77298 164248
rect 77354 164192 78260 164248
rect 77293 164190 78260 164192
rect 77293 164187 77359 164190
rect 78254 164188 78260 164190
rect 78324 164188 78330 164252
rect 78673 164250 78739 164253
rect 79542 164250 79548 164252
rect 78673 164248 79548 164250
rect 78673 164192 78678 164248
rect 78734 164192 79548 164248
rect 78673 164190 79548 164192
rect 78673 164187 78739 164190
rect 79542 164188 79548 164190
rect 79612 164188 79618 164252
rect 80053 164250 80119 164253
rect 80462 164250 80468 164252
rect 80053 164248 80468 164250
rect 80053 164192 80058 164248
rect 80114 164192 80468 164248
rect 80053 164190 80468 164192
rect 80053 164187 80119 164190
rect 80462 164188 80468 164190
rect 80532 164188 80538 164252
rect 82813 164250 82879 164253
rect 84193 164252 84259 164253
rect 83038 164250 83044 164252
rect 82813 164248 83044 164250
rect 82813 164192 82818 164248
rect 82874 164192 83044 164248
rect 82813 164190 83044 164192
rect 82813 164187 82879 164190
rect 83038 164188 83044 164190
rect 83108 164188 83114 164252
rect 84142 164188 84148 164252
rect 84212 164250 84259 164252
rect 85573 164250 85639 164253
rect 86534 164250 86540 164252
rect 84212 164248 84304 164250
rect 84254 164192 84304 164248
rect 84212 164190 84304 164192
rect 85573 164248 86540 164250
rect 85573 164192 85578 164248
rect 85634 164192 86540 164248
rect 85573 164190 86540 164192
rect 84212 164188 84259 164190
rect 84193 164187 84259 164188
rect 85573 164187 85639 164190
rect 86534 164188 86540 164190
rect 86604 164188 86610 164252
rect 86953 164250 87019 164253
rect 87638 164250 87644 164252
rect 86953 164248 87644 164250
rect 86953 164192 86958 164248
rect 87014 164192 87644 164248
rect 86953 164190 87644 164192
rect 86953 164187 87019 164190
rect 87638 164188 87644 164190
rect 87708 164188 87714 164252
rect 88425 164250 88491 164253
rect 88742 164250 88748 164252
rect 88425 164248 88748 164250
rect 88425 164192 88430 164248
rect 88486 164192 88748 164248
rect 88425 164190 88748 164192
rect 88425 164187 88491 164190
rect 88742 164188 88748 164190
rect 88812 164188 88818 164252
rect 89805 164250 89871 164253
rect 90030 164250 90036 164252
rect 89805 164248 90036 164250
rect 89805 164192 89810 164248
rect 89866 164192 90036 164248
rect 89805 164190 90036 164192
rect 89805 164187 89871 164190
rect 90030 164188 90036 164190
rect 90100 164188 90106 164252
rect 91185 164250 91251 164253
rect 91318 164250 91324 164252
rect 91185 164248 91324 164250
rect 91185 164192 91190 164248
rect 91246 164192 91324 164248
rect 91185 164190 91324 164192
rect 91185 164187 91251 164190
rect 91318 164188 91324 164190
rect 91388 164188 91394 164252
rect 92473 164250 92539 164253
rect 93342 164250 93348 164252
rect 92473 164248 93348 164250
rect 92473 164192 92478 164248
rect 92534 164192 93348 164248
rect 92473 164190 93348 164192
rect 92473 164187 92539 164190
rect 93342 164188 93348 164190
rect 93412 164188 93418 164252
rect 93853 164250 93919 164253
rect 94446 164250 94452 164252
rect 93853 164248 94452 164250
rect 93853 164192 93858 164248
rect 93914 164192 94452 164248
rect 93853 164190 94452 164192
rect 93853 164187 93919 164190
rect 94446 164188 94452 164190
rect 94516 164188 94522 164252
rect 96613 164250 96679 164253
rect 97022 164250 97028 164252
rect 96613 164248 97028 164250
rect 96613 164192 96618 164248
rect 96674 164192 97028 164248
rect 96613 164190 97028 164192
rect 96613 164187 96679 164190
rect 97022 164188 97028 164190
rect 97092 164188 97098 164252
rect 97993 164250 98059 164253
rect 98126 164250 98132 164252
rect 97993 164248 98132 164250
rect 97993 164192 97998 164248
rect 98054 164192 98132 164248
rect 97993 164190 98132 164192
rect 97993 164187 98059 164190
rect 98126 164188 98132 164190
rect 98196 164188 98202 164252
rect 100753 164250 100819 164253
rect 101806 164250 101812 164252
rect 100753 164248 101812 164250
rect 100753 164192 100758 164248
rect 100814 164192 101812 164248
rect 100753 164190 101812 164192
rect 100753 164187 100819 164190
rect 101806 164188 101812 164190
rect 101876 164188 101882 164252
rect 102133 164250 102199 164253
rect 102726 164250 102732 164252
rect 102133 164248 102732 164250
rect 102133 164192 102138 164248
rect 102194 164192 102732 164248
rect 102133 164190 102732 164192
rect 102133 164187 102199 164190
rect 102726 164188 102732 164190
rect 102796 164188 102802 164252
rect 103605 164250 103671 164253
rect 103830 164250 103836 164252
rect 103605 164248 103836 164250
rect 103605 164192 103610 164248
rect 103666 164192 103836 164248
rect 103605 164190 103836 164192
rect 103605 164187 103671 164190
rect 103830 164188 103836 164190
rect 103900 164188 103906 164252
rect 235993 164250 236059 164253
rect 237046 164250 237052 164252
rect 235993 164248 237052 164250
rect 235993 164192 235998 164248
rect 236054 164192 237052 164248
rect 235993 164190 237052 164192
rect 235993 164187 236059 164190
rect 237046 164188 237052 164190
rect 237116 164188 237122 164252
rect 237373 164250 237439 164253
rect 238150 164250 238156 164252
rect 237373 164248 238156 164250
rect 237373 164192 237378 164248
rect 237434 164192 238156 164248
rect 237373 164190 238156 164192
rect 237373 164187 237439 164190
rect 238150 164188 238156 164190
rect 238220 164188 238226 164252
rect 240133 164250 240199 164253
rect 240542 164250 240548 164252
rect 240133 164248 240548 164250
rect 240133 164192 240138 164248
rect 240194 164192 240548 164248
rect 240133 164190 240548 164192
rect 240133 164187 240199 164190
rect 240542 164188 240548 164190
rect 240612 164188 240618 164252
rect 241513 164250 241579 164253
rect 241646 164250 241652 164252
rect 241513 164248 241652 164250
rect 241513 164192 241518 164248
rect 241574 164192 241652 164248
rect 241513 164190 241652 164192
rect 241513 164187 241579 164190
rect 241646 164188 241652 164190
rect 241716 164188 241722 164252
rect 244273 164250 244339 164253
rect 245326 164250 245332 164252
rect 244273 164248 245332 164250
rect 244273 164192 244278 164248
rect 244334 164192 245332 164248
rect 244273 164190 245332 164192
rect 244273 164187 244339 164190
rect 245326 164188 245332 164190
rect 245396 164188 245402 164252
rect 245653 164250 245719 164253
rect 246430 164250 246436 164252
rect 245653 164248 246436 164250
rect 245653 164192 245658 164248
rect 245714 164192 246436 164248
rect 245653 164190 246436 164192
rect 245653 164187 245719 164190
rect 246430 164188 246436 164190
rect 246500 164188 246506 164252
rect 248413 164250 248479 164253
rect 248638 164250 248644 164252
rect 248413 164248 248644 164250
rect 248413 164192 248418 164248
rect 248474 164192 248644 164248
rect 248413 164190 248644 164192
rect 248413 164187 248479 164190
rect 248638 164188 248644 164190
rect 248708 164188 248714 164252
rect 249885 164250 249951 164253
rect 251173 164252 251239 164253
rect 250110 164250 250116 164252
rect 249885 164248 250116 164250
rect 249885 164192 249890 164248
rect 249946 164192 250116 164248
rect 249885 164190 250116 164192
rect 249885 164187 249951 164190
rect 250110 164188 250116 164190
rect 250180 164188 250186 164252
rect 251173 164250 251220 164252
rect 251128 164248 251220 164250
rect 251128 164192 251178 164248
rect 251128 164190 251220 164192
rect 251173 164188 251220 164190
rect 251284 164188 251290 164252
rect 252553 164250 252619 164253
rect 253422 164250 253428 164252
rect 252553 164248 253428 164250
rect 252553 164192 252558 164248
rect 252614 164192 253428 164248
rect 252553 164190 253428 164192
rect 251173 164187 251239 164188
rect 252553 164187 252619 164190
rect 253422 164188 253428 164190
rect 253492 164188 253498 164252
rect 253933 164250 253999 164253
rect 254526 164250 254532 164252
rect 253933 164248 254532 164250
rect 253933 164192 253938 164248
rect 253994 164192 254532 164248
rect 253933 164190 254532 164192
rect 253933 164187 253999 164190
rect 254526 164188 254532 164190
rect 254596 164188 254602 164252
rect 255405 164250 255471 164253
rect 259453 164252 259519 164253
rect 255814 164250 255820 164252
rect 255405 164248 255820 164250
rect 255405 164192 255410 164248
rect 255466 164192 255820 164248
rect 255405 164190 255820 164192
rect 255405 164187 255471 164190
rect 255814 164188 255820 164190
rect 255884 164188 255890 164252
rect 259453 164250 259500 164252
rect 259408 164248 259500 164250
rect 259408 164192 259458 164248
rect 259408 164190 259500 164192
rect 259453 164188 259500 164190
rect 259564 164188 259570 164252
rect 262213 164250 262279 164253
rect 262806 164250 262812 164252
rect 262213 164248 262812 164250
rect 262213 164192 262218 164248
rect 262274 164192 262812 164248
rect 262213 164190 262812 164192
rect 259453 164187 259519 164188
rect 262213 164187 262279 164190
rect 262806 164188 262812 164190
rect 262876 164188 262882 164252
rect 263777 164250 263843 164253
rect 263910 164250 263916 164252
rect 263777 164248 263916 164250
rect 263777 164192 263782 164248
rect 263838 164192 263916 164248
rect 263777 164190 263916 164192
rect 263777 164187 263843 164190
rect 263910 164188 263916 164190
rect 263980 164188 263986 164252
rect 266302 164188 266308 164252
rect 266372 164250 266378 164252
rect 266445 164250 266511 164253
rect 266372 164248 266511 164250
rect 266372 164192 266450 164248
rect 266506 164192 266511 164248
rect 266372 164190 266511 164192
rect 266372 164188 266378 164190
rect 266445 164187 266511 164190
rect 267733 164250 267799 164253
rect 268694 164250 268700 164252
rect 267733 164248 268700 164250
rect 267733 164192 267738 164248
rect 267794 164192 268700 164248
rect 267733 164190 268700 164192
rect 267733 164187 267799 164190
rect 268694 164188 268700 164190
rect 268764 164188 268770 164252
rect 269113 164250 269179 164253
rect 269798 164250 269804 164252
rect 269113 164248 269804 164250
rect 269113 164192 269118 164248
rect 269174 164192 269804 164248
rect 269113 164190 269804 164192
rect 269113 164187 269179 164190
rect 269798 164188 269804 164190
rect 269868 164188 269874 164252
rect 270493 164250 270559 164253
rect 271270 164250 271276 164252
rect 270493 164248 271276 164250
rect 270493 164192 270498 164248
rect 270554 164192 271276 164248
rect 270493 164190 271276 164192
rect 270493 164187 270559 164190
rect 271270 164188 271276 164190
rect 271340 164188 271346 164252
rect 273294 164188 273300 164252
rect 273364 164250 273370 164252
rect 274541 164250 274607 164253
rect 273364 164248 274607 164250
rect 273364 164192 274546 164248
rect 274602 164192 274607 164248
rect 273364 164190 274607 164192
rect 273364 164188 273370 164190
rect 274541 164187 274607 164190
rect 276657 164250 276723 164253
rect 276974 164250 276980 164252
rect 276657 164248 276980 164250
rect 276657 164192 276662 164248
rect 276718 164192 276980 164248
rect 276657 164190 276980 164192
rect 276657 164187 276723 164190
rect 276974 164188 276980 164190
rect 277044 164188 277050 164252
rect 277393 164250 277459 164253
rect 396073 164252 396139 164253
rect 278078 164250 278084 164252
rect 277393 164248 278084 164250
rect 277393 164192 277398 164248
rect 277454 164192 278084 164248
rect 277393 164190 278084 164192
rect 277393 164187 277459 164190
rect 278078 164188 278084 164190
rect 278148 164188 278154 164252
rect 396022 164250 396028 164252
rect 395982 164190 396028 164250
rect 396092 164248 396139 164252
rect 396134 164192 396139 164248
rect 396022 164188 396028 164190
rect 396092 164188 396139 164192
rect 396073 164187 396139 164188
rect 398833 164250 398899 164253
rect 399518 164250 399524 164252
rect 398833 164248 399524 164250
rect 398833 164192 398838 164248
rect 398894 164192 399524 164248
rect 398833 164190 399524 164192
rect 398833 164187 398899 164190
rect 399518 164188 399524 164190
rect 399588 164188 399594 164252
rect 400213 164250 400279 164253
rect 403065 164252 403131 164253
rect 400438 164250 400444 164252
rect 400213 164248 400444 164250
rect 400213 164192 400218 164248
rect 400274 164192 400444 164248
rect 400213 164190 400444 164192
rect 400213 164187 400279 164190
rect 400438 164188 400444 164190
rect 400508 164188 400514 164252
rect 403014 164188 403020 164252
rect 403084 164250 403131 164252
rect 405733 164250 405799 164253
rect 406510 164250 406516 164252
rect 403084 164248 403176 164250
rect 403126 164192 403176 164248
rect 403084 164190 403176 164192
rect 405733 164248 406516 164250
rect 405733 164192 405738 164248
rect 405794 164192 406516 164248
rect 405733 164190 406516 164192
rect 403084 164188 403131 164190
rect 403065 164187 403131 164188
rect 405733 164187 405799 164190
rect 406510 164188 406516 164190
rect 406580 164188 406586 164252
rect 407113 164250 407179 164253
rect 407614 164250 407620 164252
rect 407113 164248 407620 164250
rect 407113 164192 407118 164248
rect 407174 164192 407620 164248
rect 407113 164190 407620 164192
rect 407113 164187 407179 164190
rect 407614 164188 407620 164190
rect 407684 164188 407690 164252
rect 408493 164250 408559 164253
rect 409965 164252 410031 164253
rect 411253 164252 411319 164253
rect 408718 164250 408724 164252
rect 408493 164248 408724 164250
rect 408493 164192 408498 164248
rect 408554 164192 408724 164248
rect 408493 164190 408724 164192
rect 408493 164187 408559 164190
rect 408718 164188 408724 164190
rect 408788 164188 408794 164252
rect 409965 164248 410012 164252
rect 410076 164250 410082 164252
rect 409965 164192 409970 164248
rect 409965 164188 410012 164192
rect 410076 164190 410122 164250
rect 411253 164248 411300 164252
rect 411364 164250 411370 164252
rect 412725 164250 412791 164253
rect 413502 164250 413508 164252
rect 411253 164192 411258 164248
rect 410076 164188 410082 164190
rect 411253 164188 411300 164192
rect 411364 164190 411410 164250
rect 412725 164248 413508 164250
rect 412725 164192 412730 164248
rect 412786 164192 413508 164248
rect 412725 164190 413508 164192
rect 411364 164188 411370 164190
rect 409965 164187 410031 164188
rect 411253 164187 411319 164188
rect 412725 164187 412791 164190
rect 413502 164188 413508 164190
rect 413572 164188 413578 164252
rect 414013 164250 414079 164253
rect 418245 164252 418311 164253
rect 414606 164250 414612 164252
rect 414013 164248 414612 164250
rect 414013 164192 414018 164248
rect 414074 164192 414612 164248
rect 414013 164190 414612 164192
rect 414013 164187 414079 164190
rect 414606 164188 414612 164190
rect 414676 164188 414682 164252
rect 418245 164250 418292 164252
rect 418200 164248 418292 164250
rect 418200 164192 418250 164248
rect 418200 164190 418292 164192
rect 418245 164188 418292 164190
rect 418356 164188 418362 164252
rect 419533 164250 419599 164253
rect 420678 164250 420684 164252
rect 419533 164248 420684 164250
rect 419533 164192 419538 164248
rect 419594 164192 420684 164248
rect 419533 164190 420684 164192
rect 418245 164187 418311 164188
rect 419533 164187 419599 164190
rect 420678 164188 420684 164190
rect 420748 164188 420754 164252
rect 420913 164250 420979 164253
rect 421782 164250 421788 164252
rect 420913 164248 421788 164250
rect 420913 164192 420918 164248
rect 420974 164192 421788 164248
rect 420913 164190 421788 164192
rect 420913 164187 420979 164190
rect 421782 164188 421788 164190
rect 421852 164188 421858 164252
rect 422886 164188 422892 164252
rect 422956 164250 422962 164252
rect 423581 164250 423647 164253
rect 422956 164248 423647 164250
rect 422956 164192 423586 164248
rect 423642 164192 423647 164248
rect 422956 164190 423647 164192
rect 422956 164188 422962 164190
rect 423581 164187 423647 164190
rect 425053 164250 425119 164253
rect 425278 164250 425284 164252
rect 425053 164248 425284 164250
rect 425053 164192 425058 164248
rect 425114 164192 425284 164248
rect 425053 164190 425284 164192
rect 425053 164187 425119 164190
rect 425278 164188 425284 164190
rect 425348 164188 425354 164252
rect 426382 164188 426388 164252
rect 426452 164250 426458 164252
rect 427721 164250 427787 164253
rect 426452 164248 427787 164250
rect 426452 164192 427726 164248
rect 427782 164192 427787 164248
rect 426452 164190 427787 164192
rect 426452 164188 426458 164190
rect 427721 164187 427787 164190
rect 428774 164188 428780 164252
rect 428844 164250 428850 164252
rect 429101 164250 429167 164253
rect 428844 164248 429167 164250
rect 428844 164192 429106 164248
rect 429162 164192 429167 164248
rect 428844 164190 429167 164192
rect 428844 164188 428850 164190
rect 429101 164187 429167 164190
rect 430573 164250 430639 164253
rect 430982 164250 430988 164252
rect 430573 164248 430988 164250
rect 430573 164192 430578 164248
rect 430634 164192 430988 164248
rect 430573 164190 430988 164192
rect 430573 164187 430639 164190
rect 430982 164188 430988 164190
rect 431052 164188 431058 164252
rect 431953 164250 432019 164253
rect 432270 164250 432276 164252
rect 431953 164248 432276 164250
rect 431953 164192 431958 164248
rect 432014 164192 432276 164248
rect 431953 164190 432276 164192
rect 431953 164187 432019 164190
rect 432270 164188 432276 164190
rect 432340 164188 432346 164252
rect 434805 164250 434871 164253
rect 435766 164250 435772 164252
rect 434805 164248 435772 164250
rect 434805 164192 434810 164248
rect 434866 164192 435772 164248
rect 434805 164190 435772 164192
rect 434805 164187 434871 164190
rect 435766 164188 435772 164190
rect 435836 164188 435842 164252
rect 436093 164250 436159 164253
rect 436870 164250 436876 164252
rect 436093 164248 436876 164250
rect 436093 164192 436098 164248
rect 436154 164192 436876 164248
rect 436093 164190 436876 164192
rect 436093 164187 436159 164190
rect 436870 164188 436876 164190
rect 436940 164188 436946 164252
rect 439262 164188 439268 164252
rect 439332 164250 439338 164252
rect 440141 164250 440207 164253
rect 439332 164248 440207 164250
rect 439332 164192 440146 164248
rect 440202 164192 440207 164248
rect 439332 164190 440207 164192
rect 439332 164188 439338 164190
rect 440141 164187 440207 164190
rect 203006 164052 203012 164116
rect 203076 164114 203082 164116
rect 325877 164114 325943 164117
rect 203076 164112 325943 164114
rect 203076 164056 325882 164112
rect 325938 164056 325943 164112
rect 203076 164054 325943 164056
rect 203076 164052 203082 164054
rect 325877 164051 325943 164054
rect 205030 163916 205036 163980
rect 205100 163978 205106 163980
rect 320950 163978 320956 163980
rect 205100 163918 320956 163978
rect 205100 163916 205106 163918
rect 320950 163916 320956 163918
rect 321020 163916 321026 163980
rect 217358 163508 217364 163572
rect 217428 163570 217434 163572
rect 218881 163570 218947 163573
rect 217428 163568 218947 163570
rect 217428 163512 218886 163568
rect 218942 163512 218947 163568
rect 217428 163510 218947 163512
rect 217428 163508 217434 163510
rect 218881 163507 218947 163510
rect 371049 163434 371115 163437
rect 377305 163434 377371 163437
rect 371049 163432 377371 163434
rect 371049 163376 371054 163432
rect 371110 163376 377310 163432
rect 377366 163376 377371 163432
rect 371049 163374 377371 163376
rect 371049 163371 371115 163374
rect 377305 163371 377371 163374
rect 57513 163298 57579 163301
rect 57830 163298 57836 163300
rect 57513 163296 57836 163298
rect 57513 163240 57518 163296
rect 57574 163240 57836 163296
rect 57513 163238 57836 163240
rect 57513 163235 57579 163238
rect 57830 163236 57836 163238
rect 57900 163236 57906 163300
rect 377305 163028 377371 163029
rect 377254 163026 377260 163028
rect -960 162740 480 162980
rect 377214 162966 377260 163026
rect 377324 163024 377371 163028
rect 377366 162968 377371 163024
rect 377254 162964 377260 162966
rect 377324 162964 377371 162968
rect 377305 162963 377371 162964
rect 216673 162754 216739 162757
rect 217542 162754 217548 162756
rect 216673 162752 217548 162754
rect 216673 162696 216678 162752
rect 216734 162696 217548 162752
rect 216673 162694 217548 162696
rect 216673 162691 216739 162694
rect 217542 162692 217548 162694
rect 217612 162754 217618 162756
rect 218881 162754 218947 162757
rect 217612 162752 218947 162754
rect 217612 162696 218886 162752
rect 218942 162696 218947 162752
rect 217612 162694 218947 162696
rect 217612 162692 217618 162694
rect 218881 162691 218947 162694
rect 217542 162556 217548 162620
rect 217612 162618 217618 162620
rect 218605 162618 218671 162621
rect 378041 162620 378107 162621
rect 217612 162616 218671 162618
rect 217612 162560 218610 162616
rect 218666 162560 218671 162616
rect 217612 162558 218671 162560
rect 217612 162556 217618 162558
rect 218605 162555 218671 162558
rect 377990 162556 377996 162620
rect 378060 162618 378107 162620
rect 378060 162616 378152 162618
rect 378102 162560 378152 162616
rect 378060 162558 378152 162560
rect 378060 162556 378107 162558
rect 378041 162555 378107 162556
rect 580257 152690 580323 152693
rect 583520 152690 584960 152780
rect 580257 152688 584960 152690
rect 580257 152632 580262 152688
rect 580318 152632 584960 152688
rect 580257 152630 584960 152632
rect 580257 152627 580323 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect -960 149774 674 149834
rect -960 149698 480 149774
rect 614 149698 674 149774
rect -960 149684 674 149698
rect 246 149638 674 149684
rect 246 149154 306 149638
rect 370630 149154 370636 149156
rect 246 149094 370636 149154
rect 370630 149092 370636 149094
rect 370700 149092 370706 149156
rect 276013 149018 276079 149021
rect 276657 149018 276723 149021
rect 357157 149018 357223 149021
rect 276013 149016 357223 149018
rect 276013 148960 276018 149016
rect 276074 148960 276662 149016
rect 276718 148960 357162 149016
rect 357218 148960 357223 149016
rect 276013 148958 357223 148960
rect 276013 148955 276079 148958
rect 276657 148955 276723 148958
rect 357157 148955 357223 148958
rect 217358 148276 217364 148340
rect 217428 148338 217434 148340
rect 276013 148338 276079 148341
rect 217428 148336 276079 148338
rect 217428 148280 276018 148336
rect 276074 148280 276079 148336
rect 217428 148278 276079 148280
rect 217428 148276 217434 148278
rect 276013 148275 276079 148278
rect 214189 146298 214255 146301
rect 214833 146298 214899 146301
rect 269113 146298 269179 146301
rect 214189 146296 269179 146298
rect 214189 146240 214194 146296
rect 214250 146240 214838 146296
rect 214894 146240 269118 146296
rect 269174 146240 269179 146296
rect 214189 146238 269179 146240
rect 214189 146235 214255 146238
rect 214833 146235 214899 146238
rect 269113 146235 269179 146238
rect 371785 146298 371851 146301
rect 376569 146298 376635 146301
rect 371785 146296 376635 146298
rect 371785 146240 371790 146296
rect 371846 146240 376574 146296
rect 376630 146240 376635 146296
rect 371785 146238 376635 146240
rect 371785 146235 371851 146238
rect 376569 146235 376635 146238
rect 379462 146236 379468 146300
rect 379532 146298 379538 146300
rect 380893 146298 380959 146301
rect 429193 146298 429259 146301
rect 379532 146296 429259 146298
rect 379532 146240 380898 146296
rect 380954 146240 429198 146296
rect 429254 146240 429259 146296
rect 379532 146238 429259 146240
rect 379532 146236 379538 146238
rect 380893 146235 380959 146238
rect 429193 146235 429259 146238
rect 211705 146162 211771 146165
rect 214833 146162 214899 146165
rect 211705 146160 214899 146162
rect 211705 146104 211710 146160
rect 211766 146104 214838 146160
rect 214894 146104 214899 146160
rect 211705 146102 214899 146104
rect 211705 146099 211771 146102
rect 214833 146099 214899 146102
rect 218421 146162 218487 146165
rect 266537 146162 266603 146165
rect 218421 146160 266603 146162
rect 218421 146104 218426 146160
rect 218482 146104 266542 146160
rect 266598 146104 266603 146160
rect 218421 146102 266603 146104
rect 218421 146099 218487 146102
rect 266537 146099 266603 146102
rect 395337 146162 395403 146165
rect 415393 146162 415459 146165
rect 395337 146160 415459 146162
rect 395337 146104 395342 146160
rect 395398 146104 415398 146160
rect 415454 146104 415459 146160
rect 395337 146102 415459 146104
rect 395337 146099 395403 146102
rect 415393 146099 415459 146102
rect 510613 146162 510679 146165
rect 510838 146162 510844 146164
rect 510613 146160 510844 146162
rect 510613 146104 510618 146160
rect 510674 146104 510844 146160
rect 510613 146102 510844 146104
rect 510613 146099 510679 146102
rect 510838 146100 510844 146102
rect 510908 146100 510914 146164
rect 58525 146026 58591 146029
rect 91093 146026 91159 146029
rect 58525 146024 91159 146026
rect 58525 145968 58530 146024
rect 58586 145968 91098 146024
rect 91154 145968 91159 146024
rect 58525 145966 91159 145968
rect 58525 145963 58591 145966
rect 91093 145963 91159 145966
rect 54845 145890 54911 145893
rect 57646 145890 57652 145892
rect 54845 145888 57652 145890
rect 54845 145832 54850 145888
rect 54906 145832 57652 145888
rect 54845 145830 57652 145832
rect 54845 145827 54911 145830
rect 57646 145828 57652 145830
rect 57716 145890 57722 145892
rect 96613 145890 96679 145893
rect 57716 145888 96679 145890
rect 57716 145832 96618 145888
rect 96674 145832 96679 145888
rect 57716 145830 96679 145832
rect 57716 145828 57722 145830
rect 96613 145827 96679 145830
rect 211797 145890 211863 145893
rect 237373 145890 237439 145893
rect 211797 145888 237439 145890
rect 211797 145832 211802 145888
rect 211858 145832 237378 145888
rect 237434 145832 237439 145888
rect 211797 145830 237439 145832
rect 211797 145827 211863 145830
rect 237373 145827 237439 145830
rect 372521 145890 372587 145893
rect 378409 145890 378475 145893
rect 423765 145890 423831 145893
rect 372521 145888 423831 145890
rect 372521 145832 372526 145888
rect 372582 145832 378414 145888
rect 378470 145832 423770 145888
rect 423826 145832 423831 145888
rect 372521 145830 423831 145832
rect 372521 145827 372587 145830
rect 378409 145827 378475 145830
rect 423765 145827 423831 145830
rect 56501 145754 56567 145757
rect 97257 145754 97323 145757
rect 56501 145752 97323 145754
rect 56501 145696 56506 145752
rect 56562 145696 97262 145752
rect 97318 145696 97323 145752
rect 56501 145694 97323 145696
rect 56501 145691 56567 145694
rect 97257 145691 97323 145694
rect 216397 145754 216463 145757
rect 270493 145754 270559 145757
rect 216397 145752 270559 145754
rect 216397 145696 216402 145752
rect 216458 145696 270498 145752
rect 270554 145696 270559 145752
rect 216397 145694 270559 145696
rect 216397 145691 216463 145694
rect 270493 145691 270559 145694
rect 376201 145754 376267 145757
rect 376569 145754 376635 145757
rect 423673 145754 423739 145757
rect 376201 145752 423739 145754
rect 376201 145696 376206 145752
rect 376262 145696 376574 145752
rect 376630 145696 423678 145752
rect 423734 145696 423739 145752
rect 376201 145694 423739 145696
rect 376201 145691 376267 145694
rect 376569 145691 376635 145694
rect 423673 145691 423739 145694
rect 52361 145618 52427 145621
rect 54569 145618 54635 145621
rect 99373 145618 99439 145621
rect 52361 145616 99439 145618
rect 52361 145560 52366 145616
rect 52422 145560 54574 145616
rect 54630 145560 99378 145616
rect 99434 145560 99439 145616
rect 52361 145558 99439 145560
rect 52361 145555 52427 145558
rect 54569 145555 54635 145558
rect 99373 145555 99439 145558
rect 214833 145618 214899 145621
rect 271873 145618 271939 145621
rect 214833 145616 271939 145618
rect 214833 145560 214838 145616
rect 214894 145560 271878 145616
rect 271934 145560 271939 145616
rect 214833 145558 271939 145560
rect 214833 145555 214899 145558
rect 271873 145555 271939 145558
rect 369025 145618 369091 145621
rect 379053 145618 379119 145621
rect 427813 145618 427879 145621
rect 369025 145616 427879 145618
rect 369025 145560 369030 145616
rect 369086 145560 379058 145616
rect 379114 145560 427818 145616
rect 427874 145560 427879 145616
rect 369025 145558 427879 145560
rect 369025 145555 369091 145558
rect 379053 145555 379119 145558
rect 427813 145555 427879 145558
rect 190862 145420 190868 145484
rect 190932 145482 190938 145484
rect 191741 145482 191807 145485
rect 190932 145480 191807 145482
rect 190932 145424 191746 145480
rect 191802 145424 191807 145480
rect 190932 145422 191807 145424
rect 190932 145420 190938 145422
rect 191741 145419 191807 145422
rect 178534 144876 178540 144940
rect 178604 144938 178610 144940
rect 179045 144938 179111 144941
rect 179689 144940 179755 144941
rect 179638 144938 179644 144940
rect 178604 144936 179111 144938
rect 178604 144880 179050 144936
rect 179106 144880 179111 144936
rect 178604 144878 179111 144880
rect 179598 144878 179644 144938
rect 179708 144936 179755 144940
rect 179750 144880 179755 144936
rect 178604 144876 178610 144878
rect 179045 144875 179111 144878
rect 179638 144876 179644 144878
rect 179708 144876 179755 144880
rect 217174 144876 217180 144940
rect 217244 144938 217250 144940
rect 218421 144938 218487 144941
rect 338481 144940 338547 144941
rect 338430 144938 338436 144940
rect 217244 144936 218487 144938
rect 217244 144880 218426 144936
rect 218482 144880 218487 144936
rect 217244 144878 218487 144880
rect 338390 144878 338436 144938
rect 338500 144936 338547 144940
rect 338542 144880 338547 144936
rect 217244 144876 217250 144878
rect 179689 144875 179755 144876
rect 218421 144875 218487 144878
rect 338430 144876 338436 144878
rect 338500 144876 338547 144880
rect 339718 144876 339724 144940
rect 339788 144938 339794 144940
rect 340229 144938 340295 144941
rect 339788 144936 340295 144938
rect 339788 144880 340234 144936
rect 340290 144880 340295 144936
rect 339788 144878 340295 144880
rect 339788 144876 339794 144878
rect 338481 144875 338547 144876
rect 340229 144875 340295 144878
rect 350942 144876 350948 144940
rect 351012 144938 351018 144940
rect 351637 144938 351703 144941
rect 351012 144936 351703 144938
rect 351012 144880 351642 144936
rect 351698 144880 351703 144936
rect 351012 144878 351703 144880
rect 351012 144876 351018 144878
rect 351637 144875 351703 144878
rect 498510 144876 498516 144940
rect 498580 144938 498586 144940
rect 498653 144938 498719 144941
rect 499849 144940 499915 144941
rect 499798 144938 499804 144940
rect 498580 144936 498719 144938
rect 498580 144880 498658 144936
rect 498714 144880 498719 144936
rect 498580 144878 498719 144880
rect 499758 144878 499804 144938
rect 499868 144936 499915 144940
rect 499910 144880 499915 144936
rect 498580 144876 498586 144878
rect 498653 144875 498719 144878
rect 499798 144876 499804 144878
rect 499868 144876 499915 144880
rect 499849 144875 499915 144876
rect 377806 144060 377812 144124
rect 377876 144122 377882 144124
rect 440233 144122 440299 144125
rect 377876 144120 440299 144122
rect 377876 144064 440238 144120
rect 440294 144064 440299 144120
rect 377876 144062 440299 144064
rect 377876 144060 377882 144062
rect 440233 144059 440299 144062
rect 57462 140796 57468 140860
rect 57532 140858 57538 140860
rect 59445 140858 59511 140861
rect 57532 140856 59511 140858
rect 57532 140800 59450 140856
rect 59506 140800 59511 140856
rect 57532 140798 59511 140800
rect 57532 140796 57538 140798
rect 59445 140795 59511 140798
rect 358997 139362 359063 139365
rect 519261 139362 519327 139365
rect 356562 139360 359063 139362
rect 356562 139304 359002 139360
rect 359058 139304 359063 139360
rect 356562 139302 359063 139304
rect 198825 139226 198891 139229
rect 197126 139224 198891 139226
rect 197126 139220 198830 139224
rect 196604 139168 198830 139220
rect 198886 139168 198891 139224
rect 356562 139190 356622 139302
rect 358997 139299 359063 139302
rect 516558 139360 519327 139362
rect 516558 139304 519266 139360
rect 519322 139304 519327 139360
rect 516558 139302 519327 139304
rect 516558 139190 516618 139302
rect 519261 139299 519327 139302
rect 583520 139212 584960 139452
rect 196604 139166 198891 139168
rect 196604 139160 197186 139166
rect 198825 139163 198891 139166
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 580441 112842 580507 112845
rect 583520 112842 584960 112932
rect 580441 112840 584960 112842
rect 580441 112784 580446 112840
rect 580502 112784 584960 112840
rect 580441 112782 584960 112784
rect 580441 112779 580507 112782
rect 583520 112692 584960 112782
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 57053 97474 57119 97477
rect 57053 97472 60062 97474
rect 57053 97416 57058 97472
rect 57114 97416 60062 97472
rect 57053 97414 60062 97416
rect 57053 97411 57119 97414
rect 60002 96894 60062 97414
rect 217501 96930 217567 96933
rect 376937 96930 377003 96933
rect 217501 96928 219450 96930
rect 217501 96872 217506 96928
rect 217562 96924 219450 96928
rect 376937 96928 379530 96930
rect 217562 96872 220064 96924
rect 217501 96870 220064 96872
rect 217501 96867 217567 96870
rect 219390 96864 220064 96870
rect 376937 96872 376942 96928
rect 376998 96924 379530 96928
rect 376998 96872 380052 96924
rect 376937 96870 380052 96872
rect 376937 96867 377003 96870
rect 379470 96864 380052 96870
rect 56685 96522 56751 96525
rect 56685 96520 60062 96522
rect 56685 96464 56690 96520
rect 56746 96464 60062 96520
rect 56685 96462 60062 96464
rect 56685 96459 56751 96462
rect 60002 95942 60062 96462
rect 216857 95978 216923 95981
rect 377857 95978 377923 95981
rect 216857 95976 219450 95978
rect 216857 95920 216862 95976
rect 216918 95972 219450 95976
rect 377857 95976 379530 95978
rect 216918 95920 220064 95972
rect 216857 95918 220064 95920
rect 216857 95915 216923 95918
rect 219390 95912 220064 95918
rect 377857 95920 377862 95976
rect 377918 95972 379530 95976
rect 377918 95920 380052 95972
rect 377857 95918 380052 95920
rect 377857 95915 377923 95918
rect 379470 95912 380052 95918
rect 57605 93802 57671 93805
rect 217593 93802 217659 93805
rect 377765 93802 377831 93805
rect 57605 93800 60062 93802
rect 57605 93744 57610 93800
rect 57666 93744 60062 93800
rect 57605 93742 60062 93744
rect 217593 93800 219450 93802
rect 217593 93744 217598 93800
rect 217654 93796 219450 93800
rect 377765 93800 379530 93802
rect 217654 93744 220064 93796
rect 217593 93742 220064 93744
rect 57605 93739 57671 93742
rect 217593 93739 217659 93742
rect 219390 93736 220064 93742
rect 377765 93744 377770 93800
rect 377826 93796 379530 93800
rect 377826 93744 380052 93796
rect 377765 93742 380052 93744
rect 377765 93739 377831 93742
rect 379470 93736 380052 93742
rect 57145 93394 57211 93397
rect 57145 93392 60062 93394
rect 57145 93336 57150 93392
rect 57206 93336 60062 93392
rect 57145 93334 60062 93336
rect 57145 93331 57211 93334
rect 60002 92814 60062 93334
rect 217409 92850 217475 92853
rect 376845 92850 376911 92853
rect 217409 92848 219450 92850
rect 217409 92792 217414 92848
rect 217470 92844 219450 92848
rect 376845 92848 379530 92850
rect 217470 92792 220064 92844
rect 217409 92790 220064 92792
rect 217409 92787 217475 92790
rect 219390 92784 220064 92790
rect 376845 92792 376850 92848
rect 376906 92844 379530 92848
rect 376906 92792 380052 92844
rect 376845 92790 380052 92792
rect 376845 92787 376911 92790
rect 379470 92784 380052 92790
rect 57697 91082 57763 91085
rect 217869 91082 217935 91085
rect 377489 91082 377555 91085
rect 57697 91080 60062 91082
rect 57697 91024 57702 91080
rect 57758 91024 60062 91080
rect 57697 91022 60062 91024
rect 217869 91080 219450 91082
rect 217869 91024 217874 91080
rect 217930 91076 219450 91080
rect 377489 91080 379530 91082
rect 217930 91024 220064 91076
rect 217869 91022 220064 91024
rect 57697 91019 57763 91022
rect 217869 91019 217935 91022
rect 219390 91016 220064 91022
rect 377489 91024 377494 91080
rect 377550 91076 379530 91080
rect 377550 91024 380052 91076
rect 377489 91022 380052 91024
rect 377489 91019 377555 91022
rect 379470 91016 380052 91022
rect 57421 90538 57487 90541
rect 57421 90536 60062 90538
rect 57421 90480 57426 90536
rect 57482 90480 60062 90536
rect 57421 90478 60062 90480
rect 57421 90475 57487 90478
rect 60002 89958 60062 90478
rect 217777 89994 217843 89997
rect 377673 89994 377739 89997
rect 217777 89992 219450 89994
rect 217777 89936 217782 89992
rect 217838 89988 219450 89992
rect 377673 89992 379530 89994
rect 217838 89936 220064 89988
rect 217777 89934 220064 89936
rect 217777 89931 217843 89934
rect 219390 89928 220064 89934
rect 377673 89936 377678 89992
rect 377734 89988 379530 89992
rect 377734 89936 380052 89988
rect 377673 89934 380052 89936
rect 377673 89931 377739 89934
rect 379470 89928 380052 89934
rect 57789 88226 57855 88229
rect 217685 88226 217751 88229
rect 377581 88226 377647 88229
rect 57789 88224 60062 88226
rect 57789 88168 57794 88224
rect 57850 88168 60062 88224
rect 57789 88166 60062 88168
rect 217685 88224 219450 88226
rect 217685 88168 217690 88224
rect 217746 88220 219450 88224
rect 377581 88224 379530 88226
rect 217746 88168 220064 88220
rect 217685 88166 220064 88168
rect 57789 88163 57855 88166
rect 217685 88163 217751 88166
rect 219390 88160 220064 88166
rect 377581 88168 377586 88224
rect 377642 88220 379530 88224
rect 377642 88168 380052 88220
rect 377581 88166 380052 88168
rect 377581 88163 377647 88166
rect 379470 88160 380052 88166
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 359457 79930 359523 79933
rect 518985 79930 519051 79933
rect 520181 79930 520247 79933
rect 356562 79928 359523 79930
rect 356562 79872 359462 79928
rect 359518 79872 359523 79928
rect 356562 79870 359523 79872
rect 199285 79386 199351 79389
rect 197126 79384 199351 79386
rect 197126 79380 199290 79384
rect 196604 79328 199290 79380
rect 199346 79328 199351 79384
rect 356562 79350 356622 79870
rect 359457 79867 359523 79870
rect 516558 79928 520247 79930
rect 516558 79872 518990 79928
rect 519046 79872 520186 79928
rect 520242 79872 520247 79928
rect 516558 79870 520247 79872
rect 516558 79350 516618 79870
rect 518985 79867 519051 79870
rect 520181 79867 520247 79870
rect 196604 79326 199351 79328
rect 196604 79320 197186 79326
rect 199285 79323 199351 79326
rect 359273 78298 359339 78301
rect 519353 78298 519419 78301
rect 356562 78296 359339 78298
rect 356562 78240 359278 78296
rect 359334 78240 359339 78296
rect 356562 78238 359339 78240
rect 199193 77754 199259 77757
rect 197126 77752 199259 77754
rect 197126 77748 199198 77752
rect 196604 77696 199198 77748
rect 199254 77696 199259 77752
rect 356562 77718 356622 78238
rect 359273 78235 359339 78238
rect 516558 78296 519419 78298
rect 516558 78240 519358 78296
rect 519414 78240 519419 78296
rect 516558 78238 519419 78240
rect 516558 77718 516618 78238
rect 519353 78235 519419 78238
rect 196604 77694 199259 77696
rect 196604 77688 197186 77694
rect 199193 77691 199259 77694
rect 359365 76938 359431 76941
rect 356562 76936 359431 76938
rect 356562 76880 359370 76936
rect 359426 76880 359431 76936
rect 356562 76878 359431 76880
rect 198733 76394 198799 76397
rect 197126 76392 198799 76394
rect 197126 76388 198738 76392
rect 196604 76336 198738 76388
rect 198794 76336 198799 76392
rect 356562 76358 356622 76878
rect 359365 76875 359431 76878
rect 519445 76802 519511 76805
rect 516558 76800 519511 76802
rect 516558 76744 519450 76800
rect 519506 76744 519511 76800
rect 516558 76742 519511 76744
rect 516558 76358 516618 76742
rect 519445 76739 519511 76742
rect 196604 76334 198799 76336
rect 196604 76328 197186 76334
rect 198733 76331 198799 76334
rect 359181 75442 359247 75445
rect 519077 75442 519143 75445
rect 356562 75440 359247 75442
rect 356562 75384 359186 75440
rect 359242 75384 359247 75440
rect 356562 75382 359247 75384
rect 198917 74898 198983 74901
rect 197126 74896 198983 74898
rect 197126 74892 198922 74896
rect 196604 74840 198922 74892
rect 198978 74840 198983 74896
rect 356562 74862 356622 75382
rect 359181 75379 359247 75382
rect 516558 75440 519143 75442
rect 516558 75384 519082 75440
rect 519138 75384 519143 75440
rect 516558 75382 519143 75384
rect 516558 74862 516618 75382
rect 519077 75379 519143 75382
rect 196604 74838 198983 74840
rect 196604 74832 197186 74838
rect 198917 74835 198983 74838
rect 519169 74218 519235 74221
rect 516558 74216 519235 74218
rect 516558 74160 519174 74216
rect 519230 74160 519235 74216
rect 516558 74158 519235 74160
rect 359089 74082 359155 74085
rect 356562 74080 359155 74082
rect 356562 74024 359094 74080
rect 359150 74024 359155 74080
rect 356562 74022 359155 74024
rect 199101 73674 199167 73677
rect 197126 73672 199167 73674
rect 197126 73668 199106 73672
rect 196604 73616 199106 73668
rect 199162 73616 199167 73672
rect 356562 73638 356622 74022
rect 359089 74019 359155 74022
rect 516558 73638 516618 74158
rect 519169 74155 519235 74158
rect 196604 73614 199167 73616
rect 196604 73608 197186 73614
rect 199101 73611 199167 73614
rect 580349 72994 580415 72997
rect 583520 72994 584960 73084
rect 580349 72992 584960 72994
rect 580349 72936 580354 72992
rect 580410 72936 584960 72992
rect 580349 72934 584960 72936
rect 580349 72931 580415 72934
rect 583520 72844 584960 72934
rect -960 71484 480 71724
rect 57513 70138 57579 70141
rect 57513 70136 60062 70138
rect 57513 70080 57518 70136
rect 57574 70080 60062 70136
rect 57513 70078 60062 70080
rect 57513 70075 57579 70078
rect 60002 69966 60062 70078
rect 207974 69940 207980 70004
rect 208044 70002 208050 70004
rect 376937 70002 377003 70005
rect 208044 69996 219450 70002
rect 376937 70000 379530 70002
rect 208044 69942 220064 69996
rect 208044 69940 208050 69942
rect 219390 69936 220064 69942
rect 376937 69944 376942 70000
rect 376998 69996 379530 70000
rect 376998 69944 380052 69996
rect 376937 69942 380052 69944
rect 376937 69939 377003 69942
rect 379470 69936 380052 69942
rect 57881 68914 57947 68917
rect 57881 68912 60062 68914
rect 57881 68856 57886 68912
rect 57942 68856 60062 68912
rect 57881 68854 60062 68856
rect 57881 68851 57947 68854
rect 60002 68334 60062 68854
rect 216673 68370 216739 68373
rect 376937 68370 377003 68373
rect 216673 68368 219450 68370
rect 216673 68312 216678 68368
rect 216734 68364 219450 68368
rect 376937 68368 379530 68370
rect 216734 68312 220064 68364
rect 216673 68310 220064 68312
rect 216673 68307 216739 68310
rect 219390 68304 220064 68310
rect 376937 68312 376942 68368
rect 376998 68364 379530 68368
rect 376998 68312 380052 68364
rect 376937 68310 380052 68312
rect 376937 68307 377003 68310
rect 379470 68304 380052 68310
rect 216765 68098 216831 68101
rect 376017 68098 376083 68101
rect 216765 68096 219450 68098
rect 46790 67764 46796 67828
rect 46860 67826 46866 67828
rect 60002 67826 60062 68062
rect 216765 68040 216770 68096
rect 216826 68092 219450 68096
rect 376017 68096 379530 68098
rect 216826 68040 220064 68092
rect 216765 68038 220064 68040
rect 216765 68035 216831 68038
rect 219390 68032 220064 68038
rect 376017 68040 376022 68096
rect 376078 68092 379530 68096
rect 376078 68040 380052 68092
rect 376017 68038 380052 68040
rect 376017 68035 376083 68038
rect 379470 68032 380052 68038
rect 46860 67766 60062 67826
rect 46860 67764 46866 67766
rect 378174 60556 378180 60620
rect 378244 60618 378250 60620
rect 378961 60618 379027 60621
rect 378244 60616 379027 60618
rect 378244 60560 378966 60616
rect 379022 60560 379027 60616
rect 378244 60558 379027 60560
rect 378244 60556 378250 60558
rect 378961 60555 379027 60558
rect 77109 59804 77175 59805
rect 83089 59804 83155 59805
rect 84193 59804 84259 59805
rect 99465 59804 99531 59805
rect 77109 59800 77142 59804
rect 77206 59802 77212 59804
rect 77109 59744 77114 59800
rect 77109 59740 77142 59744
rect 77206 59742 77266 59802
rect 83089 59800 83126 59804
rect 83190 59802 83196 59804
rect 83089 59744 83094 59800
rect 77206 59740 77212 59742
rect 83089 59740 83126 59744
rect 83190 59742 83246 59802
rect 84193 59800 84214 59804
rect 84278 59802 84284 59804
rect 99440 59802 99446 59804
rect 84193 59744 84198 59800
rect 83190 59740 83196 59742
rect 84193 59740 84214 59744
rect 84278 59742 84350 59802
rect 99374 59742 99446 59802
rect 99510 59800 99531 59804
rect 99526 59744 99531 59800
rect 84278 59740 84284 59742
rect 99440 59740 99446 59742
rect 99510 59740 99531 59744
rect 77109 59739 77175 59740
rect 83089 59739 83155 59740
rect 84193 59739 84259 59740
rect 99465 59739 99531 59740
rect 102777 59804 102843 59805
rect 107561 59804 107627 59805
rect 255865 59804 255931 59805
rect 260649 59804 260715 59805
rect 261753 59804 261819 59805
rect 262857 59804 262923 59805
rect 102777 59800 102846 59804
rect 102777 59744 102782 59800
rect 102838 59744 102846 59800
rect 102777 59740 102846 59744
rect 102910 59802 102916 59804
rect 102910 59742 102934 59802
rect 107561 59800 107606 59804
rect 107670 59802 107676 59804
rect 107561 59744 107566 59800
rect 102910 59740 102916 59742
rect 107561 59740 107606 59744
rect 107670 59742 107718 59802
rect 255865 59800 255910 59804
rect 255974 59802 255980 59804
rect 255865 59744 255870 59800
rect 107670 59740 107676 59742
rect 255865 59740 255910 59744
rect 255974 59742 256022 59802
rect 260649 59800 260670 59804
rect 260734 59802 260740 59804
rect 260649 59744 260654 59800
rect 255974 59740 255980 59742
rect 260649 59740 260670 59744
rect 260734 59742 260806 59802
rect 260734 59740 260740 59742
rect 261752 59740 261758 59804
rect 261822 59802 261828 59804
rect 262840 59802 262846 59804
rect 261822 59742 261910 59802
rect 262766 59742 262846 59802
rect 262910 59800 262923 59804
rect 262918 59744 262923 59800
rect 261822 59740 261828 59742
rect 262840 59740 262846 59742
rect 262910 59740 262923 59744
rect 102777 59739 102843 59740
rect 107561 59739 107627 59740
rect 255865 59739 255931 59740
rect 260649 59739 260715 59740
rect 261753 59739 261819 59740
rect 262857 59739 262923 59740
rect 263869 59804 263935 59805
rect 396073 59804 396139 59805
rect 263869 59800 263934 59804
rect 263869 59744 263874 59800
rect 263930 59744 263934 59800
rect 263869 59740 263934 59744
rect 263998 59802 264004 59804
rect 396048 59802 396054 59804
rect 263998 59742 264026 59802
rect 395982 59742 396054 59802
rect 396118 59800 396139 59804
rect 396134 59744 396139 59800
rect 263998 59740 264004 59742
rect 396048 59740 396054 59742
rect 396118 59740 396139 59744
rect 263869 59739 263935 59740
rect 396073 59739 396139 59740
rect 397085 59804 397151 59805
rect 403065 59804 403131 59805
rect 413553 59804 413619 59805
rect 415853 59804 415919 59805
rect 419441 59804 419507 59805
rect 397085 59800 397142 59804
rect 397206 59802 397212 59804
rect 397085 59744 397090 59800
rect 397085 59740 397142 59744
rect 397206 59742 397242 59802
rect 403065 59800 403126 59804
rect 403065 59744 403070 59800
rect 397206 59740 397212 59742
rect 403065 59740 403126 59744
rect 403190 59802 403196 59804
rect 403190 59742 403222 59802
rect 413553 59800 413598 59804
rect 413662 59802 413668 59804
rect 413553 59744 413558 59800
rect 403190 59740 403196 59742
rect 413553 59740 413598 59744
rect 413662 59742 413710 59802
rect 415853 59800 415910 59804
rect 415974 59802 415980 59804
rect 415853 59744 415858 59800
rect 413662 59740 413668 59742
rect 415853 59740 415910 59744
rect 415974 59742 416010 59802
rect 415974 59740 415980 59742
rect 419440 59740 419446 59804
rect 419510 59802 419516 59804
rect 419510 59742 419598 59802
rect 419510 59740 419516 59742
rect 397085 59739 397151 59740
rect 403065 59739 403131 59740
rect 413553 59739 413619 59740
rect 415853 59739 415919 59740
rect 419441 59739 419507 59740
rect 100753 59668 100819 59669
rect 100702 59666 100708 59668
rect 100662 59606 100708 59666
rect 100772 59664 100819 59668
rect 100814 59608 100819 59664
rect 100702 59604 100708 59606
rect 100772 59604 100819 59608
rect 100753 59603 100819 59604
rect 103881 59668 103947 59669
rect 114369 59668 114435 59669
rect 143533 59668 143599 59669
rect 103881 59664 103934 59668
rect 103998 59666 104004 59668
rect 103881 59608 103886 59664
rect 103881 59604 103934 59608
rect 103998 59606 104038 59666
rect 114369 59664 114406 59668
rect 114470 59666 114476 59668
rect 143504 59666 143510 59668
rect 114369 59608 114374 59664
rect 103998 59604 104004 59606
rect 114369 59604 114406 59608
rect 114470 59606 114526 59666
rect 143442 59606 143510 59666
rect 143574 59664 143599 59668
rect 143594 59608 143599 59664
rect 114470 59604 114476 59606
rect 143504 59604 143510 59606
rect 143574 59604 143599 59608
rect 103881 59603 103947 59604
rect 114369 59603 114435 59604
rect 143533 59603 143599 59604
rect 256969 59668 257035 59669
rect 308489 59668 308555 59669
rect 423489 59668 423555 59669
rect 503253 59668 503319 59669
rect 256969 59664 256998 59668
rect 257062 59666 257068 59668
rect 256969 59608 256974 59664
rect 256969 59604 256998 59608
rect 257062 59606 257126 59666
rect 257062 59604 257068 59606
rect 258488 59604 258494 59668
rect 258558 59604 258564 59668
rect 308489 59664 308542 59668
rect 308606 59666 308612 59668
rect 308489 59608 308494 59664
rect 308489 59604 308542 59608
rect 308606 59606 308646 59666
rect 423489 59664 423526 59668
rect 423590 59666 423596 59668
rect 503216 59666 503222 59668
rect 423489 59608 423494 59664
rect 308606 59604 308612 59606
rect 423489 59604 423526 59608
rect 423590 59606 423646 59666
rect 503162 59606 503222 59666
rect 503286 59664 503319 59668
rect 503314 59608 503319 59664
rect 423590 59604 423596 59606
rect 503216 59604 503222 59606
rect 503286 59604 503319 59608
rect 256969 59603 257035 59604
rect 219065 59532 219131 59533
rect 219014 59530 219020 59532
rect 218974 59470 219020 59530
rect 219084 59528 219131 59532
rect 219126 59472 219131 59528
rect 219014 59468 219020 59470
rect 219084 59468 219131 59472
rect 219065 59467 219131 59468
rect 85389 59396 85455 59397
rect 95877 59396 95943 59397
rect 98085 59396 98151 59397
rect 105261 59396 105327 59397
rect 106365 59396 106431 59397
rect 85389 59392 85436 59396
rect 85500 59394 85506 59396
rect 85389 59336 85394 59392
rect 85389 59332 85436 59336
rect 85500 59334 85546 59394
rect 95877 59392 95924 59396
rect 95988 59394 95994 59396
rect 95877 59336 95882 59392
rect 85500 59332 85506 59334
rect 95877 59332 95924 59336
rect 95988 59334 96034 59394
rect 98085 59392 98132 59396
rect 98196 59394 98202 59396
rect 98085 59336 98090 59392
rect 95988 59332 95994 59334
rect 98085 59332 98132 59336
rect 98196 59334 98242 59394
rect 105261 59392 105308 59396
rect 105372 59394 105378 59396
rect 105261 59336 105266 59392
rect 98196 59332 98202 59334
rect 105261 59332 105308 59336
rect 105372 59334 105418 59394
rect 106365 59392 106412 59396
rect 106476 59394 106482 59396
rect 106365 59336 106370 59392
rect 105372 59332 105378 59334
rect 106365 59332 106412 59336
rect 106476 59334 106522 59394
rect 106476 59332 106482 59334
rect 200614 59332 200620 59396
rect 200684 59394 200690 59396
rect 258496 59394 258556 59604
rect 308489 59603 308555 59604
rect 423489 59603 423555 59604
rect 503253 59603 503319 59604
rect 583520 59516 584960 59756
rect 200684 59334 258556 59394
rect 259453 59396 259519 59397
rect 398189 59396 398255 59397
rect 410701 59396 410767 59397
rect 416957 59396 417023 59397
rect 418153 59396 418219 59397
rect 259453 59392 259500 59396
rect 259564 59394 259570 59396
rect 259453 59336 259458 59392
rect 200684 59332 200690 59334
rect 259453 59332 259500 59336
rect 259564 59334 259610 59394
rect 398189 59392 398236 59396
rect 398300 59394 398306 59396
rect 398189 59336 398194 59392
rect 259564 59332 259570 59334
rect 398189 59332 398236 59336
rect 398300 59334 398346 59394
rect 410701 59392 410748 59396
rect 410812 59394 410818 59396
rect 410701 59336 410706 59392
rect 398300 59332 398306 59334
rect 410701 59332 410748 59336
rect 410812 59334 410858 59394
rect 416957 59392 417004 59396
rect 417068 59394 417074 59396
rect 418102 59394 418108 59396
rect 416957 59336 416962 59392
rect 410812 59332 410818 59334
rect 416957 59332 417004 59336
rect 417068 59334 417114 59394
rect 418062 59334 418108 59394
rect 418172 59392 418219 59396
rect 418214 59336 418219 59392
rect 417068 59332 417074 59334
rect 418102 59332 418108 59334
rect 418172 59332 418219 59336
rect 85389 59331 85455 59332
rect 95877 59331 95943 59332
rect 98085 59331 98151 59332
rect 105261 59331 105327 59332
rect 106365 59331 106431 59332
rect 259453 59331 259519 59332
rect 398189 59331 398255 59332
rect 410701 59331 410767 59332
rect 416957 59331 417023 59332
rect 418153 59331 418219 59332
rect 421005 59396 421071 59397
rect 421741 59396 421807 59397
rect 425237 59396 425303 59397
rect 425973 59396 426039 59397
rect 428181 59396 428247 59397
rect 468477 59396 468543 59397
rect 421005 59392 421052 59396
rect 421116 59394 421122 59396
rect 421005 59336 421010 59392
rect 421005 59332 421052 59336
rect 421116 59334 421162 59394
rect 421741 59392 421788 59396
rect 421852 59394 421858 59396
rect 421741 59336 421746 59392
rect 421116 59332 421122 59334
rect 421741 59332 421788 59336
rect 421852 59334 421898 59394
rect 425237 59392 425284 59396
rect 425348 59394 425354 59396
rect 425237 59336 425242 59392
rect 421852 59332 421858 59334
rect 425237 59332 425284 59336
rect 425348 59334 425394 59394
rect 425973 59392 426020 59396
rect 426084 59394 426090 59396
rect 425973 59336 425978 59392
rect 425348 59332 425354 59334
rect 425973 59332 426020 59336
rect 426084 59334 426130 59394
rect 428181 59392 428228 59396
rect 428292 59394 428298 59396
rect 428181 59336 428186 59392
rect 426084 59332 426090 59334
rect 428181 59332 428228 59336
rect 428292 59334 428338 59394
rect 468477 59392 468524 59396
rect 468588 59394 468594 59396
rect 468477 59336 468482 59392
rect 428292 59332 428298 59334
rect 468477 59332 468524 59336
rect 468588 59334 468634 59394
rect 468588 59332 468594 59334
rect 421005 59331 421071 59332
rect 421741 59331 421807 59332
rect 425237 59331 425303 59332
rect 425973 59331 426039 59332
rect 428181 59331 428247 59332
rect 468477 59331 468543 59332
rect 148501 59260 148567 59261
rect 150893 59260 150959 59261
rect 295885 59260 295951 59261
rect 298461 59260 298527 59261
rect 303429 59260 303495 59261
rect 54702 59196 54708 59260
rect 54772 59258 54778 59260
rect 140814 59258 140820 59260
rect 54772 59198 140820 59258
rect 54772 59196 54778 59198
rect 140814 59196 140820 59198
rect 140884 59196 140890 59260
rect 148501 59256 148548 59260
rect 148612 59258 148618 59260
rect 148501 59200 148506 59256
rect 148501 59196 148548 59200
rect 148612 59198 148658 59258
rect 150893 59256 150940 59260
rect 151004 59258 151010 59260
rect 150893 59200 150898 59256
rect 148612 59196 148618 59198
rect 150893 59196 150940 59200
rect 151004 59198 151050 59258
rect 151004 59196 151010 59198
rect 205214 59196 205220 59260
rect 205284 59258 205290 59260
rect 290958 59258 290964 59260
rect 205284 59198 290964 59258
rect 205284 59196 205290 59198
rect 290958 59196 290964 59198
rect 291028 59196 291034 59260
rect 295885 59256 295932 59260
rect 295996 59258 296002 59260
rect 295885 59200 295890 59256
rect 295885 59196 295932 59200
rect 295996 59198 296042 59258
rect 298461 59256 298508 59260
rect 298572 59258 298578 59260
rect 298461 59200 298466 59256
rect 295996 59196 296002 59198
rect 298461 59196 298508 59200
rect 298572 59198 298618 59258
rect 303429 59256 303476 59260
rect 303540 59258 303546 59260
rect 303429 59200 303434 59256
rect 298572 59196 298578 59198
rect 303429 59196 303476 59200
rect 303540 59198 303586 59258
rect 303540 59196 303546 59198
rect 357934 59196 357940 59260
rect 358004 59258 358010 59260
rect 478454 59258 478460 59260
rect 358004 59198 478460 59258
rect 358004 59196 358010 59198
rect 478454 59196 478460 59198
rect 478524 59196 478530 59260
rect 148501 59195 148567 59196
rect 150893 59195 150959 59196
rect 295885 59195 295951 59196
rect 298461 59195 298527 59196
rect 303429 59195 303495 59196
rect 138381 59124 138447 59125
rect 53414 59060 53420 59124
rect 53484 59122 53490 59124
rect 135846 59122 135852 59124
rect 53484 59062 135852 59122
rect 53484 59060 53490 59062
rect 135846 59060 135852 59062
rect 135916 59060 135922 59124
rect 138381 59120 138428 59124
rect 138492 59122 138498 59124
rect 138381 59064 138386 59120
rect 138381 59060 138428 59064
rect 138492 59062 138538 59122
rect 138492 59060 138498 59062
rect 206686 59060 206692 59124
rect 206756 59122 206762 59124
rect 283414 59122 283420 59124
rect 206756 59062 283420 59122
rect 206756 59060 206762 59062
rect 283414 59060 283420 59062
rect 283484 59060 283490 59124
rect 371918 59060 371924 59124
rect 371988 59122 371994 59124
rect 485998 59122 486004 59124
rect 371988 59062 486004 59122
rect 371988 59060 371994 59062
rect 485998 59060 486004 59062
rect 486068 59060 486074 59124
rect 138381 59059 138447 59060
rect 59118 58924 59124 58988
rect 59188 58986 59194 58988
rect 125910 58986 125916 58988
rect 59188 58926 125916 58986
rect 59188 58924 59194 58926
rect 125910 58924 125916 58926
rect 125980 58924 125986 58988
rect 201350 58924 201356 58988
rect 201420 58986 201426 58988
rect 278446 58986 278452 58988
rect 201420 58926 278452 58986
rect 201420 58924 201426 58926
rect 278446 58924 278452 58926
rect 278516 58924 278522 58988
rect 374494 58924 374500 58988
rect 374564 58986 374570 58988
rect 473486 58986 473492 58988
rect 374564 58926 473492 58986
rect 374564 58924 374570 58926
rect 473486 58924 473492 58926
rect 473556 58924 473562 58988
rect 48078 58788 48084 58852
rect 48148 58850 48154 58852
rect 111006 58850 111012 58852
rect 48148 58790 111012 58850
rect 48148 58788 48154 58790
rect 111006 58788 111012 58790
rect 111076 58788 111082 58852
rect 202638 58788 202644 58852
rect 202708 58850 202714 58852
rect 276054 58850 276060 58852
rect 202708 58790 276060 58850
rect 202708 58788 202714 58790
rect 276054 58788 276060 58790
rect 276124 58788 276130 58852
rect 367870 58788 367876 58852
rect 367940 58850 367946 58852
rect 458398 58850 458404 58852
rect 367940 58790 458404 58850
rect 367940 58788 367946 58790
rect 458398 58788 458404 58790
rect 458468 58788 458474 58852
rect -960 58578 480 58668
rect 46606 58652 46612 58716
rect 46676 58714 46682 58716
rect 108246 58714 108252 58716
rect 46676 58654 108252 58714
rect 46676 58652 46682 58654
rect 108246 58652 108252 58654
rect 108316 58652 108322 58716
rect 202086 58652 202092 58716
rect 202156 58714 202162 58716
rect 250662 58714 250668 58716
rect 202156 58654 250668 58714
rect 202156 58652 202162 58654
rect 250662 58652 250668 58654
rect 250732 58652 250738 58716
rect 375966 58652 375972 58716
rect 376036 58714 376042 58716
rect 463550 58714 463556 58716
rect 376036 58654 463556 58714
rect 376036 58652 376042 58654
rect 463550 58652 463556 58654
rect 463620 58652 463626 58716
rect 3509 58578 3575 58581
rect -960 58576 3575 58578
rect -960 58520 3514 58576
rect 3570 58520 3575 58576
rect -960 58518 3575 58520
rect -960 58428 480 58518
rect 3509 58515 3575 58518
rect 59854 58516 59860 58580
rect 59924 58578 59930 58580
rect 115974 58578 115980 58580
rect 59924 58518 115980 58578
rect 59924 58516 59930 58518
rect 115974 58516 115980 58518
rect 116044 58516 116050 58580
rect 219198 58516 219204 58580
rect 219268 58578 219274 58580
rect 219341 58578 219407 58581
rect 219268 58576 219407 58578
rect 219268 58520 219346 58576
rect 219402 58520 219407 58576
rect 219268 58518 219407 58520
rect 219268 58516 219274 58518
rect 219341 58515 219407 58518
rect 222929 58578 222995 58581
rect 265198 58578 265204 58580
rect 222929 58576 265204 58578
rect 222929 58520 222934 58576
rect 222990 58520 265204 58576
rect 222929 58518 265204 58520
rect 222929 58515 222995 58518
rect 265198 58516 265204 58518
rect 265268 58516 265274 58580
rect 367686 58516 367692 58580
rect 367756 58578 367762 58580
rect 453430 58578 453436 58580
rect 367756 58518 453436 58578
rect 367756 58516 367762 58518
rect 453430 58516 453436 58518
rect 453500 58516 453506 58580
rect 59302 58380 59308 58444
rect 59372 58442 59378 58444
rect 101070 58442 101076 58444
rect 59372 58382 101076 58442
rect 59372 58380 59378 58382
rect 101070 58380 101076 58382
rect 101140 58380 101146 58444
rect 217542 58380 217548 58444
rect 217612 58442 217618 58444
rect 257838 58442 257844 58444
rect 217612 58382 257844 58442
rect 217612 58380 217618 58382
rect 257838 58380 257844 58382
rect 257908 58380 257914 58444
rect 377990 58380 377996 58444
rect 378060 58442 378066 58444
rect 420678 58442 420684 58444
rect 378060 58382 420684 58442
rect 378060 58380 378066 58382
rect 420678 58380 420684 58382
rect 420748 58380 420754 58444
rect 217174 58244 217180 58308
rect 217244 58306 217250 58308
rect 222929 58306 222995 58309
rect 217244 58304 222995 58306
rect 217244 58248 222934 58304
rect 222990 58248 222995 58304
rect 217244 58246 222995 58248
rect 217244 58244 217250 58246
rect 222929 58243 222995 58246
rect 92238 58108 92244 58172
rect 92308 58108 92314 58172
rect 113582 58108 113588 58172
rect 113652 58108 113658 58172
rect 128302 58108 128308 58172
rect 128372 58108 128378 58172
rect 153326 58108 153332 58172
rect 153396 58108 153402 58172
rect 236126 58108 236132 58172
rect 236196 58108 236202 58172
rect 272190 58108 272196 58172
rect 272260 58108 272266 58172
rect 275686 58108 275692 58172
rect 275756 58108 275762 58172
rect 300894 58108 300900 58172
rect 300964 58108 300970 58172
rect 315798 58108 315804 58172
rect 315868 58108 315874 58172
rect 325918 58108 325924 58172
rect 325988 58108 325994 58172
rect 401726 58108 401732 58172
rect 401796 58108 401802 58172
rect 455822 58108 455828 58172
rect 455892 58108 455898 58172
rect 92246 57901 92306 58108
rect 113590 57901 113650 58108
rect 76005 57900 76071 57901
rect 78213 57900 78279 57901
rect 76005 57896 76052 57900
rect 76116 57898 76122 57900
rect 76005 57840 76010 57896
rect 76005 57836 76052 57840
rect 76116 57838 76162 57898
rect 78213 57896 78260 57900
rect 78324 57898 78330 57900
rect 78673 57898 78739 57901
rect 80421 57900 80487 57901
rect 79542 57898 79548 57900
rect 78213 57840 78218 57896
rect 76116 57836 76122 57838
rect 78213 57836 78260 57840
rect 78324 57838 78370 57898
rect 78673 57896 79548 57898
rect 78673 57840 78678 57896
rect 78734 57840 79548 57896
rect 78673 57838 79548 57840
rect 78324 57836 78330 57838
rect 76005 57835 76071 57836
rect 78213 57835 78279 57836
rect 78673 57835 78739 57838
rect 79542 57836 79548 57838
rect 79612 57836 79618 57900
rect 80421 57896 80468 57900
rect 80532 57898 80538 57900
rect 81433 57898 81499 57901
rect 86493 57900 86559 57901
rect 81934 57898 81940 57900
rect 80421 57840 80426 57896
rect 80421 57836 80468 57840
rect 80532 57838 80578 57898
rect 81433 57896 81940 57898
rect 81433 57840 81438 57896
rect 81494 57840 81940 57896
rect 81433 57838 81940 57840
rect 80532 57836 80538 57838
rect 80421 57835 80487 57836
rect 81433 57835 81499 57838
rect 81934 57836 81940 57838
rect 82004 57836 82010 57900
rect 86493 57896 86540 57900
rect 86604 57898 86610 57900
rect 86953 57898 87019 57901
rect 87638 57898 87644 57900
rect 86493 57840 86498 57896
rect 86493 57836 86540 57840
rect 86604 57838 86650 57898
rect 86953 57896 87644 57898
rect 86953 57840 86958 57896
rect 87014 57840 87644 57896
rect 86953 57838 87644 57840
rect 86604 57836 86610 57838
rect 86493 57835 86559 57836
rect 86953 57835 87019 57838
rect 87638 57836 87644 57838
rect 87708 57836 87714 57900
rect 88333 57898 88399 57901
rect 89989 57900 90055 57901
rect 90725 57900 90791 57901
rect 88742 57898 88748 57900
rect 88333 57896 88748 57898
rect 88333 57840 88338 57896
rect 88394 57840 88748 57896
rect 88333 57838 88748 57840
rect 88333 57835 88399 57838
rect 88742 57836 88748 57838
rect 88812 57836 88818 57900
rect 89989 57896 90036 57900
rect 90100 57898 90106 57900
rect 89989 57840 89994 57896
rect 89989 57836 90036 57840
rect 90100 57838 90146 57898
rect 90725 57896 90772 57900
rect 90836 57898 90842 57900
rect 91185 57898 91251 57901
rect 91318 57898 91324 57900
rect 90725 57840 90730 57896
rect 90100 57836 90106 57838
rect 90725 57836 90772 57840
rect 90836 57838 90882 57898
rect 91185 57896 91324 57898
rect 91185 57840 91190 57896
rect 91246 57840 91324 57896
rect 91185 57838 91324 57840
rect 90836 57836 90842 57838
rect 89989 57835 90055 57836
rect 90725 57835 90791 57836
rect 91185 57835 91251 57838
rect 91318 57836 91324 57838
rect 91388 57836 91394 57900
rect 92197 57896 92306 57901
rect 92197 57840 92202 57896
rect 92258 57840 92306 57896
rect 92197 57838 92306 57840
rect 92473 57898 92539 57901
rect 93669 57900 93735 57901
rect 94405 57900 94471 57901
rect 98453 57900 98519 57901
rect 101765 57900 101831 57901
rect 108573 57900 108639 57901
rect 109493 57900 109559 57901
rect 111149 57900 111215 57901
rect 93342 57898 93348 57900
rect 92473 57896 93348 57898
rect 92473 57840 92478 57896
rect 92534 57840 93348 57896
rect 92473 57838 93348 57840
rect 92197 57835 92263 57838
rect 92473 57835 92539 57838
rect 93342 57836 93348 57838
rect 93412 57836 93418 57900
rect 93669 57896 93716 57900
rect 93780 57898 93786 57900
rect 93669 57840 93674 57896
rect 93669 57836 93716 57840
rect 93780 57838 93826 57898
rect 94405 57896 94452 57900
rect 94516 57898 94522 57900
rect 94405 57840 94410 57896
rect 93780 57836 93786 57838
rect 94405 57836 94452 57840
rect 94516 57838 94562 57898
rect 98453 57896 98500 57900
rect 98564 57898 98570 57900
rect 98453 57840 98458 57896
rect 94516 57836 94522 57838
rect 98453 57836 98500 57840
rect 98564 57838 98610 57898
rect 101765 57896 101812 57900
rect 101876 57898 101882 57900
rect 101765 57840 101770 57896
rect 98564 57836 98570 57838
rect 101765 57836 101812 57840
rect 101876 57838 101922 57898
rect 108573 57896 108620 57900
rect 108684 57898 108690 57900
rect 108573 57840 108578 57896
rect 101876 57836 101882 57838
rect 108573 57836 108620 57840
rect 108684 57838 108730 57898
rect 109493 57896 109540 57900
rect 109604 57898 109610 57900
rect 109493 57840 109498 57896
rect 108684 57836 108690 57838
rect 109493 57836 109540 57840
rect 109604 57838 109650 57898
rect 111149 57896 111196 57900
rect 111260 57898 111266 57900
rect 111149 57840 111154 57896
rect 109604 57836 109610 57838
rect 111149 57836 111196 57840
rect 111260 57838 111306 57898
rect 113541 57896 113650 57901
rect 113541 57840 113546 57896
rect 113602 57840 113650 57896
rect 113541 57838 113650 57840
rect 116485 57898 116551 57901
rect 117957 57900 118023 57901
rect 120717 57900 120783 57901
rect 123477 57900 123543 57901
rect 116894 57898 116900 57900
rect 116485 57896 116900 57898
rect 116485 57840 116490 57896
rect 116546 57840 116900 57896
rect 116485 57838 116900 57840
rect 111260 57836 111266 57838
rect 93669 57835 93735 57836
rect 94405 57835 94471 57836
rect 98453 57835 98519 57836
rect 101765 57835 101831 57836
rect 108573 57835 108639 57836
rect 109493 57835 109559 57836
rect 111149 57835 111215 57836
rect 113541 57835 113607 57838
rect 116485 57835 116551 57838
rect 116894 57836 116900 57838
rect 116964 57836 116970 57900
rect 117957 57896 118004 57900
rect 118068 57898 118074 57900
rect 117957 57840 117962 57896
rect 117957 57836 118004 57840
rect 118068 57838 118114 57898
rect 120717 57896 120764 57900
rect 120828 57898 120834 57900
rect 120717 57840 120722 57896
rect 118068 57836 118074 57838
rect 120717 57836 120764 57840
rect 120828 57838 120874 57898
rect 123477 57896 123524 57900
rect 123588 57898 123594 57900
rect 123477 57840 123482 57896
rect 120828 57836 120834 57838
rect 123477 57836 123524 57840
rect 123588 57838 123634 57898
rect 123588 57836 123594 57838
rect 117957 57835 118023 57836
rect 120717 57835 120783 57836
rect 123477 57835 123543 57836
rect 55070 57700 55076 57764
rect 55140 57762 55146 57764
rect 128310 57762 128370 58108
rect 153334 57901 153394 58108
rect 236134 57901 236194 58108
rect 130837 57900 130903 57901
rect 145557 57900 145623 57901
rect 130837 57896 130884 57900
rect 130948 57898 130954 57900
rect 130837 57840 130842 57896
rect 130837 57836 130884 57840
rect 130948 57838 130994 57898
rect 145557 57896 145604 57900
rect 145668 57898 145674 57900
rect 145557 57840 145562 57896
rect 130948 57836 130954 57838
rect 145557 57836 145604 57840
rect 145668 57838 145714 57898
rect 153285 57896 153394 57901
rect 153285 57840 153290 57896
rect 153346 57840 153394 57896
rect 153285 57838 153394 57840
rect 183461 57900 183527 57901
rect 183461 57896 183508 57900
rect 183572 57898 183578 57900
rect 183461 57840 183466 57896
rect 145668 57836 145674 57838
rect 130837 57835 130903 57836
rect 145557 57835 145623 57836
rect 153285 57835 153351 57838
rect 183461 57836 183508 57840
rect 183572 57838 183618 57898
rect 236085 57896 236194 57901
rect 236085 57840 236090 57896
rect 236146 57840 236194 57896
rect 236085 57838 236194 57840
rect 238109 57900 238175 57901
rect 238109 57896 238156 57900
rect 238220 57898 238226 57900
rect 238753 57898 238819 57901
rect 240501 57900 240567 57901
rect 239254 57898 239260 57900
rect 238109 57840 238114 57896
rect 183572 57836 183578 57838
rect 183461 57835 183527 57836
rect 236085 57835 236151 57838
rect 238109 57836 238156 57840
rect 238220 57838 238266 57898
rect 238753 57896 239260 57898
rect 238753 57840 238758 57896
rect 238814 57840 239260 57896
rect 238753 57838 239260 57840
rect 238220 57836 238226 57838
rect 238109 57835 238175 57836
rect 238753 57835 238819 57838
rect 239254 57836 239260 57838
rect 239324 57836 239330 57900
rect 240501 57896 240548 57900
rect 240612 57898 240618 57900
rect 241513 57898 241579 57901
rect 242893 57900 242959 57901
rect 241646 57898 241652 57900
rect 240501 57840 240506 57896
rect 240501 57836 240548 57840
rect 240612 57838 240658 57898
rect 241513 57896 241652 57898
rect 241513 57840 241518 57896
rect 241574 57840 241652 57896
rect 241513 57838 241652 57840
rect 240612 57836 240618 57838
rect 240501 57835 240567 57836
rect 241513 57835 241579 57838
rect 241646 57836 241652 57838
rect 241716 57836 241722 57900
rect 242893 57896 242940 57900
rect 243004 57898 243010 57900
rect 242893 57840 242898 57896
rect 242893 57836 242940 57840
rect 243004 57838 243050 57898
rect 243004 57836 243010 57838
rect 244222 57836 244228 57900
rect 244292 57898 244298 57900
rect 244365 57898 244431 57901
rect 244292 57896 244431 57898
rect 244292 57840 244370 57896
rect 244426 57840 244431 57896
rect 244292 57838 244431 57840
rect 244292 57836 244298 57838
rect 242893 57835 242959 57836
rect 244365 57835 244431 57838
rect 245285 57900 245351 57901
rect 245285 57896 245332 57900
rect 245396 57898 245402 57900
rect 245653 57898 245719 57901
rect 247677 57900 247743 57901
rect 246430 57898 246436 57900
rect 245285 57840 245290 57896
rect 245285 57836 245332 57840
rect 245396 57838 245442 57898
rect 245653 57896 246436 57898
rect 245653 57840 245658 57896
rect 245714 57840 246436 57896
rect 245653 57838 246436 57840
rect 245396 57836 245402 57838
rect 245285 57835 245351 57836
rect 245653 57835 245719 57838
rect 246430 57836 246436 57838
rect 246500 57836 246506 57900
rect 247677 57896 247724 57900
rect 247788 57898 247794 57900
rect 248137 57898 248203 57901
rect 248270 57898 248276 57900
rect 247677 57840 247682 57896
rect 247677 57836 247724 57840
rect 247788 57838 247834 57898
rect 248137 57896 248276 57898
rect 248137 57840 248142 57896
rect 248198 57840 248276 57896
rect 248137 57838 248276 57840
rect 247788 57836 247794 57838
rect 247677 57835 247743 57836
rect 248137 57835 248203 57838
rect 248270 57836 248276 57838
rect 248340 57836 248346 57900
rect 248413 57898 248479 57901
rect 248638 57898 248644 57900
rect 248413 57896 248644 57898
rect 248413 57840 248418 57896
rect 248474 57840 248644 57896
rect 248413 57838 248644 57840
rect 248413 57835 248479 57838
rect 248638 57836 248644 57838
rect 248708 57836 248714 57900
rect 249793 57898 249859 57901
rect 251173 57900 251239 57901
rect 250110 57898 250116 57900
rect 249793 57896 250116 57898
rect 249793 57840 249798 57896
rect 249854 57840 250116 57896
rect 249793 57838 250116 57840
rect 249793 57835 249859 57838
rect 250110 57836 250116 57838
rect 250180 57836 250186 57900
rect 251173 57898 251220 57900
rect 251128 57896 251220 57898
rect 251128 57840 251178 57896
rect 251128 57838 251220 57840
rect 251173 57836 251220 57838
rect 251284 57836 251290 57900
rect 251357 57898 251423 57901
rect 253381 57900 253447 57901
rect 252318 57898 252324 57900
rect 251357 57896 252324 57898
rect 251357 57840 251362 57896
rect 251418 57840 252324 57896
rect 251357 57838 252324 57840
rect 251173 57835 251239 57836
rect 251357 57835 251423 57838
rect 252318 57836 252324 57838
rect 252388 57836 252394 57900
rect 253381 57896 253428 57900
rect 253492 57898 253498 57900
rect 253933 57898 253999 57901
rect 271229 57900 271295 57901
rect 254526 57898 254532 57900
rect 253381 57840 253386 57896
rect 253381 57836 253428 57840
rect 253492 57838 253538 57898
rect 253933 57896 254532 57898
rect 253933 57840 253938 57896
rect 253994 57840 254532 57896
rect 253933 57838 254532 57840
rect 253492 57836 253498 57838
rect 253381 57835 253447 57836
rect 253933 57835 253999 57838
rect 254526 57836 254532 57838
rect 254596 57836 254602 57900
rect 270902 57898 270908 57900
rect 258030 57838 270908 57898
rect 183185 57764 183251 57765
rect 183134 57762 183140 57764
rect 55140 57702 128370 57762
rect 183094 57702 183140 57762
rect 183204 57760 183251 57764
rect 183246 57704 183251 57760
rect 55140 57700 55146 57702
rect 183134 57700 183140 57702
rect 183204 57700 183251 57704
rect 206134 57700 206140 57764
rect 206204 57762 206210 57764
rect 258030 57762 258090 57838
rect 270902 57836 270908 57838
rect 270972 57836 270978 57900
rect 271229 57896 271276 57900
rect 271340 57898 271346 57900
rect 271873 57898 271939 57901
rect 272198 57898 272258 58108
rect 275694 57901 275754 58108
rect 300902 57901 300962 58108
rect 271229 57840 271234 57896
rect 271229 57836 271276 57840
rect 271340 57838 271386 57898
rect 271873 57896 272258 57898
rect 271873 57840 271878 57896
rect 271934 57840 272258 57896
rect 271873 57838 272258 57840
rect 273253 57900 273319 57901
rect 273253 57896 273300 57900
rect 273364 57898 273370 57900
rect 273253 57840 273258 57896
rect 271340 57836 271346 57838
rect 271229 57835 271295 57836
rect 271873 57835 271939 57838
rect 273253 57836 273300 57840
rect 273364 57838 273410 57898
rect 275645 57896 275754 57901
rect 275645 57840 275650 57896
rect 275706 57840 275754 57896
rect 275645 57838 275754 57840
rect 278037 57900 278103 57901
rect 279049 57900 279115 57901
rect 278037 57896 278084 57900
rect 278148 57898 278154 57900
rect 278998 57898 279004 57900
rect 278037 57840 278042 57896
rect 273364 57836 273370 57838
rect 273253 57835 273319 57836
rect 275645 57835 275711 57838
rect 278037 57836 278084 57840
rect 278148 57838 278194 57898
rect 278958 57838 279004 57898
rect 279068 57896 279115 57900
rect 279110 57840 279115 57896
rect 278148 57836 278154 57838
rect 278998 57836 279004 57838
rect 279068 57836 279115 57840
rect 278037 57835 278103 57836
rect 279049 57835 279115 57836
rect 287605 57898 287671 57901
rect 293309 57900 293375 57901
rect 288198 57898 288204 57900
rect 287605 57896 288204 57898
rect 287605 57840 287610 57896
rect 287666 57840 288204 57896
rect 287605 57838 288204 57840
rect 287605 57835 287671 57838
rect 288198 57836 288204 57838
rect 288268 57836 288274 57900
rect 293309 57896 293356 57900
rect 293420 57898 293426 57900
rect 293309 57840 293314 57896
rect 293309 57836 293356 57840
rect 293420 57838 293466 57898
rect 300853 57896 300962 57901
rect 300853 57840 300858 57896
rect 300914 57840 300962 57896
rect 300853 57838 300962 57840
rect 305821 57900 305887 57901
rect 310973 57900 311039 57901
rect 313365 57900 313431 57901
rect 305821 57896 305868 57900
rect 305932 57898 305938 57900
rect 305821 57840 305826 57896
rect 293420 57836 293426 57838
rect 293309 57835 293375 57836
rect 300853 57835 300919 57838
rect 305821 57836 305868 57840
rect 305932 57838 305978 57898
rect 310973 57896 311020 57900
rect 311084 57898 311090 57900
rect 310973 57840 310978 57896
rect 305932 57836 305938 57838
rect 310973 57836 311020 57840
rect 311084 57838 311130 57898
rect 313365 57896 313412 57900
rect 313476 57898 313482 57900
rect 315021 57898 315087 57901
rect 315806 57898 315866 58108
rect 325926 57901 325986 58108
rect 313365 57840 313370 57896
rect 311084 57836 311090 57838
rect 313365 57836 313412 57840
rect 313476 57838 313522 57898
rect 315021 57896 315866 57898
rect 315021 57840 315026 57896
rect 315082 57840 315866 57896
rect 315021 57838 315866 57840
rect 318241 57898 318307 57901
rect 318374 57898 318380 57900
rect 318241 57896 318380 57898
rect 318241 57840 318246 57896
rect 318302 57840 318380 57896
rect 318241 57838 318380 57840
rect 313476 57836 313482 57838
rect 305821 57835 305887 57836
rect 310973 57835 311039 57836
rect 313365 57835 313431 57836
rect 315021 57835 315087 57838
rect 318241 57835 318307 57838
rect 318374 57836 318380 57838
rect 318444 57836 318450 57900
rect 325877 57896 325986 57901
rect 343173 57900 343239 57901
rect 343449 57900 343515 57901
rect 343173 57898 343220 57900
rect 325877 57840 325882 57896
rect 325938 57840 325986 57896
rect 325877 57838 325986 57840
rect 343128 57896 343220 57898
rect 343128 57840 343178 57896
rect 343128 57838 343220 57840
rect 325877 57835 325943 57838
rect 343173 57836 343220 57838
rect 343284 57836 343290 57900
rect 343398 57898 343404 57900
rect 343358 57838 343404 57898
rect 343468 57896 343515 57900
rect 343510 57840 343515 57896
rect 343398 57836 343404 57838
rect 343468 57836 343515 57840
rect 343173 57835 343239 57836
rect 343449 57835 343515 57836
rect 398833 57898 398899 57901
rect 400397 57900 400463 57901
rect 399518 57898 399524 57900
rect 398833 57896 399524 57898
rect 398833 57840 398838 57896
rect 398894 57840 399524 57896
rect 398833 57838 399524 57840
rect 398833 57835 398899 57838
rect 399518 57836 399524 57838
rect 399588 57836 399594 57900
rect 400397 57896 400444 57900
rect 400508 57898 400514 57900
rect 401593 57898 401659 57901
rect 401734 57898 401794 58108
rect 400397 57840 400402 57896
rect 400397 57836 400444 57840
rect 400508 57838 400554 57898
rect 401593 57896 401794 57898
rect 401593 57840 401598 57896
rect 401654 57840 401794 57896
rect 401593 57838 401794 57840
rect 404077 57900 404143 57901
rect 404077 57896 404124 57900
rect 404188 57898 404194 57900
rect 404353 57898 404419 57901
rect 405038 57898 405044 57900
rect 404077 57840 404082 57896
rect 400508 57836 400514 57838
rect 400397 57835 400463 57836
rect 401593 57835 401659 57838
rect 404077 57836 404124 57840
rect 404188 57838 404234 57898
rect 404353 57896 405044 57898
rect 404353 57840 404358 57896
rect 404414 57840 405044 57896
rect 404353 57838 405044 57840
rect 404188 57836 404194 57838
rect 404077 57835 404143 57836
rect 404353 57835 404419 57838
rect 405038 57836 405044 57838
rect 405108 57836 405114 57900
rect 405825 57898 405891 57901
rect 406510 57898 406516 57900
rect 405825 57896 406516 57898
rect 405825 57840 405830 57896
rect 405886 57840 406516 57896
rect 405825 57838 406516 57840
rect 405825 57835 405891 57838
rect 406510 57836 406516 57838
rect 406580 57836 406586 57900
rect 407113 57898 407179 57901
rect 408309 57900 408375 57901
rect 408677 57900 408743 57901
rect 407614 57898 407620 57900
rect 407113 57896 407620 57898
rect 407113 57840 407118 57896
rect 407174 57840 407620 57896
rect 407113 57838 407620 57840
rect 407113 57835 407179 57838
rect 407614 57836 407620 57838
rect 407684 57836 407690 57900
rect 408309 57896 408356 57900
rect 408420 57898 408426 57900
rect 408309 57840 408314 57896
rect 408309 57836 408356 57840
rect 408420 57838 408466 57898
rect 408677 57896 408724 57900
rect 408788 57898 408794 57900
rect 409873 57898 409939 57901
rect 410006 57898 410012 57900
rect 408677 57840 408682 57896
rect 408420 57836 408426 57838
rect 408677 57836 408724 57840
rect 408788 57838 408834 57898
rect 409873 57896 410012 57898
rect 409873 57840 409878 57896
rect 409934 57840 410012 57896
rect 409873 57838 410012 57840
rect 408788 57836 408794 57838
rect 408309 57835 408375 57836
rect 408677 57835 408743 57836
rect 409873 57835 409939 57838
rect 410006 57836 410012 57838
rect 410076 57836 410082 57900
rect 411345 57898 411411 57901
rect 413461 57900 413527 57901
rect 414565 57900 414631 57901
rect 418429 57900 418495 57901
rect 422845 57900 422911 57901
rect 412398 57898 412404 57900
rect 411345 57896 412404 57898
rect 411345 57840 411350 57896
rect 411406 57840 412404 57896
rect 411345 57838 412404 57840
rect 411345 57835 411411 57838
rect 412398 57836 412404 57838
rect 412468 57836 412474 57900
rect 413461 57896 413508 57900
rect 413572 57898 413578 57900
rect 413461 57840 413466 57896
rect 413461 57836 413508 57840
rect 413572 57838 413618 57898
rect 414565 57896 414612 57900
rect 414676 57898 414682 57900
rect 414565 57840 414570 57896
rect 413572 57836 413578 57838
rect 414565 57836 414612 57840
rect 414676 57838 414722 57898
rect 418429 57896 418476 57900
rect 418540 57898 418546 57900
rect 418429 57840 418434 57896
rect 414676 57836 414682 57838
rect 418429 57836 418476 57840
rect 418540 57838 418586 57898
rect 422845 57896 422892 57900
rect 422956 57898 422962 57900
rect 423673 57898 423739 57901
rect 423990 57898 423996 57900
rect 422845 57840 422850 57896
rect 418540 57836 418546 57838
rect 422845 57836 422892 57840
rect 422956 57838 423002 57898
rect 423673 57896 423996 57898
rect 423673 57840 423678 57896
rect 423734 57840 423996 57896
rect 423673 57838 423996 57840
rect 422956 57836 422962 57838
rect 413461 57835 413527 57836
rect 414565 57835 414631 57836
rect 418429 57835 418495 57836
rect 422845 57835 422911 57836
rect 423673 57835 423739 57838
rect 423990 57836 423996 57838
rect 424060 57836 424066 57900
rect 426382 57836 426388 57900
rect 426452 57898 426458 57900
rect 426525 57898 426591 57901
rect 427629 57900 427695 57901
rect 427629 57898 427676 57900
rect 426452 57896 426591 57898
rect 426452 57840 426530 57896
rect 426586 57840 426591 57896
rect 426452 57838 426591 57840
rect 427584 57896 427676 57898
rect 427584 57840 427634 57896
rect 427584 57838 427676 57840
rect 426452 57836 426458 57838
rect 426525 57835 426591 57838
rect 427629 57836 427676 57838
rect 427740 57836 427746 57900
rect 427813 57898 427879 57901
rect 429653 57900 429719 57901
rect 430941 57900 431007 57901
rect 428590 57898 428596 57900
rect 427813 57896 428596 57898
rect 427813 57840 427818 57896
rect 427874 57840 428596 57896
rect 427813 57838 428596 57840
rect 427629 57835 427695 57836
rect 427813 57835 427879 57838
rect 428590 57836 428596 57838
rect 428660 57836 428666 57900
rect 429653 57896 429700 57900
rect 429764 57898 429770 57900
rect 429653 57840 429658 57896
rect 429653 57836 429700 57840
rect 429764 57838 429810 57898
rect 430941 57896 430988 57900
rect 431052 57898 431058 57900
rect 431953 57898 432019 57901
rect 433333 57900 433399 57901
rect 433517 57900 433583 57901
rect 432270 57898 432276 57900
rect 430941 57840 430946 57896
rect 429764 57836 429770 57838
rect 430941 57836 430988 57840
rect 431052 57838 431098 57898
rect 431953 57896 432276 57898
rect 431953 57840 431958 57896
rect 432014 57840 432276 57896
rect 431953 57838 432276 57840
rect 431052 57836 431058 57838
rect 429653 57835 429719 57836
rect 430941 57835 431007 57836
rect 431953 57835 432019 57838
rect 432270 57836 432276 57838
rect 432340 57836 432346 57900
rect 433333 57898 433380 57900
rect 433288 57896 433380 57898
rect 433288 57840 433338 57896
rect 433288 57838 433380 57840
rect 433333 57836 433380 57838
rect 433444 57836 433450 57900
rect 433517 57896 433564 57900
rect 433628 57898 433634 57900
rect 435081 57898 435147 57901
rect 435909 57900 435975 57901
rect 438485 57900 438551 57901
rect 435766 57898 435772 57900
rect 433517 57840 433522 57896
rect 433517 57836 433564 57840
rect 433628 57838 433674 57898
rect 435081 57896 435772 57898
rect 435081 57840 435086 57896
rect 435142 57840 435772 57896
rect 435081 57838 435772 57840
rect 433628 57836 433634 57838
rect 433333 57835 433399 57836
rect 433517 57835 433583 57836
rect 435081 57835 435147 57838
rect 435766 57836 435772 57838
rect 435836 57836 435842 57900
rect 435909 57896 435956 57900
rect 436020 57898 436026 57900
rect 435909 57840 435914 57896
rect 435909 57836 435956 57840
rect 436020 57838 436066 57898
rect 438485 57896 438532 57900
rect 438596 57898 438602 57900
rect 455830 57898 455890 58108
rect 438485 57840 438490 57896
rect 436020 57836 436026 57838
rect 438485 57836 438532 57840
rect 438596 57838 438642 57898
rect 451230 57838 455890 57898
rect 460933 57900 460999 57901
rect 465901 57900 465967 57901
rect 470869 57900 470935 57901
rect 475837 57900 475903 57901
rect 480621 57900 480687 57901
rect 483381 57900 483447 57901
rect 503345 57900 503411 57901
rect 460933 57896 460980 57900
rect 461044 57898 461050 57900
rect 460933 57840 460938 57896
rect 438596 57836 438602 57838
rect 435909 57835 435975 57836
rect 438485 57835 438551 57836
rect 263593 57764 263659 57765
rect 263542 57762 263548 57764
rect 206204 57702 258090 57762
rect 263502 57702 263548 57762
rect 263612 57760 263659 57764
rect 263654 57704 263659 57760
rect 206204 57700 206210 57702
rect 263542 57700 263548 57702
rect 263612 57700 263659 57704
rect 183185 57699 183251 57700
rect 263593 57699 263659 57700
rect 265433 57762 265499 57765
rect 265934 57762 265940 57764
rect 265433 57760 265940 57762
rect 265433 57704 265438 57760
rect 265494 57704 265940 57760
rect 265433 57702 265940 57704
rect 265433 57699 265499 57702
rect 265934 57700 265940 57702
rect 266004 57700 266010 57764
rect 266445 57762 266511 57765
rect 267590 57762 267596 57764
rect 266445 57760 267596 57762
rect 266445 57704 266450 57760
rect 266506 57704 267596 57760
rect 266445 57702 267596 57704
rect 266445 57699 266511 57702
rect 267590 57700 267596 57702
rect 267660 57700 267666 57764
rect 268193 57762 268259 57765
rect 268653 57764 268719 57765
rect 268326 57762 268332 57764
rect 268193 57760 268332 57762
rect 268193 57704 268198 57760
rect 268254 57704 268332 57760
rect 268193 57702 268332 57704
rect 268193 57699 268259 57702
rect 268326 57700 268332 57702
rect 268396 57700 268402 57764
rect 268653 57760 268700 57764
rect 268764 57762 268770 57764
rect 269113 57762 269179 57765
rect 269798 57762 269804 57764
rect 268653 57704 268658 57760
rect 268653 57700 268700 57704
rect 268764 57702 268810 57762
rect 269113 57760 269804 57762
rect 269113 57704 269118 57760
rect 269174 57704 269804 57760
rect 269113 57702 269804 57704
rect 268764 57700 268770 57702
rect 268653 57699 268719 57700
rect 269113 57699 269179 57702
rect 269798 57700 269804 57702
rect 269868 57700 269874 57764
rect 273345 57762 273411 57765
rect 274398 57762 274404 57764
rect 273345 57760 274404 57762
rect 273345 57704 273350 57760
rect 273406 57704 274404 57760
rect 273345 57702 274404 57704
rect 273345 57699 273411 57702
rect 274398 57700 274404 57702
rect 274468 57700 274474 57764
rect 276013 57762 276079 57765
rect 276974 57762 276980 57764
rect 276013 57760 276980 57762
rect 276013 57704 276018 57760
rect 276074 57704 276980 57760
rect 276013 57702 276980 57704
rect 276013 57699 276079 57702
rect 276974 57700 276980 57702
rect 277044 57700 277050 57764
rect 372102 57700 372108 57764
rect 372172 57762 372178 57764
rect 451230 57762 451290 57838
rect 460933 57836 460980 57840
rect 461044 57838 461090 57898
rect 465901 57896 465948 57900
rect 466012 57898 466018 57900
rect 465901 57840 465906 57896
rect 461044 57836 461050 57838
rect 465901 57836 465948 57840
rect 466012 57838 466058 57898
rect 470869 57896 470916 57900
rect 470980 57898 470986 57900
rect 470869 57840 470874 57896
rect 466012 57836 466018 57838
rect 470869 57836 470916 57840
rect 470980 57838 471026 57898
rect 475837 57896 475884 57900
rect 475948 57898 475954 57900
rect 475837 57840 475842 57896
rect 470980 57836 470986 57838
rect 475837 57836 475884 57840
rect 475948 57838 475994 57898
rect 480621 57896 480668 57900
rect 480732 57898 480738 57900
rect 480621 57840 480626 57896
rect 475948 57836 475954 57838
rect 480621 57836 480668 57840
rect 480732 57838 480778 57898
rect 483381 57896 483428 57900
rect 483492 57898 483498 57900
rect 503294 57898 503300 57900
rect 483381 57840 483386 57896
rect 480732 57836 480738 57838
rect 483381 57836 483428 57840
rect 483492 57838 483538 57898
rect 503254 57838 503300 57898
rect 503364 57896 503411 57900
rect 503406 57840 503411 57896
rect 483492 57836 483498 57838
rect 503294 57836 503300 57838
rect 503364 57836 503411 57840
rect 460933 57835 460999 57836
rect 465901 57835 465967 57836
rect 470869 57835 470935 57836
rect 475837 57835 475903 57836
rect 480621 57835 480687 57836
rect 483381 57835 483447 57836
rect 503345 57835 503411 57836
rect 372172 57702 451290 57762
rect 372172 57700 372178 57702
rect 54886 57564 54892 57628
rect 54956 57626 54962 57628
rect 114553 57626 114619 57629
rect 115790 57626 115796 57628
rect 54956 57566 114468 57626
rect 54956 57564 54962 57566
rect 58934 57428 58940 57492
rect 59004 57490 59010 57492
rect 98637 57490 98703 57493
rect 59004 57488 98703 57490
rect 59004 57432 98642 57488
rect 98698 57432 98703 57488
rect 59004 57430 98703 57432
rect 59004 57428 59010 57430
rect 98637 57427 98703 57430
rect 111793 57490 111859 57493
rect 113173 57492 113239 57493
rect 112110 57490 112116 57492
rect 111793 57488 112116 57490
rect 111793 57432 111798 57488
rect 111854 57432 112116 57488
rect 111793 57430 112116 57432
rect 111793 57427 111859 57430
rect 112110 57428 112116 57430
rect 112180 57428 112186 57492
rect 113173 57488 113220 57492
rect 113284 57490 113290 57492
rect 114408 57490 114468 57566
rect 114553 57624 115796 57626
rect 114553 57568 114558 57624
rect 114614 57568 115796 57624
rect 114553 57566 115796 57568
rect 114553 57563 114619 57566
rect 115790 57564 115796 57566
rect 115860 57564 115866 57628
rect 118693 57626 118759 57629
rect 155953 57628 156019 57629
rect 119102 57626 119108 57628
rect 118693 57624 119108 57626
rect 118693 57568 118698 57624
rect 118754 57568 119108 57624
rect 118693 57566 119108 57568
rect 118693 57563 118759 57566
rect 119102 57564 119108 57566
rect 119172 57564 119178 57628
rect 155902 57626 155908 57628
rect 155862 57566 155908 57626
rect 155972 57624 156019 57628
rect 156014 57568 156019 57624
rect 155902 57564 155908 57566
rect 155972 57564 156019 57568
rect 155953 57563 156019 57564
rect 160093 57626 160159 57629
rect 160870 57626 160876 57628
rect 160093 57624 160876 57626
rect 160093 57568 160098 57624
rect 160154 57568 160876 57624
rect 160093 57566 160876 57568
rect 160093 57563 160159 57566
rect 160870 57564 160876 57566
rect 160940 57564 160946 57628
rect 165613 57626 165679 57629
rect 165838 57626 165844 57628
rect 165613 57624 165844 57626
rect 165613 57568 165618 57624
rect 165674 57568 165844 57624
rect 165613 57566 165844 57568
rect 165613 57563 165679 57566
rect 165838 57564 165844 57566
rect 165908 57564 165914 57628
rect 215886 57564 215892 57628
rect 215956 57626 215962 57628
rect 280838 57626 280844 57628
rect 215956 57566 280844 57626
rect 215956 57564 215962 57566
rect 280838 57564 280844 57566
rect 280908 57564 280914 57628
rect 370446 57564 370452 57628
rect 370516 57626 370522 57628
rect 451038 57626 451044 57628
rect 370516 57566 451044 57626
rect 370516 57564 370522 57566
rect 451038 57564 451044 57566
rect 451108 57564 451114 57628
rect 118366 57490 118372 57492
rect 113173 57432 113178 57488
rect 113173 57428 113220 57432
rect 113284 57430 113330 57490
rect 114408 57430 118372 57490
rect 113284 57428 113290 57430
rect 118366 57428 118372 57430
rect 118436 57428 118442 57492
rect 213126 57428 213132 57492
rect 213196 57490 213202 57492
rect 273478 57490 273484 57492
rect 213196 57430 273484 57490
rect 213196 57428 213202 57430
rect 273478 57428 273484 57430
rect 273548 57428 273554 57492
rect 360694 57428 360700 57492
rect 360764 57490 360770 57492
rect 433425 57490 433491 57493
rect 360764 57488 433491 57490
rect 360764 57432 433430 57488
rect 433486 57432 433491 57488
rect 360764 57430 433491 57432
rect 360764 57428 360770 57430
rect 113173 57427 113239 57428
rect 433425 57427 433491 57430
rect 433701 57490 433767 57493
rect 434662 57490 434668 57492
rect 433701 57488 434668 57490
rect 433701 57432 433706 57488
rect 433762 57432 434668 57488
rect 433701 57430 434668 57432
rect 433701 57427 433767 57430
rect 434662 57428 434668 57430
rect 434732 57428 434738 57492
rect 436093 57490 436159 57493
rect 436870 57490 436876 57492
rect 436093 57488 436876 57490
rect 436093 57432 436098 57488
rect 436154 57432 436876 57488
rect 436093 57430 436876 57432
rect 436093 57427 436159 57430
rect 436870 57428 436876 57430
rect 436940 57428 436946 57492
rect 438853 57490 438919 57493
rect 439078 57490 439084 57492
rect 438853 57488 439084 57490
rect 438853 57432 438858 57488
rect 438914 57432 439084 57488
rect 438853 57430 439084 57432
rect 438853 57427 438919 57430
rect 439078 57428 439084 57430
rect 439148 57428 439154 57492
rect 266353 57356 266419 57357
rect 58566 57292 58572 57356
rect 58636 57354 58642 57356
rect 103830 57354 103836 57356
rect 58636 57294 103836 57354
rect 58636 57292 58642 57294
rect 103830 57292 103836 57294
rect 103900 57292 103906 57356
rect 202270 57292 202276 57356
rect 202340 57354 202346 57356
rect 260966 57354 260972 57356
rect 202340 57294 260972 57354
rect 202340 57292 202346 57294
rect 260966 57292 260972 57294
rect 261036 57292 261042 57356
rect 266302 57354 266308 57356
rect 266262 57294 266308 57354
rect 266372 57352 266419 57356
rect 266414 57296 266419 57352
rect 266302 57292 266308 57294
rect 266372 57292 266419 57296
rect 376150 57292 376156 57356
rect 376220 57354 376226 57356
rect 448278 57354 448284 57356
rect 376220 57294 448284 57354
rect 376220 57292 376226 57294
rect 448278 57292 448284 57294
rect 448348 57292 448354 57356
rect 266353 57291 266419 57292
rect 57646 57156 57652 57220
rect 57716 57218 57722 57220
rect 98637 57218 98703 57221
rect 105854 57218 105860 57220
rect 57716 57158 93870 57218
rect 57716 57156 57722 57158
rect 88425 57084 88491 57085
rect 58750 57020 58756 57084
rect 58820 57082 58826 57084
rect 88374 57082 88380 57084
rect 58820 57022 84210 57082
rect 88334 57022 88380 57082
rect 88444 57080 88491 57084
rect 88486 57024 88491 57080
rect 58820 57020 58826 57022
rect 84150 56946 84210 57022
rect 88374 57020 88380 57022
rect 88444 57020 88491 57024
rect 93810 57082 93870 57158
rect 98637 57216 105860 57218
rect 98637 57160 98642 57216
rect 98698 57160 105860 57216
rect 98637 57158 105860 57160
rect 98637 57155 98703 57158
rect 105854 57156 105860 57158
rect 105924 57156 105930 57220
rect 203190 57156 203196 57220
rect 203260 57218 203266 57220
rect 255998 57218 256004 57220
rect 203260 57158 256004 57218
rect 203260 57156 203266 57158
rect 255998 57156 256004 57158
rect 256068 57156 256074 57220
rect 378726 57156 378732 57220
rect 378796 57218 378802 57220
rect 445886 57218 445892 57220
rect 378796 57158 445892 57218
rect 378796 57156 378802 57158
rect 445886 57156 445892 57158
rect 445956 57156 445962 57220
rect 97022 57082 97028 57084
rect 93810 57022 97028 57082
rect 97022 57020 97028 57022
rect 97092 57020 97098 57084
rect 216070 57020 216076 57084
rect 216140 57082 216146 57084
rect 253606 57082 253612 57084
rect 216140 57022 253612 57082
rect 216140 57020 216146 57022
rect 253606 57020 253612 57022
rect 253676 57020 253682 57084
rect 376334 57020 376340 57084
rect 376404 57082 376410 57084
rect 415526 57082 415532 57084
rect 376404 57022 415532 57082
rect 376404 57020 376410 57022
rect 415526 57020 415532 57022
rect 415596 57020 415602 57084
rect 430573 57082 430639 57085
rect 431166 57082 431172 57084
rect 430573 57080 431172 57082
rect 430573 57024 430578 57080
rect 430634 57024 431172 57080
rect 430573 57022 431172 57024
rect 88425 57019 88491 57020
rect 430573 57019 430639 57022
rect 431166 57020 431172 57022
rect 431236 57020 431242 57084
rect 433425 57082 433491 57085
rect 440918 57082 440924 57084
rect 433425 57080 440924 57082
rect 433425 57024 433430 57080
rect 433486 57024 440924 57080
rect 433425 57022 440924 57024
rect 433425 57019 433491 57022
rect 440918 57020 440924 57022
rect 440988 57020 440994 57084
rect 96286 56946 96292 56948
rect 84150 56886 96292 56946
rect 96286 56884 96292 56886
rect 96356 56884 96362 56948
rect 235993 56946 236059 56949
rect 411253 56948 411319 56949
rect 237046 56946 237052 56948
rect 235993 56944 237052 56946
rect 235993 56888 235998 56944
rect 236054 56888 237052 56944
rect 235993 56886 237052 56888
rect 235993 56883 236059 56886
rect 237046 56884 237052 56886
rect 237116 56884 237122 56948
rect 411253 56944 411300 56948
rect 411364 56946 411370 56948
rect 411253 56888 411258 56944
rect 411253 56884 411300 56888
rect 411364 56886 411410 56946
rect 411364 56884 411370 56886
rect 411253 56883 411319 56884
rect 443494 56810 443500 56812
rect 431910 56750 443500 56810
rect 52310 56612 52316 56676
rect 52380 56674 52386 56676
rect 133454 56674 133460 56676
rect 52380 56614 133460 56674
rect 52380 56612 52386 56614
rect 133454 56612 133460 56614
rect 133524 56612 133530 56676
rect 163262 56612 163268 56676
rect 163332 56612 163338 56676
rect 211654 56612 211660 56676
rect 211724 56674 211730 56676
rect 285990 56674 285996 56676
rect 211724 56614 285996 56674
rect 211724 56612 211730 56614
rect 285990 56612 285996 56614
rect 286060 56612 286066 56676
rect 320950 56612 320956 56676
rect 321020 56612 321026 56676
rect 323342 56612 323348 56676
rect 323412 56612 323418 56676
rect 358118 56612 358124 56676
rect 358188 56674 358194 56676
rect 431910 56674 431970 56750
rect 443494 56748 443500 56750
rect 443564 56748 443570 56812
rect 358188 56614 431970 56674
rect 358188 56612 358194 56614
rect 438342 56612 438348 56676
rect 438412 56612 438418 56676
rect 53598 56476 53604 56540
rect 53668 56538 53674 56540
rect 163270 56538 163330 56612
rect 53668 56478 163330 56538
rect 53668 56476 53674 56478
rect 205398 56476 205404 56540
rect 205468 56538 205474 56540
rect 320958 56538 321018 56612
rect 205468 56478 321018 56538
rect 205468 56476 205474 56478
rect 48630 56340 48636 56404
rect 48700 56402 48706 56404
rect 158478 56402 158484 56404
rect 48700 56342 158484 56402
rect 48700 56340 48706 56342
rect 158478 56340 158484 56342
rect 158548 56340 158554 56404
rect 209630 56340 209636 56404
rect 209700 56402 209706 56404
rect 323350 56402 323410 56612
rect 377254 56476 377260 56540
rect 377324 56538 377330 56540
rect 438350 56538 438410 56612
rect 377324 56478 438410 56538
rect 377324 56476 377330 56478
rect 209700 56342 323410 56402
rect 209700 56340 209706 56342
rect 52126 56204 52132 56268
rect 52196 56266 52202 56268
rect 153285 56266 153351 56269
rect 52196 56264 153351 56266
rect 52196 56208 153290 56264
rect 153346 56208 153351 56264
rect 52196 56206 153351 56208
rect 52196 56204 52202 56206
rect 153285 56203 153351 56206
rect 206870 56204 206876 56268
rect 206940 56266 206946 56268
rect 315021 56266 315087 56269
rect 206940 56264 315087 56266
rect 206940 56208 315026 56264
rect 315082 56208 315087 56264
rect 206940 56206 315087 56208
rect 206940 56204 206946 56206
rect 315021 56203 315087 56206
rect 57830 56068 57836 56132
rect 57900 56130 57906 56132
rect 116485 56130 116551 56133
rect 57900 56128 116551 56130
rect 57900 56072 116490 56128
rect 116546 56072 116551 56128
rect 57900 56070 116551 56072
rect 57900 56068 57906 56070
rect 116485 56067 116551 56070
rect 197854 56068 197860 56132
rect 197924 56130 197930 56132
rect 265433 56130 265499 56133
rect 197924 56128 265499 56130
rect 197924 56072 265438 56128
rect 265494 56072 265499 56128
rect 197924 56070 265499 56072
rect 197924 56068 197930 56070
rect 265433 56067 265499 56070
rect 50654 55116 50660 55180
rect 50724 55178 50730 55180
rect 165613 55178 165679 55181
rect 50724 55176 165679 55178
rect 50724 55120 165618 55176
rect 165674 55120 165679 55176
rect 50724 55118 165679 55120
rect 50724 55116 50730 55118
rect 165613 55115 165679 55118
rect 212165 55178 212231 55181
rect 273345 55178 273411 55181
rect 212165 55176 273411 55178
rect 212165 55120 212170 55176
rect 212226 55120 273350 55176
rect 273406 55120 273411 55176
rect 212165 55118 273411 55120
rect 212165 55115 212231 55118
rect 273345 55115 273411 55118
rect 377806 55116 377812 55180
rect 377876 55178 377882 55180
rect 438853 55178 438919 55181
rect 377876 55176 438919 55178
rect 377876 55120 438858 55176
rect 438914 55120 438919 55176
rect 377876 55118 438919 55120
rect 377876 55116 377882 55118
rect 438853 55115 438919 55118
rect 50470 54980 50476 55044
rect 50540 55042 50546 55044
rect 160093 55042 160159 55045
rect 50540 55040 160159 55042
rect 50540 54984 160098 55040
rect 160154 54984 160159 55040
rect 50540 54982 160159 54984
rect 50540 54980 50546 54982
rect 160093 54979 160159 54982
rect 217358 54980 217364 55044
rect 217428 55042 217434 55044
rect 276013 55042 276079 55045
rect 217428 55040 276079 55042
rect 217428 54984 276018 55040
rect 276074 54984 276079 55040
rect 217428 54982 276079 54984
rect 217428 54980 217434 54982
rect 276013 54979 276079 54982
rect 379462 54980 379468 55044
rect 379532 55042 379538 55044
rect 427813 55042 427879 55045
rect 379532 55040 427879 55042
rect 379532 54984 427818 55040
rect 427874 54984 427879 55040
rect 379532 54982 427879 54984
rect 379532 54980 379538 54982
rect 427813 54979 427879 54982
rect 50838 54844 50844 54908
rect 50908 54906 50914 54908
rect 155953 54906 156019 54909
rect 50908 54904 156019 54906
rect 50908 54848 155958 54904
rect 156014 54848 156019 54904
rect 50908 54846 156019 54848
rect 50908 54844 50914 54846
rect 155953 54843 156019 54846
rect 57462 54708 57468 54772
rect 57532 54770 57538 54772
rect 118693 54770 118759 54773
rect 57532 54768 118759 54770
rect 57532 54712 118698 54768
rect 118754 54712 118759 54768
rect 57532 54710 118759 54712
rect 57532 54708 57538 54710
rect 118693 54707 118759 54710
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 580257 33146 580323 33149
rect 583520 33146 584960 33236
rect 580257 33144 584960 33146
rect 580257 33088 580262 33144
rect 580318 33088 584960 33144
rect 580257 33086 584960 33088
rect 580257 33083 580323 33086
rect 583520 32996 584960 33086
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19410 480 19500
rect 2773 19410 2839 19413
rect -960 19408 2839 19410
rect -960 19352 2778 19408
rect 2834 19352 2839 19408
rect -960 19350 2839 19352
rect -960 19260 480 19350
rect 2773 19347 2839 19350
rect -960 6340 480 6580
rect 583520 6476 584960 6716
rect 143533 4042 143599 4045
rect 208894 4042 208900 4044
rect 143533 4040 208900 4042
rect 143533 3984 143538 4040
rect 143594 3984 208900 4040
rect 143533 3982 208900 3984
rect 143533 3979 143599 3982
rect 208894 3980 208900 3982
rect 208964 3980 208970 4044
rect 136449 3906 136515 3909
rect 204846 3906 204852 3908
rect 136449 3904 204852 3906
rect 136449 3848 136454 3904
rect 136510 3848 204852 3904
rect 136449 3846 204852 3848
rect 136449 3843 136515 3846
rect 204846 3844 204852 3846
rect 204916 3844 204922 3908
rect 140037 3770 140103 3773
rect 210366 3770 210372 3772
rect 140037 3768 210372 3770
rect 140037 3712 140042 3768
rect 140098 3712 210372 3768
rect 140037 3710 210372 3712
rect 140037 3707 140103 3710
rect 210366 3708 210372 3710
rect 210436 3708 210442 3772
rect 150617 3634 150683 3637
rect 371734 3634 371740 3636
rect 150617 3632 371740 3634
rect 150617 3576 150622 3632
rect 150678 3576 371740 3632
rect 150617 3574 371740 3576
rect 150617 3571 150683 3574
rect 371734 3572 371740 3574
rect 371804 3572 371810 3636
rect 132953 3498 133019 3501
rect 363454 3498 363460 3500
rect 132953 3496 363460 3498
rect 132953 3440 132958 3496
rect 133014 3440 363460 3496
rect 132953 3438 363460 3440
rect 132953 3435 133019 3438
rect 363454 3436 363460 3438
rect 363524 3436 363530 3500
rect 129365 3362 129431 3365
rect 364926 3362 364932 3364
rect 129365 3360 364932 3362
rect 129365 3304 129370 3360
rect 129426 3304 364932 3360
rect 129365 3302 364932 3304
rect 129365 3299 129431 3302
rect 364926 3300 364932 3302
rect 364996 3300 365002 3364
<< via3 >>
rect 54340 646172 54404 646236
rect 51580 646036 51644 646100
rect 53052 645900 53116 645964
rect 476068 639916 476132 639980
rect 488580 639916 488644 639980
rect 506612 639916 506676 639980
rect 436140 606324 436204 606388
rect 436140 534516 436204 534580
rect 370636 529076 370700 529140
rect 371740 526356 371804 526420
rect 363460 496028 363524 496092
rect 476068 496028 476132 496092
rect 364932 493308 364996 493372
rect 208900 491812 208964 491876
rect 488580 491812 488644 491876
rect 60228 491132 60292 491196
rect 198228 491132 198292 491196
rect 216628 491132 216692 491196
rect 219940 491132 220004 491196
rect 357940 491132 358004 491196
rect 199332 490996 199396 491060
rect 202644 490996 202708 491060
rect 206692 490996 206756 491060
rect 216812 490996 216876 491060
rect 371924 490996 371988 491060
rect 54892 490860 54956 490924
rect 196572 490860 196636 490924
rect 201356 490860 201420 490924
rect 205220 490860 205284 490924
rect 367876 490860 367940 490924
rect 55076 490724 55140 490788
rect 197860 490724 197924 490788
rect 219020 490724 219084 490788
rect 367692 490724 367756 490788
rect 46796 490588 46860 490652
rect 200620 490588 200684 490652
rect 50844 490512 50908 490516
rect 50844 490456 50894 490512
rect 50894 490456 50908 490512
rect 50844 490452 50908 490456
rect 52316 490452 52380 490516
rect 202092 490452 202156 490516
rect 205404 490452 205468 490516
rect 213316 490588 213380 490652
rect 218836 490588 218900 490652
rect 374500 490588 374564 490652
rect 217548 490452 217612 490516
rect 219204 490452 219268 490516
rect 375972 490452 376036 490516
rect 59308 490316 59372 490380
rect 198044 490316 198108 490380
rect 200988 490316 201052 490380
rect 206876 490316 206940 490380
rect 209636 490316 209700 490380
rect 59124 490180 59188 490244
rect 198412 490180 198476 490244
rect 55628 490044 55692 490108
rect 213132 489092 213196 489156
rect 378916 489092 378980 489156
rect 57100 488276 57164 488340
rect 44036 487732 44100 487796
rect 358124 487732 358188 487796
rect 378732 486372 378796 486436
rect 209820 485012 209884 485076
rect 376156 485012 376220 485076
rect 207980 483788 208044 483852
rect 211660 483652 211724 483716
rect 360700 483652 360764 483716
rect 57468 482428 57532 482492
rect 211844 482428 211908 482492
rect 47716 482292 47780 482356
rect 214052 482292 214116 482356
rect 372660 482292 372724 482356
rect 44956 482156 45020 482220
rect 202276 482156 202340 482220
rect 210372 482156 210436 482220
rect 379468 481068 379532 481132
rect 215892 480932 215956 480996
rect 376340 480932 376404 480996
rect 204852 480796 204916 480860
rect 216076 479436 216140 479500
rect 378180 479436 378244 479500
rect 208348 478076 208412 478140
rect 359412 478076 359476 478140
rect 213868 476852 213932 476916
rect 206140 476716 206204 476780
rect 360148 476716 360212 476780
rect 377260 475492 377324 475556
rect 215340 475356 215404 475420
rect 372108 475356 372172 475420
rect 216260 474404 216324 474468
rect 203196 474268 203260 474332
rect 214236 474132 214300 474196
rect 196756 473996 196820 474060
rect 370452 473996 370516 474060
rect 506612 472636 506676 472700
rect 202460 472500 202524 472564
rect 378364 472500 378428 472564
rect 203012 471820 203076 471884
rect 44772 471684 44836 471748
rect 205036 471684 205100 471748
rect 57836 471548 57900 471612
rect 217180 471548 217244 471612
rect 359596 471412 359660 471476
rect 377444 471276 377508 471340
rect 47900 471140 47964 471204
rect 377628 471140 377692 471204
rect 58940 469780 59004 469844
rect 199516 468964 199580 469028
rect 48084 468828 48148 468892
rect 200804 468828 200868 468892
rect 46612 468692 46676 468756
rect 210556 468692 210620 468756
rect 53604 468556 53668 468620
rect 50660 468420 50724 468484
rect 359780 468420 359844 468484
rect 58756 467060 58820 467124
rect 206324 467060 206388 467124
rect 178356 466516 178420 466580
rect 179644 466516 179708 466580
rect 190868 466576 190932 466580
rect 190868 466520 190918 466576
rect 190918 466520 190932 466576
rect 190868 466516 190932 466520
rect 338436 466576 338500 466580
rect 338436 466520 338486 466576
rect 338486 466520 338500 466576
rect 338436 466516 338500 466520
rect 339724 466576 339788 466580
rect 339724 466520 339774 466576
rect 339774 466520 339788 466576
rect 339724 466516 339788 466520
rect 350948 466576 351012 466580
rect 350948 466520 350998 466576
rect 350998 466520 351012 466576
rect 350948 466516 351012 466520
rect 498516 466576 498580 466580
rect 498516 466520 498530 466576
rect 498530 466520 498580 466576
rect 498516 466516 498580 466520
rect 499804 466576 499868 466580
rect 499804 466520 499818 466576
rect 499818 466520 499868 466576
rect 499804 466516 499868 466520
rect 510844 466576 510908 466580
rect 510844 466520 510894 466576
rect 510894 466520 510908 466576
rect 510844 466516 510908 466520
rect 53420 466380 53484 466444
rect 54708 466244 54772 466308
rect 53236 466108 53300 466172
rect 198964 466108 199028 466172
rect 51948 465972 52012 466036
rect 208164 465972 208228 466036
rect 52132 465836 52196 465900
rect 377812 465836 377876 465900
rect 48636 465700 48700 465764
rect 198780 465700 198844 465764
rect 58572 465564 58636 465628
rect 50476 465156 50540 465220
rect 57652 464340 57716 464404
rect 359964 410484 360028 410548
rect 216812 396612 216876 396676
rect 57468 390628 57532 390692
rect 53236 388452 53300 388516
rect 55628 380972 55692 381036
rect 198412 380972 198476 381036
rect 200988 380972 201052 381036
rect 84214 380836 84278 380900
rect 83126 380700 83190 380764
rect 217548 380700 217612 380764
rect 323366 380836 323430 380900
rect 413598 380896 413662 380900
rect 413598 380840 413614 380896
rect 413614 380840 413662 380896
rect 413598 380836 413662 380840
rect 421078 380896 421142 380900
rect 421078 380840 421102 380896
rect 421102 380840 421142 380896
rect 421078 380836 421142 380840
rect 425974 380896 426038 380900
rect 425974 380840 425978 380896
rect 425978 380840 426034 380896
rect 426034 380840 426038 380896
rect 425974 380836 426038 380840
rect 433590 380896 433654 380900
rect 433590 380840 433614 380896
rect 433614 380840 433654 380896
rect 433590 380836 433654 380840
rect 436038 380896 436102 380900
rect 436038 380840 436062 380896
rect 436062 380840 436102 380896
rect 436038 380836 436102 380840
rect 236054 380700 236118 380764
rect 237142 380760 237206 380764
rect 237142 380704 237158 380760
rect 237158 380704 237206 380760
rect 237142 380700 237206 380704
rect 243126 380760 243190 380764
rect 243126 380704 243138 380760
rect 243138 380704 243190 380760
rect 243126 380700 243190 380704
rect 248294 380700 248358 380764
rect 254550 380700 254614 380764
rect 255910 380760 255974 380764
rect 255910 380704 255926 380760
rect 255926 380704 255974 380760
rect 255910 380700 255974 380704
rect 313438 380760 313502 380764
rect 313438 380704 313462 380760
rect 313462 380704 313502 380760
rect 313438 380700 313502 380704
rect 438486 380760 438550 380764
rect 438486 380704 438490 380760
rect 438490 380704 438546 380760
rect 438546 380704 438550 380760
rect 438486 380700 438550 380704
rect 440934 380760 440998 380764
rect 440934 380704 440938 380760
rect 440938 380704 440998 380760
rect 440934 380700 440998 380704
rect 443518 380700 443582 380764
rect 448278 380760 448342 380764
rect 448278 380704 448298 380760
rect 448298 380704 448342 380760
rect 448278 380700 448342 380704
rect 94550 380564 94614 380628
rect 95924 380292 95988 380356
rect 111012 380352 111076 380356
rect 111012 380296 111026 380352
rect 111026 380296 111076 380352
rect 111012 380292 111076 380296
rect 113588 380352 113652 380356
rect 113588 380296 113602 380352
rect 113602 380296 113652 380352
rect 113588 380292 113652 380296
rect 115980 380352 116044 380356
rect 115980 380296 115994 380352
rect 115994 380296 116044 380352
rect 115980 380292 116044 380296
rect 118372 380352 118436 380356
rect 118372 380296 118386 380352
rect 118386 380296 118436 380352
rect 118372 380292 118436 380296
rect 120948 380352 121012 380356
rect 120948 380296 120998 380352
rect 120998 380296 121012 380352
rect 120948 380292 121012 380296
rect 123524 380352 123588 380356
rect 123524 380296 123538 380352
rect 123538 380296 123588 380352
rect 123524 380292 123588 380296
rect 128308 380352 128372 380356
rect 128308 380296 128358 380352
rect 128358 380296 128372 380352
rect 128308 380292 128372 380296
rect 135852 380352 135916 380356
rect 135852 380296 135902 380352
rect 135902 380296 135916 380352
rect 135852 380292 135916 380296
rect 143580 380352 143644 380356
rect 143580 380296 143630 380352
rect 143630 380296 143644 380352
rect 143580 380292 143644 380296
rect 148548 380352 148612 380356
rect 148548 380296 148598 380352
rect 148598 380296 148612 380352
rect 148548 380292 148612 380296
rect 155908 380352 155972 380356
rect 155908 380296 155958 380352
rect 155958 380296 155972 380352
rect 155908 380292 155972 380296
rect 158484 380352 158548 380356
rect 158484 380296 158534 380352
rect 158534 380296 158548 380352
rect 158484 380292 158548 380296
rect 160876 380352 160940 380356
rect 160876 380296 160926 380352
rect 160926 380296 160940 380352
rect 160876 380292 160940 380296
rect 163452 380352 163516 380356
rect 163452 380296 163502 380352
rect 163502 380296 163516 380352
rect 163452 380292 163516 380296
rect 166028 380352 166092 380356
rect 166028 380296 166078 380352
rect 166078 380296 166092 380352
rect 166028 380292 166092 380296
rect 216628 380156 216692 380220
rect 256998 380564 257062 380628
rect 258086 380624 258150 380628
rect 258086 380568 258134 380624
rect 258134 380568 258150 380624
rect 258086 380564 258150 380568
rect 261758 380624 261822 380628
rect 261758 380568 261814 380624
rect 261814 380568 261822 380624
rect 261758 380564 261822 380568
rect 271006 380624 271070 380628
rect 271006 380568 271014 380624
rect 271014 380568 271070 380624
rect 271006 380564 271070 380568
rect 315886 380624 315950 380628
rect 315886 380568 315910 380624
rect 315910 380568 315950 380624
rect 315886 380564 315950 380568
rect 404214 380624 404278 380628
rect 404214 380568 404230 380624
rect 404230 380568 404278 380624
rect 404214 380564 404278 380568
rect 405438 380624 405502 380628
rect 405438 380568 405462 380624
rect 405462 380568 405502 380624
rect 405438 380564 405502 380568
rect 413462 380624 413526 380628
rect 413462 380568 413466 380624
rect 413466 380568 413522 380624
rect 413522 380568 413526 380624
rect 413462 380564 413526 380568
rect 445966 380624 446030 380628
rect 445966 380568 445998 380624
rect 445998 380568 446030 380624
rect 445966 380564 446030 380568
rect 503358 380624 503422 380628
rect 503358 380568 503406 380624
rect 503406 380568 503422 380624
rect 503358 380564 503422 380568
rect 244228 380488 244292 380492
rect 244228 380432 244278 380488
rect 244278 380432 244292 380488
rect 244228 380428 244292 380432
rect 247540 380292 247604 380356
rect 359596 380156 359660 380220
rect 427492 380156 427556 380220
rect 259500 380020 259564 380084
rect 217364 379672 217428 379676
rect 217364 379616 217378 379672
rect 217378 379616 217428 379672
rect 217364 379612 217428 379616
rect 51948 379476 52012 379540
rect 209820 379476 209884 379540
rect 218836 379476 218900 379540
rect 360148 379476 360212 379540
rect 77156 379400 77220 379404
rect 77156 379344 77206 379400
rect 77206 379344 77220 379400
rect 77156 379340 77220 379344
rect 80468 379400 80532 379404
rect 80468 379344 80482 379400
rect 80482 379344 80532 379400
rect 80468 379340 80532 379344
rect 85436 379400 85500 379404
rect 85436 379344 85486 379400
rect 85486 379344 85500 379400
rect 85436 379340 85500 379344
rect 86540 379400 86604 379404
rect 86540 379344 86590 379400
rect 86590 379344 86604 379400
rect 86540 379340 86604 379344
rect 88380 379400 88444 379404
rect 88380 379344 88394 379400
rect 88394 379344 88444 379400
rect 88380 379340 88444 379344
rect 88748 379400 88812 379404
rect 88748 379344 88798 379400
rect 88798 379344 88812 379400
rect 88748 379340 88812 379344
rect 90772 379400 90836 379404
rect 90772 379344 90786 379400
rect 90786 379344 90836 379400
rect 90772 379340 90836 379344
rect 91324 379400 91388 379404
rect 91324 379344 91374 379400
rect 91374 379344 91388 379400
rect 91324 379340 91388 379344
rect 92428 379400 92492 379404
rect 92428 379344 92442 379400
rect 92442 379344 92492 379400
rect 92428 379340 92492 379344
rect 93348 379340 93412 379404
rect 96108 379400 96172 379404
rect 96108 379344 96122 379400
rect 96122 379344 96172 379400
rect 96108 379340 96172 379344
rect 98500 379400 98564 379404
rect 98500 379344 98514 379400
rect 98514 379344 98564 379400
rect 98500 379340 98564 379344
rect 101076 379400 101140 379404
rect 101076 379344 101090 379400
rect 101090 379344 101140 379400
rect 101076 379340 101140 379344
rect 103284 379340 103348 379404
rect 105860 379340 105924 379404
rect 108252 379400 108316 379404
rect 108252 379344 108266 379400
rect 108266 379344 108316 379400
rect 108252 379340 108316 379344
rect 108804 379400 108868 379404
rect 108804 379344 108854 379400
rect 108854 379344 108868 379400
rect 108804 379340 108868 379344
rect 109724 379400 109788 379404
rect 109724 379344 109774 379400
rect 109774 379344 109788 379400
rect 109724 379340 109788 379344
rect 111196 379400 111260 379404
rect 111196 379344 111246 379400
rect 111246 379344 111260 379400
rect 111196 379340 111260 379344
rect 112300 379400 112364 379404
rect 112300 379344 112350 379400
rect 112350 379344 112364 379400
rect 112300 379340 112364 379344
rect 113404 379400 113468 379404
rect 113404 379344 113454 379400
rect 113454 379344 113468 379400
rect 113404 379340 113468 379344
rect 114508 379400 114572 379404
rect 114508 379344 114522 379400
rect 114522 379344 114572 379400
rect 114508 379340 114572 379344
rect 115796 379400 115860 379404
rect 115796 379344 115846 379400
rect 115846 379344 115860 379400
rect 115796 379340 115860 379344
rect 117084 379400 117148 379404
rect 117084 379344 117134 379400
rect 117134 379344 117148 379400
rect 117084 379340 117148 379344
rect 141004 379400 141068 379404
rect 141004 379344 141054 379400
rect 141054 379344 141068 379400
rect 141004 379340 141068 379344
rect 145972 379400 146036 379404
rect 145972 379344 146022 379400
rect 146022 379344 146036 379400
rect 145972 379340 146036 379344
rect 150940 379400 151004 379404
rect 150940 379344 150990 379400
rect 150990 379344 151004 379400
rect 150940 379340 151004 379344
rect 153516 379400 153580 379404
rect 153516 379344 153566 379400
rect 153566 379344 153580 379400
rect 153516 379340 153580 379344
rect 239628 379400 239692 379404
rect 239628 379344 239642 379400
rect 239642 379344 239692 379400
rect 239628 379340 239692 379344
rect 245332 379340 245396 379404
rect 246436 379340 246500 379404
rect 248644 379400 248708 379404
rect 248644 379344 248658 379400
rect 248658 379344 248708 379400
rect 248644 379340 248708 379344
rect 250116 379400 250180 379404
rect 250116 379344 250130 379400
rect 250130 379344 250180 379400
rect 250116 379340 250180 379344
rect 251220 379400 251284 379404
rect 251220 379344 251234 379400
rect 251234 379344 251284 379400
rect 251220 379340 251284 379344
rect 252324 379400 252388 379404
rect 252324 379344 252338 379400
rect 252338 379344 252388 379400
rect 252324 379340 252388 379344
rect 253428 379400 253492 379404
rect 253428 379344 253442 379400
rect 253442 379344 253492 379400
rect 253428 379340 253492 379344
rect 263916 379400 263980 379404
rect 263916 379344 263930 379400
rect 263930 379344 263980 379400
rect 263916 379340 263980 379344
rect 265204 379340 265268 379404
rect 268700 379340 268764 379404
rect 269804 379400 269868 379404
rect 269804 379344 269818 379400
rect 269818 379344 269868 379400
rect 269804 379340 269868 379344
rect 271092 379400 271156 379404
rect 271092 379344 271106 379400
rect 271106 379344 271156 379400
rect 271092 379340 271156 379344
rect 272196 379400 272260 379404
rect 272196 379344 272210 379400
rect 272210 379344 272260 379400
rect 272196 379340 272260 379344
rect 273300 379400 273364 379404
rect 273300 379344 273314 379400
rect 273314 379344 273364 379400
rect 273300 379340 273364 379344
rect 275692 379400 275756 379404
rect 275692 379344 275742 379400
rect 275742 379344 275756 379400
rect 275692 379340 275756 379344
rect 285996 379400 286060 379404
rect 285996 379344 286010 379400
rect 286010 379344 286060 379400
rect 285996 379340 286060 379344
rect 288204 379340 288268 379404
rect 290964 379340 291028 379404
rect 293356 379400 293420 379404
rect 293356 379344 293370 379400
rect 293370 379344 293420 379400
rect 293356 379340 293420 379344
rect 295932 379400 295996 379404
rect 295932 379344 295946 379400
rect 295946 379344 295996 379400
rect 295932 379340 295996 379344
rect 298508 379340 298572 379404
rect 305868 379400 305932 379404
rect 305868 379344 305882 379400
rect 305882 379344 305932 379400
rect 305868 379340 305932 379344
rect 308444 379340 308508 379404
rect 311020 379400 311084 379404
rect 311020 379344 311034 379400
rect 311034 379344 311084 379400
rect 311020 379340 311084 379344
rect 318380 379340 318444 379404
rect 320956 379400 321020 379404
rect 320956 379344 320970 379400
rect 320970 379344 321020 379400
rect 320956 379340 321020 379344
rect 325924 379400 325988 379404
rect 325924 379344 325938 379400
rect 325938 379344 325988 379400
rect 325924 379340 325988 379344
rect 396028 379400 396092 379404
rect 396028 379344 396078 379400
rect 396078 379344 396092 379400
rect 396028 379340 396092 379344
rect 397132 379340 397196 379404
rect 398236 379400 398300 379404
rect 398236 379344 398250 379400
rect 398250 379344 398300 379400
rect 398236 379340 398300 379344
rect 399524 379400 399588 379404
rect 399524 379344 399538 379400
rect 399538 379344 399588 379400
rect 399524 379340 399588 379344
rect 406516 379340 406580 379404
rect 407620 379400 407684 379404
rect 407620 379344 407634 379400
rect 407634 379344 407684 379400
rect 407620 379340 407684 379344
rect 408356 379400 408420 379404
rect 408356 379344 408370 379400
rect 408370 379344 408420 379400
rect 408356 379340 408420 379344
rect 410748 379340 410812 379404
rect 411300 379400 411364 379404
rect 411300 379344 411314 379400
rect 411314 379344 411364 379400
rect 411300 379340 411364 379344
rect 412404 379400 412468 379404
rect 412404 379344 412418 379400
rect 412418 379344 412468 379400
rect 412404 379340 412468 379344
rect 420684 379400 420748 379404
rect 420684 379344 420698 379400
rect 420698 379344 420748 379400
rect 420684 379340 420748 379344
rect 428228 379400 428292 379404
rect 428228 379344 428242 379400
rect 428242 379344 428292 379400
rect 428228 379340 428292 379344
rect 431172 379400 431236 379404
rect 431172 379344 431186 379400
rect 431186 379344 431236 379400
rect 431172 379340 431236 379344
rect 434300 379400 434364 379404
rect 434300 379344 434314 379400
rect 434314 379344 434364 379400
rect 434300 379340 434364 379344
rect 437980 379400 438044 379404
rect 437980 379344 437994 379400
rect 437994 379344 438044 379400
rect 437980 379340 438044 379344
rect 451044 379400 451108 379404
rect 451044 379344 451058 379400
rect 451058 379344 451108 379400
rect 451044 379340 451108 379344
rect 453436 379340 453500 379404
rect 455828 379340 455892 379404
rect 460980 379400 461044 379404
rect 460980 379344 460994 379400
rect 460994 379344 461044 379400
rect 460980 379340 461044 379344
rect 463556 379400 463620 379404
rect 463556 379344 463570 379400
rect 463570 379344 463620 379400
rect 463556 379340 463620 379344
rect 473492 379400 473556 379404
rect 473492 379344 473506 379400
rect 473506 379344 473556 379400
rect 473492 379340 473556 379344
rect 480852 379340 480916 379404
rect 486004 379400 486068 379404
rect 486004 379344 486018 379400
rect 486018 379344 486068 379400
rect 486004 379340 486068 379344
rect 503300 379340 503364 379404
rect 78260 379204 78324 379268
rect 81756 379204 81820 379268
rect 90036 379204 90100 379268
rect 44772 379068 44836 379132
rect 93716 379204 93780 379268
rect 99420 379264 99484 379268
rect 99420 379208 99470 379264
rect 99470 379208 99484 379264
rect 99420 379204 99484 379208
rect 102916 379264 102980 379268
rect 102916 379208 102966 379264
rect 102966 379208 102980 379264
rect 102916 379204 102980 379208
rect 104020 379204 104084 379268
rect 118188 379204 118252 379268
rect 238156 379264 238220 379268
rect 238156 379208 238206 379264
rect 238206 379208 238220 379264
rect 238156 379204 238220 379208
rect 78260 378932 78324 378996
rect 274404 379204 274468 379268
rect 276060 379264 276124 379268
rect 276060 379208 276110 379264
rect 276110 379208 276124 379264
rect 276060 379204 276124 379208
rect 276980 379264 277044 379268
rect 276980 379208 277030 379264
rect 277030 379208 277044 379264
rect 276980 379204 277044 379208
rect 278452 379264 278516 379268
rect 278452 379208 278466 379264
rect 278466 379208 278516 379264
rect 278452 379204 278516 379208
rect 280844 379264 280908 379268
rect 280844 379208 280858 379264
rect 280858 379208 280908 379264
rect 280844 379204 280908 379208
rect 283420 379204 283484 379268
rect 300900 379264 300964 379268
rect 300900 379208 300914 379264
rect 300914 379208 300964 379264
rect 300900 379204 300964 379208
rect 401732 379204 401796 379268
rect 403020 379264 403084 379268
rect 403020 379208 403034 379264
rect 403034 379208 403084 379264
rect 403020 379204 403084 379208
rect 414612 379264 414676 379268
rect 414612 379208 414626 379264
rect 414626 379208 414676 379264
rect 414612 379204 414676 379208
rect 415900 379264 415964 379268
rect 415900 379208 415914 379264
rect 415914 379208 415964 379264
rect 415900 379204 415964 379208
rect 416084 379264 416148 379268
rect 416084 379208 416098 379264
rect 416098 379208 416148 379264
rect 416084 379204 416148 379208
rect 278084 379068 278148 379132
rect 343404 379128 343468 379132
rect 343404 379072 343454 379128
rect 343454 379072 343468 379128
rect 343404 379068 343468 379072
rect 400444 379068 400508 379132
rect 273484 378992 273548 378996
rect 273484 378936 273498 378992
rect 273498 378936 273548 378992
rect 273484 378932 273548 378936
rect 303476 378932 303540 378996
rect 343220 378932 343284 378996
rect 423444 379204 423508 379268
rect 419396 379128 419460 379132
rect 419396 379072 419410 379128
rect 419410 379072 419460 379128
rect 419396 379068 419460 379072
rect 465948 379068 466012 379132
rect 470916 378992 470980 378996
rect 470916 378936 470930 378992
rect 470930 378936 470980 378992
rect 79548 378796 79612 378860
rect 250668 378856 250732 378860
rect 470916 378932 470980 378936
rect 250668 378800 250682 378856
rect 250682 378800 250732 378856
rect 250668 378796 250732 378800
rect 377628 378796 377692 378860
rect 429700 378796 429764 378860
rect 468524 378796 468588 378860
rect 475884 378796 475948 378860
rect 478460 378796 478524 378860
rect 483428 378856 483492 378860
rect 483428 378800 483442 378856
rect 483442 378800 483492 378856
rect 483428 378796 483492 378800
rect 240548 378660 240612 378724
rect 377444 378660 377508 378724
rect 433380 378660 433444 378724
rect 76052 378524 76116 378588
rect 97028 378584 97092 378588
rect 97028 378528 97078 378584
rect 97078 378528 97092 378584
rect 97028 378524 97092 378528
rect 98132 378524 98196 378588
rect 101812 378584 101876 378588
rect 101812 378528 101862 378584
rect 101862 378528 101876 378584
rect 101812 378524 101876 378528
rect 107516 378584 107580 378588
rect 107516 378528 107566 378584
rect 107566 378528 107580 378584
rect 107516 378524 107580 378528
rect 119108 378524 119172 378588
rect 208348 378524 208412 378588
rect 125916 378448 125980 378452
rect 125916 378392 125966 378448
rect 125966 378392 125980 378448
rect 125916 378388 125980 378392
rect 131068 378448 131132 378452
rect 131068 378392 131082 378448
rect 131082 378392 131132 378448
rect 131068 378388 131132 378392
rect 133460 378448 133524 378452
rect 133460 378392 133510 378448
rect 133510 378392 133524 378448
rect 133460 378388 133524 378392
rect 138428 378448 138492 378452
rect 138428 378392 138478 378448
rect 138478 378392 138492 378448
rect 138428 378388 138492 378392
rect 183508 378388 183572 378452
rect 241836 378388 241900 378452
rect 253612 378388 253676 378452
rect 256004 378448 256068 378452
rect 258396 378584 258460 378588
rect 258396 378528 258410 378584
rect 258410 378528 258460 378584
rect 258396 378524 258460 378528
rect 260604 378584 260668 378588
rect 260604 378528 260618 378584
rect 260618 378528 260668 378584
rect 260604 378524 260668 378528
rect 260972 378584 261036 378588
rect 260972 378528 260986 378584
rect 260986 378528 261036 378584
rect 260972 378524 261036 378528
rect 262812 378584 262876 378588
rect 262812 378528 262826 378584
rect 262826 378528 262876 378584
rect 262812 378524 262876 378528
rect 263548 378584 263612 378588
rect 263548 378528 263598 378584
rect 263598 378528 263612 378584
rect 263548 378524 263612 378528
rect 265940 378584 266004 378588
rect 265940 378528 265954 378584
rect 265954 378528 266004 378584
rect 265940 378524 266004 378528
rect 266308 378584 266372 378588
rect 266308 378528 266358 378584
rect 266358 378528 266372 378584
rect 266308 378524 266372 378528
rect 267596 378584 267660 378588
rect 267596 378528 267610 378584
rect 267610 378528 267660 378584
rect 267596 378524 267660 378528
rect 268332 378524 268396 378588
rect 408724 378584 408788 378588
rect 408724 378528 408738 378584
rect 408738 378528 408788 378584
rect 408724 378524 408788 378528
rect 418476 378584 418540 378588
rect 418476 378528 418490 378584
rect 418490 378528 418540 378584
rect 418476 378524 418540 378528
rect 421788 378584 421852 378588
rect 421788 378528 421802 378584
rect 421802 378528 421852 378584
rect 421788 378524 421852 378528
rect 430988 378524 431052 378588
rect 436876 378524 436940 378588
rect 256004 378392 256018 378448
rect 256018 378392 256068 378448
rect 256004 378388 256068 378392
rect 100708 378312 100772 378316
rect 100708 378256 100758 378312
rect 100758 378256 100772 378312
rect 100708 378252 100772 378256
rect 183140 378252 183204 378316
rect 422892 378252 422956 378316
rect 87644 378116 87708 378180
rect 279004 378116 279068 378180
rect 410012 378176 410076 378180
rect 410012 378120 410026 378176
rect 410026 378120 410076 378176
rect 410012 378116 410076 378120
rect 417004 378176 417068 378180
rect 417004 378120 417018 378176
rect 417018 378120 417068 378176
rect 417004 378116 417068 378120
rect 418108 378176 418172 378180
rect 418108 378120 418158 378176
rect 418158 378120 418172 378176
rect 418108 378116 418172 378120
rect 423996 378176 424060 378180
rect 423996 378120 424010 378176
rect 424010 378120 424060 378176
rect 423996 378116 424060 378120
rect 425284 378116 425348 378180
rect 426388 378176 426452 378180
rect 426388 378120 426438 378176
rect 426438 378120 426452 378176
rect 426388 378116 426452 378120
rect 428596 378116 428660 378180
rect 432276 378176 432340 378180
rect 432276 378120 432290 378176
rect 432290 378120 432340 378176
rect 432276 378116 432340 378120
rect 435772 378116 435836 378180
rect 439084 378116 439148 378180
rect 458404 378116 458468 378180
rect 57100 377980 57164 378044
rect 105308 377980 105372 378044
rect 106412 377844 106476 377908
rect 211844 377980 211908 378044
rect 213316 377980 213380 378044
rect 215340 377980 215404 378044
rect 359780 377980 359844 378044
rect 372660 377844 372724 377908
rect 214236 376620 214300 376684
rect 214052 376484 214116 376548
rect 359964 375940 360028 376004
rect 217548 375668 217612 375732
rect 376708 375320 376772 375324
rect 376708 375264 376758 375320
rect 376758 375264 376772 375320
rect 376708 375260 376772 375264
rect 377812 375260 377876 375324
rect 216628 374640 216692 374644
rect 216628 374584 216678 374640
rect 216678 374584 216692 374640
rect 216628 374580 216692 374584
rect 178540 358864 178604 358868
rect 178540 358808 178590 358864
rect 178590 358808 178604 358864
rect 178540 358804 178604 358808
rect 179644 358864 179708 358868
rect 179644 358808 179694 358864
rect 179694 358808 179708 358864
rect 179644 358804 179708 358808
rect 190868 358864 190932 358868
rect 190868 358808 190918 358864
rect 190918 358808 190932 358864
rect 190868 358804 190932 358808
rect 338436 358864 338500 358868
rect 338436 358808 338486 358864
rect 338486 358808 338500 358864
rect 338436 358804 338500 358808
rect 339724 358864 339788 358868
rect 339724 358808 339774 358864
rect 339774 358808 339788 358864
rect 339724 358804 339788 358808
rect 350948 358804 351012 358868
rect 498516 358804 498580 358868
rect 499804 358804 499868 358868
rect 510844 358864 510908 358868
rect 510844 358808 510894 358864
rect 510894 358808 510908 358864
rect 510844 358804 510908 358808
rect 57468 357308 57532 357372
rect 53052 304948 53116 305012
rect 95910 273804 95974 273868
rect 130998 273728 131062 273732
rect 130998 273672 131026 273728
rect 131026 273672 131062 273728
rect 130998 273668 131062 273672
rect 145958 273728 146022 273732
rect 145958 273672 145986 273728
rect 145986 273672 146022 273728
rect 145958 273668 146022 273672
rect 440934 273728 440998 273732
rect 440934 273672 440938 273728
rect 440938 273672 440998 273728
rect 440934 273668 440998 273672
rect 133446 273592 133510 273596
rect 133446 273536 133474 273592
rect 133474 273536 133510 273592
rect 133446 273532 133510 273536
rect 135894 273592 135958 273596
rect 135894 273536 135902 273592
rect 135902 273536 135958 273592
rect 135894 273532 135958 273536
rect 138478 273592 138542 273596
rect 138478 273536 138534 273592
rect 138534 273536 138542 273592
rect 138478 273532 138542 273536
rect 140926 273532 140990 273596
rect 250742 273592 250806 273596
rect 250742 273536 250774 273592
rect 250774 273536 250806 273592
rect 250742 273532 250806 273536
rect 272230 273592 272294 273596
rect 272230 273536 272246 273592
rect 272246 273536 272294 273592
rect 272230 273532 272294 273536
rect 280934 273592 280998 273596
rect 280934 273536 280950 273592
rect 280950 273536 280998 273592
rect 280934 273532 280998 273536
rect 416046 273592 416110 273596
rect 416046 273536 416098 273592
rect 416098 273536 416110 273592
rect 416046 273532 416110 273536
rect 427606 273592 427670 273596
rect 427606 273536 427634 273592
rect 427634 273536 427670 273592
rect 427606 273532 427670 273536
rect 433318 273592 433382 273596
rect 433318 273536 433338 273592
rect 433338 273536 433382 273592
rect 433318 273532 433382 273536
rect 273300 273456 273364 273460
rect 273300 273400 273314 273456
rect 273314 273400 273364 273456
rect 273300 273396 273364 273400
rect 376892 273260 376956 273324
rect 377996 273260 378060 273324
rect 378364 273260 378428 273324
rect 430988 273320 431052 273324
rect 430988 273264 431002 273320
rect 431002 273264 431052 273320
rect 430988 273260 431052 273264
rect 77156 273184 77220 273188
rect 77156 273128 77170 273184
rect 77170 273128 77220 273184
rect 77156 273124 77220 273128
rect 88380 273184 88444 273188
rect 88380 273128 88394 273184
rect 88394 273128 88444 273184
rect 88380 273124 88444 273128
rect 90772 273184 90836 273188
rect 90772 273128 90786 273184
rect 90786 273128 90836 273184
rect 90772 273124 90836 273128
rect 93716 273184 93780 273188
rect 93716 273128 93730 273184
rect 93730 273128 93780 273184
rect 93716 273124 93780 273128
rect 98132 273184 98196 273188
rect 98132 273128 98146 273184
rect 98146 273128 98196 273184
rect 98132 273124 98196 273128
rect 101812 273124 101876 273188
rect 196756 273124 196820 273188
rect 198044 273124 198108 273188
rect 318380 273124 318444 273188
rect 486004 273124 486068 273188
rect 112116 272988 112180 273052
rect 198228 272988 198292 273052
rect 311020 272988 311084 273052
rect 483244 272988 483308 273052
rect 98500 272912 98564 272916
rect 98500 272856 98514 272912
rect 98514 272856 98564 272912
rect 95924 272776 95988 272780
rect 95924 272720 95938 272776
rect 95938 272720 95988 272776
rect 95924 272716 95988 272720
rect 98500 272852 98564 272856
rect 99420 272912 99484 272916
rect 99420 272856 99434 272912
rect 99434 272856 99484 272912
rect 99420 272852 99484 272856
rect 199332 272852 199396 272916
rect 305868 272852 305932 272916
rect 359412 272852 359476 272916
rect 423444 272912 423508 272916
rect 423444 272856 423458 272912
rect 423458 272856 423508 272912
rect 100708 272716 100772 272780
rect 199516 272716 199580 272780
rect 283420 272776 283484 272780
rect 283420 272720 283434 272776
rect 283434 272720 283484 272776
rect 118004 272580 118068 272644
rect 196572 272580 196636 272644
rect 278452 272580 278516 272644
rect 283420 272716 283484 272720
rect 288204 272776 288268 272780
rect 288204 272720 288218 272776
rect 288218 272720 288268 272776
rect 288204 272716 288268 272720
rect 290964 272776 291028 272780
rect 290964 272720 290978 272776
rect 290978 272720 291028 272776
rect 290964 272716 291028 272720
rect 295932 272776 295996 272780
rect 295932 272720 295946 272776
rect 295946 272720 295996 272776
rect 295932 272716 295996 272720
rect 377996 272716 378060 272780
rect 422892 272716 422956 272780
rect 423444 272852 423508 272856
rect 423812 272912 423876 272916
rect 423812 272856 423826 272912
rect 423826 272856 423876 272912
rect 423812 272852 423876 272856
rect 426388 272912 426452 272916
rect 426388 272856 426438 272912
rect 426438 272856 426452 272912
rect 426388 272852 426452 272856
rect 428228 272912 428292 272916
rect 428228 272856 428242 272912
rect 428242 272856 428292 272912
rect 428228 272852 428292 272856
rect 468524 272912 468588 272916
rect 468524 272856 468538 272912
rect 468538 272856 468588 272912
rect 468524 272852 468588 272856
rect 470916 272912 470980 272916
rect 470916 272856 470930 272912
rect 470930 272856 470980 272912
rect 470916 272852 470980 272856
rect 426020 272716 426084 272780
rect 478460 272776 478524 272780
rect 478460 272720 478474 272776
rect 478474 272720 478524 272776
rect 478460 272716 478524 272720
rect 480852 272776 480916 272780
rect 480852 272720 480866 272776
rect 480866 272720 480916 272776
rect 480852 272716 480916 272720
rect 285996 272580 286060 272644
rect 298508 272640 298572 272644
rect 298508 272584 298522 272640
rect 298522 272584 298572 272640
rect 298508 272580 298572 272584
rect 300900 272640 300964 272644
rect 300900 272584 300914 272640
rect 300914 272584 300964 272640
rect 300900 272580 300964 272584
rect 473492 272640 473556 272644
rect 473492 272584 473506 272640
rect 473506 272584 473556 272640
rect 473492 272580 473556 272584
rect 475884 272640 475948 272644
rect 475884 272584 475898 272640
rect 475898 272584 475948 272640
rect 475884 272580 475948 272584
rect 57468 272444 57532 272508
rect 119108 272444 119172 272508
rect 217180 272444 217244 272508
rect 293356 272444 293420 272508
rect 83044 272368 83108 272372
rect 83044 272312 83058 272368
rect 83058 272312 83108 272368
rect 83044 272308 83108 272312
rect 101812 272308 101876 272372
rect 85436 272232 85500 272236
rect 85436 272176 85450 272232
rect 85450 272176 85500 272232
rect 85436 272172 85500 272176
rect 113588 272232 113652 272236
rect 113588 272176 113602 272232
rect 113602 272176 113652 272232
rect 113588 272172 113652 272176
rect 235948 272232 236012 272236
rect 235948 272176 235998 272232
rect 235998 272176 236012 272232
rect 235948 272172 236012 272176
rect 401732 272232 401796 272236
rect 401732 272176 401746 272232
rect 401746 272176 401796 272232
rect 401732 272172 401796 272176
rect 455828 272232 455892 272236
rect 455828 272176 455842 272232
rect 455842 272176 455892 272232
rect 455828 272172 455892 272176
rect 76052 271764 76116 271828
rect 83964 271764 84028 271828
rect 88748 271764 88812 271828
rect 94452 271764 94516 271828
rect 102732 271764 102796 271828
rect 108252 271764 108316 271828
rect 125916 271764 125980 271828
rect 143580 271824 143644 271828
rect 143580 271768 143594 271824
rect 143594 271768 143644 271824
rect 143580 271764 143644 271768
rect 154068 271764 154132 271828
rect 155908 271764 155972 271828
rect 158484 271764 158548 271828
rect 213868 271764 213932 271828
rect 256188 271764 256252 271828
rect 263548 271824 263612 271828
rect 263548 271768 263598 271824
rect 263598 271768 263612 271824
rect 263548 271764 263612 271768
rect 265940 271764 266004 271828
rect 268332 271764 268396 271828
rect 270908 271764 270972 271828
rect 273484 271764 273548 271828
rect 275324 271764 275388 271828
rect 276244 271764 276308 271828
rect 276980 271764 277044 271828
rect 278084 271764 278148 271828
rect 303476 271764 303540 271828
rect 308628 271764 308692 271828
rect 404124 271764 404188 271828
rect 425284 271764 425348 271828
rect 428596 271764 428660 271828
rect 439268 271764 439332 271828
rect 448284 271764 448348 271828
rect 451044 271764 451108 271828
rect 453436 271764 453500 271828
rect 458404 271764 458468 271828
rect 460980 271824 461044 271828
rect 460980 271768 460994 271824
rect 460994 271768 461044 271824
rect 460980 271764 461044 271768
rect 80468 271628 80532 271692
rect 103836 271628 103900 271692
rect 111012 271628 111076 271692
rect 120764 271628 120828 271692
rect 123524 271628 123588 271692
rect 160876 271628 160940 271692
rect 163452 271628 163516 271692
rect 166028 271628 166092 271692
rect 198964 271628 199028 271692
rect 325556 271628 325620 271692
rect 343220 271628 343284 271692
rect 465948 271628 466012 271692
rect 101076 271492 101140 271556
rect 115980 271552 116044 271556
rect 115980 271496 115994 271552
rect 115994 271496 116044 271552
rect 115980 271492 116044 271496
rect 118372 271492 118436 271556
rect 150940 271492 151004 271556
rect 198780 271492 198844 271556
rect 315068 271492 315132 271556
rect 343404 271552 343468 271556
rect 343404 271496 343454 271552
rect 343454 271496 343468 271552
rect 343404 271492 343468 271496
rect 379468 271492 379532 271556
rect 413692 271492 413756 271556
rect 443500 271492 443564 271556
rect 503484 271492 503548 271556
rect 78260 271356 78324 271420
rect 91508 271356 91572 271420
rect 105860 271356 105924 271420
rect 183140 271356 183204 271420
rect 313412 271356 313476 271420
rect 377260 271356 377324 271420
rect 408172 271356 408236 271420
rect 418476 271356 418540 271420
rect 435956 271356 436020 271420
rect 445892 271356 445956 271420
rect 503116 271356 503180 271420
rect 81940 271220 82004 271284
rect 107516 271220 107580 271284
rect 258396 271220 258460 271284
rect 260972 271220 261036 271284
rect 279004 271220 279068 271284
rect 397132 271220 397196 271284
rect 47716 271084 47780 271148
rect 109540 271084 109604 271148
rect 128676 271084 128740 271148
rect 183508 271144 183572 271148
rect 183508 271088 183522 271144
rect 183522 271088 183572 271144
rect 183508 271084 183572 271088
rect 239260 271084 239324 271148
rect 248276 271084 248340 271148
rect 253612 271084 253676 271148
rect 262076 271084 262140 271148
rect 266308 271144 266372 271148
rect 266308 271088 266358 271144
rect 266358 271088 266372 271144
rect 266308 271084 266372 271088
rect 268700 271084 268764 271148
rect 271276 271084 271340 271148
rect 417004 271220 417068 271284
rect 433564 271220 433628 271284
rect 438532 271220 438596 271284
rect 421052 271084 421116 271148
rect 79548 270948 79612 271012
rect 105308 270948 105372 271012
rect 320956 270948 321020 271012
rect 410748 270948 410812 271012
rect 429700 270948 429764 271012
rect 438348 270948 438412 271012
rect 97028 270812 97092 270876
rect 116900 270812 116964 270876
rect 148548 270812 148612 270876
rect 253428 270812 253492 270876
rect 265756 270812 265820 270876
rect 462636 270812 462700 270876
rect 86540 270676 86604 270740
rect 90036 270676 90100 270740
rect 93348 270676 93412 270740
rect 245332 270676 245396 270740
rect 252324 270676 252388 270740
rect 260604 270676 260668 270740
rect 267596 270676 267660 270740
rect 411300 270736 411364 270740
rect 411300 270680 411350 270736
rect 411350 270680 411364 270736
rect 411300 270676 411364 270680
rect 432276 270676 432340 270740
rect 87644 270540 87708 270604
rect 91324 270540 91388 270604
rect 104020 270540 104084 270604
rect 106412 270600 106476 270604
rect 106412 270544 106426 270600
rect 106426 270544 106476 270600
rect 106412 270540 106476 270544
rect 108620 270540 108684 270604
rect 111196 270540 111260 270604
rect 113220 270600 113284 270604
rect 113220 270544 113234 270600
rect 113234 270544 113284 270600
rect 113220 270540 113284 270544
rect 114508 270600 114572 270604
rect 114508 270544 114522 270600
rect 114522 270544 114572 270600
rect 114508 270540 114572 270544
rect 115796 270600 115860 270604
rect 115796 270544 115846 270600
rect 115846 270544 115860 270600
rect 115796 270540 115860 270544
rect 237052 270540 237116 270604
rect 238156 270540 238220 270604
rect 242940 270600 243004 270604
rect 242940 270544 242954 270600
rect 242954 270544 243004 270600
rect 242940 270540 243004 270544
rect 244228 270540 244292 270604
rect 246436 270540 246500 270604
rect 247724 270540 247788 270604
rect 248644 270540 248708 270604
rect 250116 270540 250180 270604
rect 251220 270600 251284 270604
rect 251220 270544 251234 270600
rect 251234 270544 251284 270600
rect 251220 270540 251284 270544
rect 254532 270540 254596 270604
rect 255820 270540 255884 270604
rect 256924 270540 256988 270604
rect 258396 270540 258460 270604
rect 259500 270600 259564 270604
rect 259500 270544 259514 270600
rect 259514 270544 259564 270600
rect 259500 270540 259564 270544
rect 262812 270540 262876 270604
rect 263916 270540 263980 270604
rect 269804 270540 269868 270604
rect 274404 270540 274468 270604
rect 396028 270600 396092 270604
rect 396028 270544 396078 270600
rect 396078 270544 396092 270600
rect 396028 270540 396092 270544
rect 397500 270600 397564 270604
rect 397500 270544 397514 270600
rect 397514 270544 397564 270600
rect 397500 270540 397564 270544
rect 399524 270540 399588 270604
rect 400444 270540 400508 270604
rect 403020 270600 403084 270604
rect 403020 270544 403034 270600
rect 403034 270544 403084 270600
rect 403020 270540 403084 270544
rect 405044 270540 405108 270604
rect 406516 270540 406580 270604
rect 407620 270540 407684 270604
rect 408724 270540 408788 270604
rect 410012 270540 410076 270604
rect 412404 270540 412468 270604
rect 413324 270540 413388 270604
rect 414428 270540 414492 270604
rect 415532 270540 415596 270604
rect 418292 270540 418356 270604
rect 419212 270540 419276 270604
rect 420684 270540 420748 270604
rect 421788 270540 421852 270604
rect 436876 270540 436940 270604
rect 323348 270404 323412 270468
rect 435772 270404 435836 270468
rect 241652 270268 241716 270332
rect 240548 270132 240612 270196
rect 217364 270056 217428 270060
rect 217364 270000 217378 270056
rect 217378 270000 217428 270056
rect 217364 269996 217428 270000
rect 434668 269860 434732 269924
rect 431172 269724 431236 269788
rect 217548 268364 217612 268428
rect 54340 253948 54404 254012
rect 339724 253404 339788 253468
rect 179644 253268 179708 253332
rect 499804 253268 499868 253332
rect 178540 253132 178604 253196
rect 350948 253132 351012 253196
rect 338436 252996 338500 253060
rect 498516 252724 498580 252788
rect 190868 252588 190932 252652
rect 510844 252648 510908 252652
rect 510844 252592 510894 252648
rect 510894 252592 510908 252648
rect 510844 252588 510908 252592
rect 57468 252452 57532 252516
rect 216628 252452 216692 252516
rect 217364 252452 217428 252516
rect 217548 251772 217612 251836
rect 377996 251772 378060 251836
rect 44956 251092 45020 251156
rect 44036 250956 44100 251020
rect 51580 201452 51644 201516
rect 219940 167044 220004 167108
rect 57652 166908 57716 166972
rect 148364 166908 148428 166972
rect 206324 166908 206388 166972
rect 57836 166772 57900 166836
rect 98500 166696 98564 166700
rect 98500 166640 98514 166696
rect 98514 166640 98564 166696
rect 98500 166636 98564 166640
rect 101076 166696 101140 166700
rect 101076 166640 101090 166696
rect 101090 166640 101140 166696
rect 101076 166636 101140 166640
rect 105860 166696 105924 166700
rect 105860 166640 105874 166696
rect 105874 166640 105924 166696
rect 105860 166636 105924 166640
rect 108252 166696 108316 166700
rect 108252 166640 108266 166696
rect 108266 166640 108316 166696
rect 108252 166636 108316 166640
rect 138478 166832 138542 166836
rect 138478 166776 138534 166832
rect 138534 166776 138542 166832
rect 138478 166772 138542 166776
rect 143510 166832 143574 166836
rect 143510 166776 143538 166832
rect 143538 166776 143574 166832
rect 143510 166772 143574 166776
rect 145958 166832 146022 166836
rect 145958 166776 145986 166832
rect 145986 166776 146022 166832
rect 145958 166772 146022 166776
rect 210556 166772 210620 166836
rect 140926 166636 140990 166700
rect 163366 166696 163430 166700
rect 163366 166640 163374 166696
rect 163374 166640 163430 166696
rect 163366 166636 163430 166640
rect 165950 166636 166014 166700
rect 208164 166636 208228 166700
rect 113318 166560 113382 166564
rect 113318 166504 113326 166560
rect 113326 166504 113382 166560
rect 113318 166500 113382 166504
rect 150940 166560 151004 166564
rect 150940 166504 150954 166560
rect 150954 166504 151004 166560
rect 150940 166500 151004 166504
rect 153332 166560 153396 166564
rect 153332 166504 153346 166560
rect 153346 166504 153396 166560
rect 153332 166500 153396 166504
rect 253612 166560 253676 166564
rect 253612 166504 253626 166560
rect 253626 166504 253676 166560
rect 253612 166500 253676 166504
rect 265940 166560 266004 166564
rect 265940 166504 265954 166560
rect 265954 166504 266004 166560
rect 265940 166500 266004 166504
rect 270908 166560 270972 166564
rect 270908 166504 270922 166560
rect 270922 166504 270972 166560
rect 270908 166500 270972 166504
rect 288278 166696 288342 166700
rect 288278 166640 288310 166696
rect 288310 166640 288342 166696
rect 288278 166636 288342 166640
rect 295894 166696 295958 166700
rect 298478 166832 298542 166836
rect 298478 166776 298522 166832
rect 298522 166776 298542 166832
rect 298478 166772 298542 166776
rect 303510 166832 303574 166836
rect 303510 166776 303526 166832
rect 303526 166776 303574 166832
rect 303510 166772 303574 166776
rect 313438 166772 313502 166836
rect 416046 166832 416110 166836
rect 416046 166776 416098 166832
rect 416098 166776 416110 166832
rect 416046 166772 416110 166776
rect 418476 166832 418540 166836
rect 418476 166776 418490 166832
rect 418490 166776 418540 166832
rect 418476 166772 418540 166776
rect 423444 166832 423508 166836
rect 423444 166776 423458 166832
rect 423458 166776 423508 166832
rect 423444 166772 423508 166776
rect 426020 166832 426084 166836
rect 426020 166776 426034 166832
rect 426034 166776 426084 166832
rect 426020 166772 426084 166776
rect 470990 166832 471054 166836
rect 470990 166776 471022 166832
rect 471022 166776 471054 166832
rect 470990 166772 471054 166776
rect 473438 166832 473502 166836
rect 473438 166776 473450 166832
rect 473450 166776 473502 166832
rect 473438 166772 473502 166776
rect 475886 166832 475950 166836
rect 475886 166776 475898 166832
rect 475898 166776 475950 166832
rect 475886 166772 475950 166776
rect 478470 166832 478534 166836
rect 478470 166776 478474 166832
rect 478474 166776 478534 166832
rect 478470 166772 478534 166776
rect 480918 166832 480982 166836
rect 480918 166776 480958 166832
rect 480958 166776 480982 166832
rect 480918 166772 480982 166776
rect 295894 166640 295946 166696
rect 295946 166640 295958 166696
rect 295894 166636 295958 166640
rect 305958 166636 306022 166700
rect 308542 166696 308606 166700
rect 308542 166640 308550 166696
rect 308550 166640 308606 166696
rect 308542 166636 308606 166640
rect 315886 166696 315950 166700
rect 315886 166640 315910 166696
rect 315910 166640 315950 166696
rect 315886 166636 315950 166640
rect 483366 166696 483430 166700
rect 483366 166640 483386 166696
rect 483386 166640 483430 166696
rect 483366 166636 483430 166640
rect 485950 166696 486014 166700
rect 485950 166640 485962 166696
rect 485962 166640 486014 166696
rect 485950 166636 486014 166640
rect 290998 166500 291062 166564
rect 413598 166560 413662 166564
rect 413598 166504 413614 166560
rect 413614 166504 413662 166560
rect 413598 166500 413662 166504
rect 503222 166560 503286 166564
rect 503222 166504 503258 166560
rect 503258 166504 503286 166560
rect 503222 166500 503286 166504
rect 96108 166288 96172 166292
rect 96108 166232 96122 166288
rect 96122 166232 96172 166288
rect 96108 166228 96172 166232
rect 408172 166288 408236 166292
rect 408172 166232 408186 166288
rect 408186 166232 408236 166288
rect 408172 166228 408236 166232
rect 428228 166288 428292 166292
rect 428228 166232 428242 166288
rect 428242 166232 428292 166288
rect 428228 166228 428292 166232
rect 81756 165548 81820 165612
rect 85436 165548 85500 165612
rect 90772 165548 90836 165612
rect 92428 165548 92492 165612
rect 95740 165548 95804 165612
rect 99420 165608 99484 165612
rect 99420 165552 99434 165608
rect 99434 165552 99484 165608
rect 99420 165548 99484 165552
rect 103468 165608 103532 165612
rect 103468 165552 103518 165608
rect 103518 165552 103532 165608
rect 103468 165548 103532 165552
rect 109724 165608 109788 165612
rect 109724 165552 109738 165608
rect 109738 165552 109788 165608
rect 109724 165548 109788 165552
rect 111012 165548 111076 165612
rect 111196 165608 111260 165612
rect 111196 165552 111210 165608
rect 111210 165552 111260 165608
rect 111196 165548 111260 165552
rect 112116 165548 112180 165612
rect 113588 165608 113652 165612
rect 113588 165552 113602 165608
rect 113602 165552 113652 165608
rect 113588 165548 113652 165552
rect 115980 165608 116044 165612
rect 115980 165552 115994 165608
rect 115994 165552 116044 165608
rect 115980 165548 116044 165552
rect 116900 165548 116964 165612
rect 118004 165548 118068 165612
rect 118372 165608 118436 165612
rect 118372 165552 118386 165608
rect 118386 165552 118436 165608
rect 118372 165548 118436 165552
rect 120948 165608 121012 165612
rect 120948 165552 120962 165608
rect 120962 165552 121012 165608
rect 120948 165548 121012 165552
rect 123524 165608 123588 165612
rect 123524 165552 123538 165608
rect 123538 165552 123588 165608
rect 123524 165548 123588 165552
rect 125916 165608 125980 165612
rect 125916 165552 125930 165608
rect 125930 165552 125980 165608
rect 125916 165548 125980 165552
rect 128492 165548 128556 165612
rect 130884 165548 130948 165612
rect 133460 165548 133524 165612
rect 183140 165608 183204 165612
rect 183140 165552 183190 165608
rect 183190 165552 183204 165608
rect 183140 165548 183204 165552
rect 236132 165608 236196 165612
rect 236132 165552 236146 165608
rect 236146 165552 236196 165608
rect 236132 165548 236196 165552
rect 239628 165548 239692 165612
rect 243124 165548 243188 165612
rect 247540 165548 247604 165612
rect 258028 165548 258092 165612
rect 261708 165548 261772 165612
rect 273484 165608 273548 165612
rect 273484 165552 273498 165608
rect 273498 165552 273548 165608
rect 273484 165548 273548 165552
rect 276060 165608 276124 165612
rect 276060 165552 276074 165608
rect 276074 165552 276124 165608
rect 276060 165548 276124 165552
rect 278452 165608 278516 165612
rect 278452 165552 278466 165608
rect 278466 165552 278516 165608
rect 278452 165548 278516 165552
rect 280844 165608 280908 165612
rect 280844 165552 280858 165608
rect 280858 165552 280908 165608
rect 280844 165548 280908 165552
rect 285996 165608 286060 165612
rect 285996 165552 286010 165608
rect 286010 165552 286060 165608
rect 285996 165548 286060 165552
rect 293356 165608 293420 165612
rect 293356 165552 293370 165608
rect 293370 165552 293420 165608
rect 293356 165548 293420 165552
rect 300900 165608 300964 165612
rect 300900 165552 300914 165608
rect 300914 165552 300964 165608
rect 300900 165548 300964 165552
rect 311020 165608 311084 165612
rect 311020 165552 311034 165608
rect 311034 165552 311084 165608
rect 311020 165548 311084 165552
rect 325924 165608 325988 165612
rect 325924 165552 325938 165608
rect 325938 165552 325988 165608
rect 325924 165548 325988 165552
rect 343220 165608 343284 165612
rect 343220 165552 343270 165608
rect 343270 165552 343284 165608
rect 343220 165548 343284 165552
rect 398236 165548 398300 165612
rect 401732 165548 401796 165612
rect 405412 165548 405476 165612
rect 410748 165548 410812 165612
rect 415900 165548 415964 165612
rect 417004 165548 417068 165612
rect 419396 165548 419460 165612
rect 423812 165608 423876 165612
rect 423812 165552 423826 165608
rect 423826 165552 423876 165608
rect 423812 165548 423876 165552
rect 427492 165548 427556 165612
rect 433380 165548 433444 165612
rect 435956 165548 436020 165612
rect 437980 165548 438044 165612
rect 440924 165548 440988 165612
rect 443500 165548 443564 165612
rect 448284 165548 448348 165612
rect 451044 165548 451108 165612
rect 453436 165548 453500 165612
rect 455828 165548 455892 165612
rect 458404 165608 458468 165612
rect 458404 165552 458418 165608
rect 458418 165552 458468 165608
rect 458404 165548 458468 165552
rect 155908 165412 155972 165476
rect 318380 165412 318444 165476
rect 468524 165412 468588 165476
rect 158484 165276 158548 165340
rect 216260 165276 216324 165340
rect 283420 165276 283484 165340
rect 465948 165276 466012 165340
rect 135852 165140 135916 165204
rect 200804 165140 200868 165204
rect 260972 165140 261036 165204
rect 263732 165140 263796 165204
rect 265388 165140 265452 165204
rect 272196 165140 272260 165204
rect 275692 165140 275756 165204
rect 279188 165140 279252 165204
rect 378916 165140 378980 165204
rect 463556 165140 463620 165204
rect 47900 165004 47964 165068
rect 93716 165004 93780 165068
rect 119108 165004 119172 165068
rect 183508 165064 183572 165068
rect 183508 165008 183522 165064
rect 183522 165008 183572 165064
rect 183508 165004 183572 165008
rect 268332 165004 268396 165068
rect 438532 165004 438596 165068
rect 445892 165004 445956 165068
rect 105308 164868 105372 164932
rect 106412 164868 106476 164932
rect 114508 164928 114572 164932
rect 114508 164872 114522 164928
rect 114522 164872 114572 164928
rect 114508 164868 114572 164872
rect 248276 164868 248340 164932
rect 250668 164868 250732 164932
rect 256188 164868 256252 164932
rect 258396 164868 258460 164932
rect 343404 164868 343468 164932
rect 421052 164868 421116 164932
rect 433564 164868 433628 164932
rect 88380 164792 88444 164796
rect 88380 164736 88394 164792
rect 88394 164736 88444 164792
rect 88380 164732 88444 164736
rect 107516 164732 107580 164796
rect 202460 164732 202524 164796
rect 323348 164732 323412 164796
rect 460980 164732 461044 164796
rect 160876 164596 160940 164660
rect 434668 164596 434732 164660
rect 503300 164596 503364 164660
rect 100708 164520 100772 164524
rect 100708 164464 100758 164520
rect 100758 164464 100772 164520
rect 100708 164460 100772 164464
rect 108620 164460 108684 164524
rect 115796 164460 115860 164524
rect 77156 164324 77220 164388
rect 244412 164384 244476 164388
rect 244412 164328 244426 164384
rect 244426 164328 244476 164384
rect 244412 164324 244476 164328
rect 252324 164324 252388 164388
rect 256924 164324 256988 164388
rect 260604 164324 260668 164388
rect 267596 164324 267660 164388
rect 274404 164324 274468 164388
rect 397132 164324 397196 164388
rect 404124 164324 404188 164388
rect 412404 164324 412468 164388
rect 429700 164324 429764 164388
rect 431172 164324 431236 164388
rect 57468 164188 57532 164252
rect 76052 164188 76116 164252
rect 78260 164188 78324 164252
rect 79548 164188 79612 164252
rect 80468 164188 80532 164252
rect 83044 164188 83108 164252
rect 84148 164248 84212 164252
rect 84148 164192 84198 164248
rect 84198 164192 84212 164248
rect 84148 164188 84212 164192
rect 86540 164188 86604 164252
rect 87644 164188 87708 164252
rect 88748 164188 88812 164252
rect 90036 164188 90100 164252
rect 91324 164188 91388 164252
rect 93348 164188 93412 164252
rect 94452 164188 94516 164252
rect 97028 164188 97092 164252
rect 98132 164188 98196 164252
rect 101812 164188 101876 164252
rect 102732 164188 102796 164252
rect 103836 164188 103900 164252
rect 237052 164188 237116 164252
rect 238156 164188 238220 164252
rect 240548 164188 240612 164252
rect 241652 164188 241716 164252
rect 245332 164188 245396 164252
rect 246436 164188 246500 164252
rect 248644 164188 248708 164252
rect 250116 164188 250180 164252
rect 251220 164248 251284 164252
rect 251220 164192 251234 164248
rect 251234 164192 251284 164248
rect 251220 164188 251284 164192
rect 253428 164188 253492 164252
rect 254532 164188 254596 164252
rect 255820 164188 255884 164252
rect 259500 164248 259564 164252
rect 259500 164192 259514 164248
rect 259514 164192 259564 164248
rect 259500 164188 259564 164192
rect 262812 164188 262876 164252
rect 263916 164188 263980 164252
rect 266308 164188 266372 164252
rect 268700 164188 268764 164252
rect 269804 164188 269868 164252
rect 271276 164188 271340 164252
rect 273300 164188 273364 164252
rect 276980 164188 277044 164252
rect 278084 164188 278148 164252
rect 396028 164248 396092 164252
rect 396028 164192 396078 164248
rect 396078 164192 396092 164248
rect 396028 164188 396092 164192
rect 399524 164188 399588 164252
rect 400444 164188 400508 164252
rect 403020 164248 403084 164252
rect 403020 164192 403070 164248
rect 403070 164192 403084 164248
rect 403020 164188 403084 164192
rect 406516 164188 406580 164252
rect 407620 164188 407684 164252
rect 408724 164188 408788 164252
rect 410012 164248 410076 164252
rect 410012 164192 410026 164248
rect 410026 164192 410076 164248
rect 410012 164188 410076 164192
rect 411300 164248 411364 164252
rect 411300 164192 411314 164248
rect 411314 164192 411364 164248
rect 411300 164188 411364 164192
rect 413508 164188 413572 164252
rect 414612 164188 414676 164252
rect 418292 164248 418356 164252
rect 418292 164192 418306 164248
rect 418306 164192 418356 164248
rect 418292 164188 418356 164192
rect 420684 164188 420748 164252
rect 421788 164188 421852 164252
rect 422892 164188 422956 164252
rect 425284 164188 425348 164252
rect 426388 164188 426452 164252
rect 428780 164188 428844 164252
rect 430988 164188 431052 164252
rect 432276 164188 432340 164252
rect 435772 164188 435836 164252
rect 436876 164188 436940 164252
rect 439268 164188 439332 164252
rect 203012 164052 203076 164116
rect 205036 163916 205100 163980
rect 320956 163916 321020 163980
rect 217364 163508 217428 163572
rect 57836 163236 57900 163300
rect 377260 163024 377324 163028
rect 377260 162968 377310 163024
rect 377310 162968 377324 163024
rect 377260 162964 377324 162968
rect 217548 162692 217612 162756
rect 217548 162556 217612 162620
rect 377996 162616 378060 162620
rect 377996 162560 378046 162616
rect 378046 162560 378060 162616
rect 377996 162556 378060 162560
rect 370636 149092 370700 149156
rect 217364 148276 217428 148340
rect 379468 146236 379532 146300
rect 510844 146100 510908 146164
rect 57652 145828 57716 145892
rect 190868 145420 190932 145484
rect 178540 144876 178604 144940
rect 179644 144936 179708 144940
rect 179644 144880 179694 144936
rect 179694 144880 179708 144936
rect 179644 144876 179708 144880
rect 217180 144876 217244 144940
rect 338436 144936 338500 144940
rect 338436 144880 338486 144936
rect 338486 144880 338500 144936
rect 338436 144876 338500 144880
rect 339724 144876 339788 144940
rect 350948 144876 351012 144940
rect 498516 144876 498580 144940
rect 499804 144936 499868 144940
rect 499804 144880 499854 144936
rect 499854 144880 499868 144936
rect 499804 144876 499868 144880
rect 377812 144060 377876 144124
rect 57468 140796 57532 140860
rect 207980 69940 208044 70004
rect 46796 67764 46860 67828
rect 378180 60556 378244 60620
rect 77142 59800 77206 59804
rect 77142 59744 77170 59800
rect 77170 59744 77206 59800
rect 77142 59740 77206 59744
rect 83126 59800 83190 59804
rect 83126 59744 83150 59800
rect 83150 59744 83190 59800
rect 83126 59740 83190 59744
rect 84214 59800 84278 59804
rect 84214 59744 84254 59800
rect 84254 59744 84278 59800
rect 84214 59740 84278 59744
rect 99446 59800 99510 59804
rect 99446 59744 99470 59800
rect 99470 59744 99510 59800
rect 99446 59740 99510 59744
rect 102846 59740 102910 59804
rect 107606 59800 107670 59804
rect 107606 59744 107622 59800
rect 107622 59744 107670 59800
rect 107606 59740 107670 59744
rect 255910 59800 255974 59804
rect 255910 59744 255926 59800
rect 255926 59744 255974 59800
rect 255910 59740 255974 59744
rect 260670 59800 260734 59804
rect 260670 59744 260710 59800
rect 260710 59744 260734 59800
rect 260670 59740 260734 59744
rect 261758 59800 261822 59804
rect 261758 59744 261814 59800
rect 261814 59744 261822 59800
rect 261758 59740 261822 59744
rect 262846 59800 262910 59804
rect 262846 59744 262862 59800
rect 262862 59744 262910 59800
rect 262846 59740 262910 59744
rect 263934 59740 263998 59804
rect 396054 59800 396118 59804
rect 396054 59744 396078 59800
rect 396078 59744 396118 59800
rect 396054 59740 396118 59744
rect 397142 59800 397206 59804
rect 397142 59744 397146 59800
rect 397146 59744 397206 59800
rect 397142 59740 397206 59744
rect 403126 59740 403190 59804
rect 413598 59800 413662 59804
rect 413598 59744 413614 59800
rect 413614 59744 413662 59800
rect 413598 59740 413662 59744
rect 415910 59800 415974 59804
rect 415910 59744 415914 59800
rect 415914 59744 415974 59800
rect 415910 59740 415974 59744
rect 419446 59800 419510 59804
rect 419446 59744 419502 59800
rect 419502 59744 419510 59800
rect 419446 59740 419510 59744
rect 100708 59664 100772 59668
rect 100708 59608 100758 59664
rect 100758 59608 100772 59664
rect 100708 59604 100772 59608
rect 103934 59664 103998 59668
rect 103934 59608 103942 59664
rect 103942 59608 103998 59664
rect 103934 59604 103998 59608
rect 114406 59664 114470 59668
rect 114406 59608 114430 59664
rect 114430 59608 114470 59664
rect 114406 59604 114470 59608
rect 143510 59664 143574 59668
rect 143510 59608 143538 59664
rect 143538 59608 143574 59664
rect 143510 59604 143574 59608
rect 256998 59664 257062 59668
rect 256998 59608 257030 59664
rect 257030 59608 257062 59664
rect 256998 59604 257062 59608
rect 258494 59604 258558 59668
rect 308542 59664 308606 59668
rect 308542 59608 308550 59664
rect 308550 59608 308606 59664
rect 308542 59604 308606 59608
rect 423526 59664 423590 59668
rect 423526 59608 423550 59664
rect 423550 59608 423590 59664
rect 423526 59604 423590 59608
rect 503222 59664 503286 59668
rect 503222 59608 503258 59664
rect 503258 59608 503286 59664
rect 503222 59604 503286 59608
rect 219020 59528 219084 59532
rect 219020 59472 219070 59528
rect 219070 59472 219084 59528
rect 219020 59468 219084 59472
rect 85436 59392 85500 59396
rect 85436 59336 85450 59392
rect 85450 59336 85500 59392
rect 85436 59332 85500 59336
rect 95924 59392 95988 59396
rect 95924 59336 95938 59392
rect 95938 59336 95988 59392
rect 95924 59332 95988 59336
rect 98132 59392 98196 59396
rect 98132 59336 98146 59392
rect 98146 59336 98196 59392
rect 98132 59332 98196 59336
rect 105308 59392 105372 59396
rect 105308 59336 105322 59392
rect 105322 59336 105372 59392
rect 105308 59332 105372 59336
rect 106412 59392 106476 59396
rect 106412 59336 106426 59392
rect 106426 59336 106476 59392
rect 106412 59332 106476 59336
rect 200620 59332 200684 59396
rect 259500 59392 259564 59396
rect 259500 59336 259514 59392
rect 259514 59336 259564 59392
rect 259500 59332 259564 59336
rect 398236 59392 398300 59396
rect 398236 59336 398250 59392
rect 398250 59336 398300 59392
rect 398236 59332 398300 59336
rect 410748 59392 410812 59396
rect 410748 59336 410762 59392
rect 410762 59336 410812 59392
rect 410748 59332 410812 59336
rect 417004 59392 417068 59396
rect 417004 59336 417018 59392
rect 417018 59336 417068 59392
rect 417004 59332 417068 59336
rect 418108 59392 418172 59396
rect 418108 59336 418158 59392
rect 418158 59336 418172 59392
rect 418108 59332 418172 59336
rect 421052 59392 421116 59396
rect 421052 59336 421066 59392
rect 421066 59336 421116 59392
rect 421052 59332 421116 59336
rect 421788 59392 421852 59396
rect 421788 59336 421802 59392
rect 421802 59336 421852 59392
rect 421788 59332 421852 59336
rect 425284 59392 425348 59396
rect 425284 59336 425298 59392
rect 425298 59336 425348 59392
rect 425284 59332 425348 59336
rect 426020 59392 426084 59396
rect 426020 59336 426034 59392
rect 426034 59336 426084 59392
rect 426020 59332 426084 59336
rect 428228 59392 428292 59396
rect 428228 59336 428242 59392
rect 428242 59336 428292 59392
rect 428228 59332 428292 59336
rect 468524 59392 468588 59396
rect 468524 59336 468538 59392
rect 468538 59336 468588 59392
rect 468524 59332 468588 59336
rect 54708 59196 54772 59260
rect 140820 59196 140884 59260
rect 148548 59256 148612 59260
rect 148548 59200 148562 59256
rect 148562 59200 148612 59256
rect 148548 59196 148612 59200
rect 150940 59256 151004 59260
rect 150940 59200 150954 59256
rect 150954 59200 151004 59256
rect 150940 59196 151004 59200
rect 205220 59196 205284 59260
rect 290964 59196 291028 59260
rect 295932 59256 295996 59260
rect 295932 59200 295946 59256
rect 295946 59200 295996 59256
rect 295932 59196 295996 59200
rect 298508 59256 298572 59260
rect 298508 59200 298522 59256
rect 298522 59200 298572 59256
rect 298508 59196 298572 59200
rect 303476 59256 303540 59260
rect 303476 59200 303490 59256
rect 303490 59200 303540 59256
rect 303476 59196 303540 59200
rect 357940 59196 358004 59260
rect 478460 59196 478524 59260
rect 53420 59060 53484 59124
rect 135852 59060 135916 59124
rect 138428 59120 138492 59124
rect 138428 59064 138442 59120
rect 138442 59064 138492 59120
rect 138428 59060 138492 59064
rect 206692 59060 206756 59124
rect 283420 59060 283484 59124
rect 371924 59060 371988 59124
rect 486004 59060 486068 59124
rect 59124 58924 59188 58988
rect 125916 58924 125980 58988
rect 201356 58924 201420 58988
rect 278452 58924 278516 58988
rect 374500 58924 374564 58988
rect 473492 58924 473556 58988
rect 48084 58788 48148 58852
rect 111012 58788 111076 58852
rect 202644 58788 202708 58852
rect 276060 58788 276124 58852
rect 367876 58788 367940 58852
rect 458404 58788 458468 58852
rect 46612 58652 46676 58716
rect 108252 58652 108316 58716
rect 202092 58652 202156 58716
rect 250668 58652 250732 58716
rect 375972 58652 376036 58716
rect 463556 58652 463620 58716
rect 59860 58516 59924 58580
rect 115980 58516 116044 58580
rect 219204 58516 219268 58580
rect 265204 58516 265268 58580
rect 367692 58516 367756 58580
rect 453436 58516 453500 58580
rect 59308 58380 59372 58444
rect 101076 58380 101140 58444
rect 217548 58380 217612 58444
rect 257844 58380 257908 58444
rect 377996 58380 378060 58444
rect 420684 58380 420748 58444
rect 217180 58244 217244 58308
rect 92244 58108 92308 58172
rect 113588 58108 113652 58172
rect 128308 58108 128372 58172
rect 153332 58108 153396 58172
rect 236132 58108 236196 58172
rect 272196 58108 272260 58172
rect 275692 58108 275756 58172
rect 300900 58108 300964 58172
rect 315804 58108 315868 58172
rect 325924 58108 325988 58172
rect 401732 58108 401796 58172
rect 455828 58108 455892 58172
rect 76052 57896 76116 57900
rect 76052 57840 76066 57896
rect 76066 57840 76116 57896
rect 76052 57836 76116 57840
rect 78260 57896 78324 57900
rect 78260 57840 78274 57896
rect 78274 57840 78324 57896
rect 78260 57836 78324 57840
rect 79548 57836 79612 57900
rect 80468 57896 80532 57900
rect 80468 57840 80482 57896
rect 80482 57840 80532 57896
rect 80468 57836 80532 57840
rect 81940 57836 82004 57900
rect 86540 57896 86604 57900
rect 86540 57840 86554 57896
rect 86554 57840 86604 57896
rect 86540 57836 86604 57840
rect 87644 57836 87708 57900
rect 88748 57836 88812 57900
rect 90036 57896 90100 57900
rect 90036 57840 90050 57896
rect 90050 57840 90100 57896
rect 90036 57836 90100 57840
rect 90772 57896 90836 57900
rect 90772 57840 90786 57896
rect 90786 57840 90836 57896
rect 90772 57836 90836 57840
rect 91324 57836 91388 57900
rect 93348 57836 93412 57900
rect 93716 57896 93780 57900
rect 93716 57840 93730 57896
rect 93730 57840 93780 57896
rect 93716 57836 93780 57840
rect 94452 57896 94516 57900
rect 94452 57840 94466 57896
rect 94466 57840 94516 57896
rect 94452 57836 94516 57840
rect 98500 57896 98564 57900
rect 98500 57840 98514 57896
rect 98514 57840 98564 57896
rect 98500 57836 98564 57840
rect 101812 57896 101876 57900
rect 101812 57840 101826 57896
rect 101826 57840 101876 57896
rect 101812 57836 101876 57840
rect 108620 57896 108684 57900
rect 108620 57840 108634 57896
rect 108634 57840 108684 57896
rect 108620 57836 108684 57840
rect 109540 57896 109604 57900
rect 109540 57840 109554 57896
rect 109554 57840 109604 57896
rect 109540 57836 109604 57840
rect 111196 57896 111260 57900
rect 111196 57840 111210 57896
rect 111210 57840 111260 57896
rect 111196 57836 111260 57840
rect 116900 57836 116964 57900
rect 118004 57896 118068 57900
rect 118004 57840 118018 57896
rect 118018 57840 118068 57896
rect 118004 57836 118068 57840
rect 120764 57896 120828 57900
rect 120764 57840 120778 57896
rect 120778 57840 120828 57896
rect 120764 57836 120828 57840
rect 123524 57896 123588 57900
rect 123524 57840 123538 57896
rect 123538 57840 123588 57896
rect 123524 57836 123588 57840
rect 55076 57700 55140 57764
rect 130884 57896 130948 57900
rect 130884 57840 130898 57896
rect 130898 57840 130948 57896
rect 130884 57836 130948 57840
rect 145604 57896 145668 57900
rect 145604 57840 145618 57896
rect 145618 57840 145668 57896
rect 145604 57836 145668 57840
rect 183508 57896 183572 57900
rect 183508 57840 183522 57896
rect 183522 57840 183572 57896
rect 183508 57836 183572 57840
rect 238156 57896 238220 57900
rect 238156 57840 238170 57896
rect 238170 57840 238220 57896
rect 238156 57836 238220 57840
rect 239260 57836 239324 57900
rect 240548 57896 240612 57900
rect 240548 57840 240562 57896
rect 240562 57840 240612 57896
rect 240548 57836 240612 57840
rect 241652 57836 241716 57900
rect 242940 57896 243004 57900
rect 242940 57840 242954 57896
rect 242954 57840 243004 57896
rect 242940 57836 243004 57840
rect 244228 57836 244292 57900
rect 245332 57896 245396 57900
rect 245332 57840 245346 57896
rect 245346 57840 245396 57896
rect 245332 57836 245396 57840
rect 246436 57836 246500 57900
rect 247724 57896 247788 57900
rect 247724 57840 247738 57896
rect 247738 57840 247788 57896
rect 247724 57836 247788 57840
rect 248276 57836 248340 57900
rect 248644 57836 248708 57900
rect 250116 57836 250180 57900
rect 251220 57896 251284 57900
rect 251220 57840 251234 57896
rect 251234 57840 251284 57896
rect 251220 57836 251284 57840
rect 252324 57836 252388 57900
rect 253428 57896 253492 57900
rect 253428 57840 253442 57896
rect 253442 57840 253492 57896
rect 253428 57836 253492 57840
rect 254532 57836 254596 57900
rect 183140 57760 183204 57764
rect 183140 57704 183190 57760
rect 183190 57704 183204 57760
rect 183140 57700 183204 57704
rect 206140 57700 206204 57764
rect 270908 57836 270972 57900
rect 271276 57896 271340 57900
rect 271276 57840 271290 57896
rect 271290 57840 271340 57896
rect 271276 57836 271340 57840
rect 273300 57896 273364 57900
rect 273300 57840 273314 57896
rect 273314 57840 273364 57896
rect 273300 57836 273364 57840
rect 278084 57896 278148 57900
rect 278084 57840 278098 57896
rect 278098 57840 278148 57896
rect 278084 57836 278148 57840
rect 279004 57896 279068 57900
rect 279004 57840 279054 57896
rect 279054 57840 279068 57896
rect 279004 57836 279068 57840
rect 288204 57836 288268 57900
rect 293356 57896 293420 57900
rect 293356 57840 293370 57896
rect 293370 57840 293420 57896
rect 293356 57836 293420 57840
rect 305868 57896 305932 57900
rect 305868 57840 305882 57896
rect 305882 57840 305932 57896
rect 305868 57836 305932 57840
rect 311020 57896 311084 57900
rect 311020 57840 311034 57896
rect 311034 57840 311084 57896
rect 311020 57836 311084 57840
rect 313412 57896 313476 57900
rect 313412 57840 313426 57896
rect 313426 57840 313476 57896
rect 313412 57836 313476 57840
rect 318380 57836 318444 57900
rect 343220 57896 343284 57900
rect 343220 57840 343234 57896
rect 343234 57840 343284 57896
rect 343220 57836 343284 57840
rect 343404 57896 343468 57900
rect 343404 57840 343454 57896
rect 343454 57840 343468 57896
rect 343404 57836 343468 57840
rect 399524 57836 399588 57900
rect 400444 57896 400508 57900
rect 400444 57840 400458 57896
rect 400458 57840 400508 57896
rect 400444 57836 400508 57840
rect 404124 57896 404188 57900
rect 404124 57840 404138 57896
rect 404138 57840 404188 57896
rect 404124 57836 404188 57840
rect 405044 57836 405108 57900
rect 406516 57836 406580 57900
rect 407620 57836 407684 57900
rect 408356 57896 408420 57900
rect 408356 57840 408370 57896
rect 408370 57840 408420 57896
rect 408356 57836 408420 57840
rect 408724 57896 408788 57900
rect 408724 57840 408738 57896
rect 408738 57840 408788 57896
rect 408724 57836 408788 57840
rect 410012 57836 410076 57900
rect 412404 57836 412468 57900
rect 413508 57896 413572 57900
rect 413508 57840 413522 57896
rect 413522 57840 413572 57896
rect 413508 57836 413572 57840
rect 414612 57896 414676 57900
rect 414612 57840 414626 57896
rect 414626 57840 414676 57896
rect 414612 57836 414676 57840
rect 418476 57896 418540 57900
rect 418476 57840 418490 57896
rect 418490 57840 418540 57896
rect 418476 57836 418540 57840
rect 422892 57896 422956 57900
rect 422892 57840 422906 57896
rect 422906 57840 422956 57896
rect 422892 57836 422956 57840
rect 423996 57836 424060 57900
rect 426388 57836 426452 57900
rect 427676 57896 427740 57900
rect 427676 57840 427690 57896
rect 427690 57840 427740 57896
rect 427676 57836 427740 57840
rect 428596 57836 428660 57900
rect 429700 57896 429764 57900
rect 429700 57840 429714 57896
rect 429714 57840 429764 57896
rect 429700 57836 429764 57840
rect 430988 57896 431052 57900
rect 430988 57840 431002 57896
rect 431002 57840 431052 57896
rect 430988 57836 431052 57840
rect 432276 57836 432340 57900
rect 433380 57896 433444 57900
rect 433380 57840 433394 57896
rect 433394 57840 433444 57896
rect 433380 57836 433444 57840
rect 433564 57896 433628 57900
rect 433564 57840 433578 57896
rect 433578 57840 433628 57896
rect 433564 57836 433628 57840
rect 435772 57836 435836 57900
rect 435956 57896 436020 57900
rect 435956 57840 435970 57896
rect 435970 57840 436020 57896
rect 435956 57836 436020 57840
rect 438532 57896 438596 57900
rect 438532 57840 438546 57896
rect 438546 57840 438596 57896
rect 438532 57836 438596 57840
rect 460980 57896 461044 57900
rect 460980 57840 460994 57896
rect 460994 57840 461044 57896
rect 263548 57760 263612 57764
rect 263548 57704 263598 57760
rect 263598 57704 263612 57760
rect 263548 57700 263612 57704
rect 265940 57700 266004 57764
rect 267596 57700 267660 57764
rect 268332 57700 268396 57764
rect 268700 57760 268764 57764
rect 268700 57704 268714 57760
rect 268714 57704 268764 57760
rect 268700 57700 268764 57704
rect 269804 57700 269868 57764
rect 274404 57700 274468 57764
rect 276980 57700 277044 57764
rect 372108 57700 372172 57764
rect 460980 57836 461044 57840
rect 465948 57896 466012 57900
rect 465948 57840 465962 57896
rect 465962 57840 466012 57896
rect 465948 57836 466012 57840
rect 470916 57896 470980 57900
rect 470916 57840 470930 57896
rect 470930 57840 470980 57896
rect 470916 57836 470980 57840
rect 475884 57896 475948 57900
rect 475884 57840 475898 57896
rect 475898 57840 475948 57896
rect 475884 57836 475948 57840
rect 480668 57896 480732 57900
rect 480668 57840 480682 57896
rect 480682 57840 480732 57896
rect 480668 57836 480732 57840
rect 483428 57896 483492 57900
rect 483428 57840 483442 57896
rect 483442 57840 483492 57896
rect 483428 57836 483492 57840
rect 503300 57896 503364 57900
rect 503300 57840 503350 57896
rect 503350 57840 503364 57896
rect 503300 57836 503364 57840
rect 54892 57564 54956 57628
rect 58940 57428 59004 57492
rect 112116 57428 112180 57492
rect 113220 57488 113284 57492
rect 115796 57564 115860 57628
rect 119108 57564 119172 57628
rect 155908 57624 155972 57628
rect 155908 57568 155958 57624
rect 155958 57568 155972 57624
rect 155908 57564 155972 57568
rect 160876 57564 160940 57628
rect 165844 57564 165908 57628
rect 215892 57564 215956 57628
rect 280844 57564 280908 57628
rect 370452 57564 370516 57628
rect 451044 57564 451108 57628
rect 113220 57432 113234 57488
rect 113234 57432 113284 57488
rect 113220 57428 113284 57432
rect 118372 57428 118436 57492
rect 213132 57428 213196 57492
rect 273484 57428 273548 57492
rect 360700 57428 360764 57492
rect 434668 57428 434732 57492
rect 436876 57428 436940 57492
rect 439084 57428 439148 57492
rect 58572 57292 58636 57356
rect 103836 57292 103900 57356
rect 202276 57292 202340 57356
rect 260972 57292 261036 57356
rect 266308 57352 266372 57356
rect 266308 57296 266358 57352
rect 266358 57296 266372 57352
rect 266308 57292 266372 57296
rect 376156 57292 376220 57356
rect 448284 57292 448348 57356
rect 57652 57156 57716 57220
rect 58756 57020 58820 57084
rect 88380 57080 88444 57084
rect 88380 57024 88430 57080
rect 88430 57024 88444 57080
rect 88380 57020 88444 57024
rect 105860 57156 105924 57220
rect 203196 57156 203260 57220
rect 256004 57156 256068 57220
rect 378732 57156 378796 57220
rect 445892 57156 445956 57220
rect 97028 57020 97092 57084
rect 216076 57020 216140 57084
rect 253612 57020 253676 57084
rect 376340 57020 376404 57084
rect 415532 57020 415596 57084
rect 431172 57020 431236 57084
rect 440924 57020 440988 57084
rect 96292 56884 96356 56948
rect 237052 56884 237116 56948
rect 411300 56944 411364 56948
rect 411300 56888 411314 56944
rect 411314 56888 411364 56944
rect 411300 56884 411364 56888
rect 52316 56612 52380 56676
rect 133460 56612 133524 56676
rect 163268 56612 163332 56676
rect 211660 56612 211724 56676
rect 285996 56612 286060 56676
rect 320956 56612 321020 56676
rect 323348 56612 323412 56676
rect 358124 56612 358188 56676
rect 443500 56748 443564 56812
rect 438348 56612 438412 56676
rect 53604 56476 53668 56540
rect 205404 56476 205468 56540
rect 48636 56340 48700 56404
rect 158484 56340 158548 56404
rect 209636 56340 209700 56404
rect 377260 56476 377324 56540
rect 52132 56204 52196 56268
rect 206876 56204 206940 56268
rect 57836 56068 57900 56132
rect 197860 56068 197924 56132
rect 50660 55116 50724 55180
rect 377812 55116 377876 55180
rect 50476 54980 50540 55044
rect 217364 54980 217428 55044
rect 379468 54980 379532 55044
rect 50844 54844 50908 54908
rect 57468 54708 57532 54772
rect 208900 3980 208964 4044
rect 204852 3844 204916 3908
rect 210372 3708 210436 3772
rect 371740 3572 371804 3636
rect 363460 3436 363524 3500
rect 364932 3300 364996 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 44035 487796 44101 487797
rect 44035 487732 44036 487796
rect 44100 487732 44101 487796
rect 44035 487731 44101 487732
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 44038 251021 44098 487731
rect 44955 482220 45021 482221
rect 44955 482156 44956 482220
rect 45020 482156 45021 482220
rect 44955 482155 45021 482156
rect 44771 471748 44837 471749
rect 44771 471684 44772 471748
rect 44836 471684 44837 471748
rect 44771 471683 44837 471684
rect 44774 379133 44834 471683
rect 44771 379132 44837 379133
rect 44771 379068 44772 379132
rect 44836 379068 44837 379132
rect 44771 379067 44837 379068
rect 44958 251157 45018 482155
rect 45234 478894 45854 514338
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 54339 646236 54405 646237
rect 54339 646172 54340 646236
rect 54404 646172 54405 646236
rect 54339 646171 54405 646172
rect 51579 646100 51645 646101
rect 51579 646036 51580 646100
rect 51644 646036 51645 646100
rect 51579 646035 51645 646036
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 46795 490652 46861 490653
rect 46795 490588 46796 490652
rect 46860 490588 46861 490652
rect 46795 490587 46861 490588
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 46611 468756 46677 468757
rect 46611 468692 46612 468756
rect 46676 468692 46677 468756
rect 46611 468691 46677 468692
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 44955 251156 45021 251157
rect 44955 251092 44956 251156
rect 45020 251092 45021 251156
rect 44955 251091 45021 251092
rect 44035 251020 44101 251021
rect 44035 250956 44036 251020
rect 44100 250956 44101 251020
rect 44035 250955 44101 250956
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 46614 58717 46674 468691
rect 46798 67829 46858 490587
rect 48954 482614 49574 518058
rect 50843 490516 50909 490517
rect 50843 490452 50844 490516
rect 50908 490452 50909 490516
rect 50843 490451 50909 490452
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 47715 482356 47781 482357
rect 47715 482292 47716 482356
rect 47780 482292 47781 482356
rect 47715 482291 47781 482292
rect 48954 482294 49574 482378
rect 47718 271149 47778 482291
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 47899 471204 47965 471205
rect 47899 471140 47900 471204
rect 47964 471140 47965 471204
rect 47899 471139 47965 471140
rect 47715 271148 47781 271149
rect 47715 271084 47716 271148
rect 47780 271084 47781 271148
rect 47715 271083 47781 271084
rect 47902 165069 47962 471139
rect 48083 468892 48149 468893
rect 48083 468828 48084 468892
rect 48148 468828 48149 468892
rect 48083 468827 48149 468828
rect 47899 165068 47965 165069
rect 47899 165004 47900 165068
rect 47964 165004 47965 165068
rect 47899 165003 47965 165004
rect 46795 67828 46861 67829
rect 46795 67764 46796 67828
rect 46860 67764 46861 67828
rect 46795 67763 46861 67764
rect 48086 58853 48146 468827
rect 48635 465764 48701 465765
rect 48635 465700 48636 465764
rect 48700 465700 48701 465764
rect 48635 465699 48701 465700
rect 48083 58852 48149 58853
rect 48083 58788 48084 58852
rect 48148 58788 48149 58852
rect 48083 58787 48149 58788
rect 46611 58716 46677 58717
rect 46611 58652 46612 58716
rect 46676 58652 46677 58716
rect 46611 58651 46677 58652
rect 48638 56405 48698 465699
rect 48954 446614 49574 482058
rect 50659 468484 50725 468485
rect 50659 468420 50660 468484
rect 50724 468420 50725 468484
rect 50659 468419 50725 468420
rect 50475 465220 50541 465221
rect 50475 465156 50476 465220
rect 50540 465156 50541 465220
rect 50475 465155 50541 465156
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48635 56404 48701 56405
rect 48635 56340 48636 56404
rect 48700 56340 48701 56404
rect 48635 56339 48701 56340
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 50614 49574 86058
rect 50478 55045 50538 465155
rect 50662 55181 50722 468419
rect 50659 55180 50725 55181
rect 50659 55116 50660 55180
rect 50724 55116 50725 55180
rect 50659 55115 50725 55116
rect 50475 55044 50541 55045
rect 50475 54980 50476 55044
rect 50540 54980 50541 55044
rect 50475 54979 50541 54980
rect 50846 54909 50906 490451
rect 51582 201517 51642 646035
rect 53051 645964 53117 645965
rect 53051 645900 53052 645964
rect 53116 645900 53117 645964
rect 53051 645899 53117 645900
rect 52315 490516 52381 490517
rect 52315 490452 52316 490516
rect 52380 490452 52381 490516
rect 52315 490451 52381 490452
rect 51947 466036 52013 466037
rect 51947 465972 51948 466036
rect 52012 465972 52013 466036
rect 51947 465971 52013 465972
rect 51950 379541 52010 465971
rect 52131 465900 52197 465901
rect 52131 465836 52132 465900
rect 52196 465836 52197 465900
rect 52131 465835 52197 465836
rect 51947 379540 52013 379541
rect 51947 379476 51948 379540
rect 52012 379476 52013 379540
rect 51947 379475 52013 379476
rect 51579 201516 51645 201517
rect 51579 201452 51580 201516
rect 51644 201452 51645 201516
rect 51579 201451 51645 201452
rect 52134 56269 52194 465835
rect 52318 56677 52378 490451
rect 53054 305013 53114 645899
rect 53603 468620 53669 468621
rect 53603 468556 53604 468620
rect 53668 468556 53669 468620
rect 53603 468555 53669 468556
rect 53419 466444 53485 466445
rect 53419 466380 53420 466444
rect 53484 466380 53485 466444
rect 53419 466379 53485 466380
rect 53235 466172 53301 466173
rect 53235 466108 53236 466172
rect 53300 466108 53301 466172
rect 53235 466107 53301 466108
rect 53238 388517 53298 466107
rect 53235 388516 53301 388517
rect 53235 388452 53236 388516
rect 53300 388452 53301 388516
rect 53235 388451 53301 388452
rect 53051 305012 53117 305013
rect 53051 304948 53052 305012
rect 53116 304948 53117 305012
rect 53051 304947 53117 304948
rect 53422 59125 53482 466379
rect 53419 59124 53485 59125
rect 53419 59060 53420 59124
rect 53484 59060 53485 59124
rect 53419 59059 53485 59060
rect 52315 56676 52381 56677
rect 52315 56612 52316 56676
rect 52380 56612 52381 56676
rect 52315 56611 52381 56612
rect 53606 56541 53666 468555
rect 54342 254013 54402 646171
rect 55794 633454 56414 668898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 645099 60134 672618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 645099 63854 676338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 645099 67574 680058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 645099 74414 650898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 645099 78134 654618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 645099 81854 658338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 645099 85574 662058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 645099 92414 668898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 645099 96134 672618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 645099 99854 676338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 645099 103574 680058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 645099 110414 650898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 645099 114134 654618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 645099 117854 658338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 645099 121574 662058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 79568 633454 79888 633486
rect 79568 633218 79610 633454
rect 79846 633218 79888 633454
rect 79568 633134 79888 633218
rect 79568 632898 79610 633134
rect 79846 632898 79888 633134
rect 79568 632866 79888 632898
rect 110288 633454 110608 633486
rect 110288 633218 110330 633454
rect 110566 633218 110608 633454
rect 110288 633134 110608 633218
rect 110288 632898 110330 633134
rect 110566 632898 110608 633134
rect 110288 632866 110608 632898
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 64208 615454 64528 615486
rect 64208 615218 64250 615454
rect 64486 615218 64528 615454
rect 64208 615134 64528 615218
rect 64208 614898 64250 615134
rect 64486 614898 64528 615134
rect 64208 614866 64528 614898
rect 94928 615454 95248 615486
rect 94928 615218 94970 615454
rect 95206 615218 95248 615454
rect 94928 615134 95248 615218
rect 94928 614898 94970 615134
rect 95206 614898 95248 615134
rect 94928 614866 95248 614898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 79568 597454 79888 597486
rect 79568 597218 79610 597454
rect 79846 597218 79888 597454
rect 79568 597134 79888 597218
rect 79568 596898 79610 597134
rect 79846 596898 79888 597134
rect 79568 596866 79888 596898
rect 110288 597454 110608 597486
rect 110288 597218 110330 597454
rect 110566 597218 110608 597454
rect 110288 597134 110608 597218
rect 110288 596898 110330 597134
rect 110566 596898 110608 597134
rect 110288 596866 110608 596898
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 59514 565174 60134 578000
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 555000 60134 564618
rect 63234 568894 63854 578000
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 555000 63854 568338
rect 66954 572614 67574 578000
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 555000 67574 572058
rect 73794 562394 74414 578000
rect 73794 562158 73826 562394
rect 74062 562158 74146 562394
rect 74382 562158 74414 562394
rect 73794 562074 74414 562158
rect 73794 561838 73826 562074
rect 74062 561838 74146 562074
rect 74382 561838 74414 562074
rect 73794 555000 74414 561838
rect 77514 566114 78134 578000
rect 77514 565878 77546 566114
rect 77782 565878 77866 566114
rect 78102 565878 78134 566114
rect 77514 565794 78134 565878
rect 77514 565558 77546 565794
rect 77782 565558 77866 565794
rect 78102 565558 78134 565794
rect 77514 555000 78134 565558
rect 81234 567954 81854 578000
rect 81234 567718 81266 567954
rect 81502 567718 81586 567954
rect 81822 567718 81854 567954
rect 81234 567634 81854 567718
rect 81234 567398 81266 567634
rect 81502 567398 81586 567634
rect 81822 567398 81854 567634
rect 81234 555000 81854 567398
rect 84954 571674 85574 578000
rect 84954 571438 84986 571674
rect 85222 571438 85306 571674
rect 85542 571438 85574 571674
rect 84954 571354 85574 571438
rect 84954 571118 84986 571354
rect 85222 571118 85306 571354
rect 85542 571118 85574 571354
rect 84954 555000 85574 571118
rect 91794 561454 92414 578000
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 555000 92414 560898
rect 95514 565174 96134 578000
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 555000 96134 564618
rect 99234 568894 99854 578000
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 555000 99854 568338
rect 102954 572614 103574 578000
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 555000 103574 572058
rect 109794 562394 110414 578000
rect 109794 562158 109826 562394
rect 110062 562158 110146 562394
rect 110382 562158 110414 562394
rect 109794 562074 110414 562158
rect 109794 561838 109826 562074
rect 110062 561838 110146 562074
rect 110382 561838 110414 562074
rect 109794 555000 110414 561838
rect 113514 566114 114134 578000
rect 113514 565878 113546 566114
rect 113782 565878 113866 566114
rect 114102 565878 114134 566114
rect 113514 565794 114134 565878
rect 113514 565558 113546 565794
rect 113782 565558 113866 565794
rect 114102 565558 114134 565794
rect 113514 555000 114134 565558
rect 117234 567954 117854 578000
rect 117234 567718 117266 567954
rect 117502 567718 117586 567954
rect 117822 567718 117854 567954
rect 117234 567634 117854 567718
rect 117234 567398 117266 567634
rect 117502 567398 117586 567634
rect 117822 567398 117854 567634
rect 117234 555000 117854 567398
rect 120954 571674 121574 578000
rect 120954 571438 120986 571674
rect 121222 571438 121306 571674
rect 121542 571438 121574 571674
rect 120954 571354 121574 571438
rect 120954 571118 120986 571354
rect 121222 571118 121306 571354
rect 121542 571118 121574 571354
rect 120954 555000 121574 571118
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 555000 128414 560898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 555000 132134 564618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 555000 135854 568338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 555000 139574 572058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 645099 150134 654618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 645099 153854 658338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 645099 157574 662058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 645099 164414 668898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 645099 168134 672618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 645099 171854 676338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 645099 175574 680058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 645099 182414 650898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 645099 186134 654618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 645099 189854 658338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 645099 193574 662058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 645099 200414 668898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 645099 204134 672618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 645099 207854 676338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 645099 211574 680058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 169568 633454 169888 633486
rect 169568 633218 169610 633454
rect 169846 633218 169888 633454
rect 169568 633134 169888 633218
rect 169568 632898 169610 633134
rect 169846 632898 169888 633134
rect 169568 632866 169888 632898
rect 200288 633454 200608 633486
rect 200288 633218 200330 633454
rect 200566 633218 200608 633454
rect 200288 633134 200608 633218
rect 200288 632898 200330 633134
rect 200566 632898 200608 633134
rect 200288 632866 200608 632898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 154208 615454 154528 615486
rect 154208 615218 154250 615454
rect 154486 615218 154528 615454
rect 154208 615134 154528 615218
rect 154208 614898 154250 615134
rect 154486 614898 154528 615134
rect 154208 614866 154528 614898
rect 184928 615454 185248 615486
rect 184928 615218 184970 615454
rect 185206 615218 185248 615454
rect 184928 615134 185248 615218
rect 184928 614898 184970 615134
rect 185206 614898 185248 615134
rect 184928 614866 185248 614898
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 169568 597454 169888 597486
rect 169568 597218 169610 597454
rect 169846 597218 169888 597454
rect 169568 597134 169888 597218
rect 169568 596898 169610 597134
rect 169846 596898 169888 597134
rect 169568 596866 169888 596898
rect 200288 597454 200608 597486
rect 200288 597218 200330 597454
rect 200566 597218 200608 597454
rect 200288 597134 200608 597218
rect 200288 596898 200330 597134
rect 200566 596898 200608 597134
rect 200288 596866 200608 596898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 562394 146414 578898
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 145794 562158 145826 562394
rect 146062 562158 146146 562394
rect 146382 562158 146414 562394
rect 145794 562074 146414 562158
rect 145794 561838 145826 562074
rect 146062 561838 146146 562074
rect 146382 561838 146414 562074
rect 145794 555000 146414 561838
rect 149514 566114 150134 578000
rect 149514 565878 149546 566114
rect 149782 565878 149866 566114
rect 150102 565878 150134 566114
rect 149514 565794 150134 565878
rect 149514 565558 149546 565794
rect 149782 565558 149866 565794
rect 150102 565558 150134 565794
rect 149514 555000 150134 565558
rect 153234 567954 153854 578000
rect 153234 567718 153266 567954
rect 153502 567718 153586 567954
rect 153822 567718 153854 567954
rect 153234 567634 153854 567718
rect 153234 567398 153266 567634
rect 153502 567398 153586 567634
rect 153822 567398 153854 567634
rect 153234 555000 153854 567398
rect 156954 571674 157574 578000
rect 156954 571438 156986 571674
rect 157222 571438 157306 571674
rect 157542 571438 157574 571674
rect 156954 571354 157574 571438
rect 156954 571118 156986 571354
rect 157222 571118 157306 571354
rect 157542 571118 157574 571354
rect 156954 555000 157574 571118
rect 163794 561454 164414 578000
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 555000 164414 560898
rect 167514 565174 168134 578000
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 555000 168134 564618
rect 171234 568894 171854 578000
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 555000 171854 568338
rect 174954 572614 175574 578000
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 555000 175574 572058
rect 181794 562394 182414 578000
rect 181794 562158 181826 562394
rect 182062 562158 182146 562394
rect 182382 562158 182414 562394
rect 181794 562074 182414 562158
rect 181794 561838 181826 562074
rect 182062 561838 182146 562074
rect 182382 561838 182414 562074
rect 181794 555000 182414 561838
rect 185514 566114 186134 578000
rect 185514 565878 185546 566114
rect 185782 565878 185866 566114
rect 186102 565878 186134 566114
rect 185514 565794 186134 565878
rect 185514 565558 185546 565794
rect 185782 565558 185866 565794
rect 186102 565558 186134 565794
rect 185514 555000 186134 565558
rect 189234 567954 189854 578000
rect 189234 567718 189266 567954
rect 189502 567718 189586 567954
rect 189822 567718 189854 567954
rect 189234 567634 189854 567718
rect 189234 567398 189266 567634
rect 189502 567398 189586 567634
rect 189822 567398 189854 567634
rect 189234 555000 189854 567398
rect 192954 571674 193574 578000
rect 192954 571438 192986 571674
rect 193222 571438 193306 571674
rect 193542 571438 193574 571674
rect 192954 571354 193574 571438
rect 192954 571118 192986 571354
rect 193222 571118 193306 571354
rect 193542 571118 193574 571354
rect 192954 555000 193574 571118
rect 199794 561454 200414 578000
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 555000 200414 560898
rect 203514 565174 204134 578000
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 555000 204134 564618
rect 207234 568894 207854 578000
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 555000 207854 568338
rect 210954 572614 211574 578000
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 555000 211574 572058
rect 217794 562394 218414 578898
rect 217794 562158 217826 562394
rect 218062 562158 218146 562394
rect 218382 562158 218414 562394
rect 217794 562074 218414 562158
rect 217794 561838 217826 562074
rect 218062 561838 218146 562074
rect 218382 561838 218414 562074
rect 217794 555000 218414 561838
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 566114 222134 582618
rect 221514 565878 221546 566114
rect 221782 565878 221866 566114
rect 222102 565878 222134 566114
rect 221514 565794 222134 565878
rect 221514 565558 221546 565794
rect 221782 565558 221866 565794
rect 222102 565558 222134 565794
rect 221514 555000 222134 565558
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 567954 225854 586338
rect 225234 567718 225266 567954
rect 225502 567718 225586 567954
rect 225822 567718 225854 567954
rect 225234 567634 225854 567718
rect 225234 567398 225266 567634
rect 225502 567398 225586 567634
rect 225822 567398 225854 567634
rect 225234 555000 225854 567398
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 571674 229574 590058
rect 228954 571438 228986 571674
rect 229222 571438 229306 571674
rect 229542 571438 229574 571674
rect 228954 571354 229574 571438
rect 228954 571118 228986 571354
rect 229222 571118 229306 571354
rect 229542 571118 229574 571354
rect 228954 555000 229574 571118
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 645099 240134 672618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 645099 243854 676338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 645099 247574 680058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 645099 254414 650898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 645099 258134 654618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 645099 261854 658338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 645099 265574 662058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 645099 272414 668898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 645099 276134 672618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 645099 279854 676338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 645099 283574 680058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 645099 290414 650898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 645099 294134 654618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 645099 297854 658338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 645099 301574 662058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 259568 633454 259888 633486
rect 259568 633218 259610 633454
rect 259846 633218 259888 633454
rect 259568 633134 259888 633218
rect 259568 632898 259610 633134
rect 259846 632898 259888 633134
rect 259568 632866 259888 632898
rect 290288 633454 290608 633486
rect 290288 633218 290330 633454
rect 290566 633218 290608 633454
rect 290288 633134 290608 633218
rect 290288 632898 290330 633134
rect 290566 632898 290608 633134
rect 290288 632866 290608 632898
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 244208 615454 244528 615486
rect 244208 615218 244250 615454
rect 244486 615218 244528 615454
rect 244208 615134 244528 615218
rect 244208 614898 244250 615134
rect 244486 614898 244528 615134
rect 244208 614866 244528 614898
rect 274928 615454 275248 615486
rect 274928 615218 274970 615454
rect 275206 615218 275248 615454
rect 274928 615134 275248 615218
rect 274928 614898 274970 615134
rect 275206 614898 275248 615134
rect 274928 614866 275248 614898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 259568 597454 259888 597486
rect 259568 597218 259610 597454
rect 259846 597218 259888 597454
rect 259568 597134 259888 597218
rect 259568 596898 259610 597134
rect 259846 596898 259888 597134
rect 259568 596866 259888 596898
rect 290288 597454 290608 597486
rect 290288 597218 290330 597454
rect 290566 597218 290608 597454
rect 290288 597134 290608 597218
rect 290288 596898 290330 597134
rect 290566 596898 290608 597134
rect 290288 596866 290608 596898
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 555000 236414 560898
rect 239514 565174 240134 578000
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 555000 240134 564618
rect 243234 568894 243854 578000
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 555000 243854 568338
rect 246954 572614 247574 578000
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 555000 247574 572058
rect 253794 562394 254414 578000
rect 253794 562158 253826 562394
rect 254062 562158 254146 562394
rect 254382 562158 254414 562394
rect 253794 562074 254414 562158
rect 253794 561838 253826 562074
rect 254062 561838 254146 562074
rect 254382 561838 254414 562074
rect 253794 555000 254414 561838
rect 257514 566114 258134 578000
rect 257514 565878 257546 566114
rect 257782 565878 257866 566114
rect 258102 565878 258134 566114
rect 257514 565794 258134 565878
rect 257514 565558 257546 565794
rect 257782 565558 257866 565794
rect 258102 565558 258134 565794
rect 257514 555000 258134 565558
rect 261234 567954 261854 578000
rect 261234 567718 261266 567954
rect 261502 567718 261586 567954
rect 261822 567718 261854 567954
rect 261234 567634 261854 567718
rect 261234 567398 261266 567634
rect 261502 567398 261586 567634
rect 261822 567398 261854 567634
rect 261234 555000 261854 567398
rect 264954 571674 265574 578000
rect 264954 571438 264986 571674
rect 265222 571438 265306 571674
rect 265542 571438 265574 571674
rect 264954 571354 265574 571438
rect 264954 571118 264986 571354
rect 265222 571118 265306 571354
rect 265542 571118 265574 571354
rect 264954 555000 265574 571118
rect 271794 561454 272414 578000
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 555000 272414 560898
rect 275514 565174 276134 578000
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 555000 276134 564618
rect 279234 568894 279854 578000
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 555000 279854 568338
rect 282954 572614 283574 578000
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 555000 283574 572058
rect 289794 562394 290414 578000
rect 289794 562158 289826 562394
rect 290062 562158 290146 562394
rect 290382 562158 290414 562394
rect 289794 562074 290414 562158
rect 289794 561838 289826 562074
rect 290062 561838 290146 562074
rect 290382 561838 290414 562074
rect 289794 555000 290414 561838
rect 293514 566114 294134 578000
rect 293514 565878 293546 566114
rect 293782 565878 293866 566114
rect 294102 565878 294134 566114
rect 293514 565794 294134 565878
rect 293514 565558 293546 565794
rect 293782 565558 293866 565794
rect 294102 565558 294134 565794
rect 293514 555000 294134 565558
rect 297234 567954 297854 578000
rect 297234 567718 297266 567954
rect 297502 567718 297586 567954
rect 297822 567718 297854 567954
rect 297234 567634 297854 567718
rect 297234 567398 297266 567634
rect 297502 567398 297586 567634
rect 297822 567398 297854 567634
rect 297234 555000 297854 567398
rect 300954 571674 301574 578000
rect 300954 571438 300986 571674
rect 301222 571438 301306 571674
rect 301542 571438 301574 571674
rect 300954 571354 301574 571438
rect 300954 571118 300986 571354
rect 301222 571118 301306 571354
rect 301542 571118 301574 571354
rect 300954 555000 301574 571118
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 64208 543454 64528 543486
rect 64208 543218 64250 543454
rect 64486 543218 64528 543454
rect 64208 543134 64528 543218
rect 64208 542898 64250 543134
rect 64486 542898 64528 543134
rect 64208 542866 64528 542898
rect 94928 543454 95248 543486
rect 94928 543218 94970 543454
rect 95206 543218 95248 543454
rect 94928 543134 95248 543218
rect 94928 542898 94970 543134
rect 95206 542898 95248 543134
rect 94928 542866 95248 542898
rect 125648 543454 125968 543486
rect 125648 543218 125690 543454
rect 125926 543218 125968 543454
rect 125648 543134 125968 543218
rect 125648 542898 125690 543134
rect 125926 542898 125968 543134
rect 125648 542866 125968 542898
rect 156368 543454 156688 543486
rect 156368 543218 156410 543454
rect 156646 543218 156688 543454
rect 156368 543134 156688 543218
rect 156368 542898 156410 543134
rect 156646 542898 156688 543134
rect 156368 542866 156688 542898
rect 187088 543454 187408 543486
rect 187088 543218 187130 543454
rect 187366 543218 187408 543454
rect 187088 543134 187408 543218
rect 187088 542898 187130 543134
rect 187366 542898 187408 543134
rect 187088 542866 187408 542898
rect 217808 543454 218128 543486
rect 217808 543218 217850 543454
rect 218086 543218 218128 543454
rect 217808 543134 218128 543218
rect 217808 542898 217850 543134
rect 218086 542898 218128 543134
rect 217808 542866 218128 542898
rect 248528 543454 248848 543486
rect 248528 543218 248570 543454
rect 248806 543218 248848 543454
rect 248528 543134 248848 543218
rect 248528 542898 248570 543134
rect 248806 542898 248848 543134
rect 248528 542866 248848 542898
rect 279248 543454 279568 543486
rect 279248 543218 279290 543454
rect 279526 543218 279568 543454
rect 279248 543134 279568 543218
rect 279248 542898 279290 543134
rect 279526 542898 279568 543134
rect 279248 542866 279568 542898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 54891 490924 54957 490925
rect 54891 490860 54892 490924
rect 54956 490860 54957 490924
rect 54891 490859 54957 490860
rect 54707 466308 54773 466309
rect 54707 466244 54708 466308
rect 54772 466244 54773 466308
rect 54707 466243 54773 466244
rect 54339 254012 54405 254013
rect 54339 253948 54340 254012
rect 54404 253948 54405 254012
rect 54339 253947 54405 253948
rect 54710 59261 54770 466243
rect 54707 59260 54773 59261
rect 54707 59196 54708 59260
rect 54772 59196 54773 59260
rect 54707 59195 54773 59196
rect 54894 57629 54954 490859
rect 55075 490788 55141 490789
rect 55075 490724 55076 490788
rect 55140 490724 55141 490788
rect 55075 490723 55141 490724
rect 55078 57765 55138 490723
rect 55627 490108 55693 490109
rect 55627 490044 55628 490108
rect 55692 490044 55693 490108
rect 55627 490043 55693 490044
rect 55630 381037 55690 490043
rect 55794 489454 56414 524898
rect 79568 525454 79888 525486
rect 79568 525218 79610 525454
rect 79846 525218 79888 525454
rect 79568 525134 79888 525218
rect 79568 524898 79610 525134
rect 79846 524898 79888 525134
rect 79568 524866 79888 524898
rect 110288 525454 110608 525486
rect 110288 525218 110330 525454
rect 110566 525218 110608 525454
rect 110288 525134 110608 525218
rect 110288 524898 110330 525134
rect 110566 524898 110608 525134
rect 110288 524866 110608 524898
rect 141008 525454 141328 525486
rect 141008 525218 141050 525454
rect 141286 525218 141328 525454
rect 141008 525134 141328 525218
rect 141008 524898 141050 525134
rect 141286 524898 141328 525134
rect 141008 524866 141328 524898
rect 171728 525454 172048 525486
rect 171728 525218 171770 525454
rect 172006 525218 172048 525454
rect 171728 525134 172048 525218
rect 171728 524898 171770 525134
rect 172006 524898 172048 525134
rect 171728 524866 172048 524898
rect 202448 525454 202768 525486
rect 202448 525218 202490 525454
rect 202726 525218 202768 525454
rect 202448 525134 202768 525218
rect 202448 524898 202490 525134
rect 202726 524898 202768 525134
rect 202448 524866 202768 524898
rect 233168 525454 233488 525486
rect 233168 525218 233210 525454
rect 233446 525218 233488 525454
rect 233168 525134 233488 525218
rect 233168 524898 233210 525134
rect 233446 524898 233488 525134
rect 233168 524866 233488 524898
rect 263888 525454 264208 525486
rect 263888 525218 263930 525454
rect 264166 525218 264208 525454
rect 263888 525134 264208 525218
rect 263888 524898 263930 525134
rect 264166 524898 264208 525134
rect 263888 524866 264208 524898
rect 294608 525454 294928 525486
rect 294608 525218 294650 525454
rect 294886 525218 294928 525454
rect 294608 525134 294928 525218
rect 294608 524898 294650 525134
rect 294886 524898 294928 525134
rect 294608 524866 294928 524898
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 64208 507454 64528 507486
rect 64208 507218 64250 507454
rect 64486 507218 64528 507454
rect 64208 507134 64528 507218
rect 64208 506898 64250 507134
rect 64486 506898 64528 507134
rect 64208 506866 64528 506898
rect 94928 507454 95248 507486
rect 94928 507218 94970 507454
rect 95206 507218 95248 507454
rect 94928 507134 95248 507218
rect 94928 506898 94970 507134
rect 95206 506898 95248 507134
rect 94928 506866 95248 506898
rect 125648 507454 125968 507486
rect 125648 507218 125690 507454
rect 125926 507218 125968 507454
rect 125648 507134 125968 507218
rect 125648 506898 125690 507134
rect 125926 506898 125968 507134
rect 125648 506866 125968 506898
rect 156368 507454 156688 507486
rect 156368 507218 156410 507454
rect 156646 507218 156688 507454
rect 156368 507134 156688 507218
rect 156368 506898 156410 507134
rect 156646 506898 156688 507134
rect 156368 506866 156688 506898
rect 187088 507454 187408 507486
rect 187088 507218 187130 507454
rect 187366 507218 187408 507454
rect 187088 507134 187408 507218
rect 187088 506898 187130 507134
rect 187366 506898 187408 507134
rect 187088 506866 187408 506898
rect 217808 507454 218128 507486
rect 217808 507218 217850 507454
rect 218086 507218 218128 507454
rect 217808 507134 218128 507218
rect 217808 506898 217850 507134
rect 218086 506898 218128 507134
rect 217808 506866 218128 506898
rect 248528 507454 248848 507486
rect 248528 507218 248570 507454
rect 248806 507218 248848 507454
rect 248528 507134 248848 507218
rect 248528 506898 248570 507134
rect 248806 506898 248848 507134
rect 248528 506866 248848 506898
rect 279248 507454 279568 507486
rect 279248 507218 279290 507454
rect 279526 507218 279568 507454
rect 279248 507134 279568 507218
rect 279248 506898 279290 507134
rect 279526 506898 279568 507134
rect 279248 506866 279568 506898
rect 208899 491876 208965 491877
rect 208899 491812 208900 491876
rect 208964 491812 208965 491876
rect 208899 491811 208965 491812
rect 60227 491196 60293 491197
rect 60227 491132 60228 491196
rect 60292 491132 60293 491196
rect 60227 491131 60293 491132
rect 198227 491196 198293 491197
rect 198227 491132 198228 491196
rect 198292 491132 198293 491196
rect 198227 491131 198293 491132
rect 59307 490380 59373 490381
rect 59307 490316 59308 490380
rect 59372 490316 59373 490380
rect 59307 490315 59373 490316
rect 59123 490244 59189 490245
rect 59123 490180 59124 490244
rect 59188 490180 59189 490244
rect 59123 490179 59189 490180
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 57099 488340 57165 488341
rect 57099 488276 57100 488340
rect 57164 488276 57165 488340
rect 57099 488275 57165 488276
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55627 381036 55693 381037
rect 55627 380972 55628 381036
rect 55692 380972 55693 381036
rect 55627 380971 55693 380972
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 57102 378045 57162 488275
rect 57467 482492 57533 482493
rect 57467 482428 57468 482492
rect 57532 482428 57533 482492
rect 57467 482427 57533 482428
rect 57470 390693 57530 482427
rect 57835 471612 57901 471613
rect 57835 471548 57836 471612
rect 57900 471548 57901 471612
rect 57835 471547 57901 471548
rect 57651 464404 57717 464405
rect 57651 464340 57652 464404
rect 57716 464340 57717 464404
rect 57651 464339 57717 464340
rect 57467 390692 57533 390693
rect 57467 390628 57468 390692
rect 57532 390628 57533 390692
rect 57467 390627 57533 390628
rect 57099 378044 57165 378045
rect 57099 377980 57100 378044
rect 57164 377980 57165 378044
rect 57099 377979 57165 377980
rect 57467 357372 57533 357373
rect 57467 357308 57468 357372
rect 57532 357308 57533 357372
rect 57467 357307 57533 357308
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 57470 272509 57530 357307
rect 57467 272508 57533 272509
rect 57467 272444 57468 272508
rect 57532 272444 57533 272508
rect 57467 272443 57533 272444
rect 57467 252516 57533 252517
rect 57467 252452 57468 252516
rect 57532 252452 57533 252516
rect 57467 252451 57533 252452
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 57470 164253 57530 252451
rect 57654 166973 57714 464339
rect 57651 166972 57717 166973
rect 57651 166908 57652 166972
rect 57716 166908 57717 166972
rect 57651 166907 57717 166908
rect 57838 166837 57898 471547
rect 58939 469844 59005 469845
rect 58939 469780 58940 469844
rect 59004 469780 59005 469844
rect 58939 469779 59005 469780
rect 58755 467124 58821 467125
rect 58755 467060 58756 467124
rect 58820 467060 58821 467124
rect 58755 467059 58821 467060
rect 58571 465628 58637 465629
rect 58571 465564 58572 465628
rect 58636 465564 58637 465628
rect 58571 465563 58637 465564
rect 57835 166836 57901 166837
rect 57835 166772 57836 166836
rect 57900 166772 57901 166836
rect 57835 166771 57901 166772
rect 57467 164252 57533 164253
rect 57467 164188 57468 164252
rect 57532 164188 57533 164252
rect 57467 164187 57533 164188
rect 57835 163300 57901 163301
rect 57835 163236 57836 163300
rect 57900 163236 57901 163300
rect 57835 163235 57901 163236
rect 57651 145892 57717 145893
rect 57651 145828 57652 145892
rect 57716 145828 57717 145892
rect 57651 145827 57717 145828
rect 57467 140860 57533 140861
rect 57467 140796 57468 140860
rect 57532 140796 57533 140860
rect 57467 140795 57533 140796
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55075 57764 55141 57765
rect 55075 57700 55076 57764
rect 55140 57700 55141 57764
rect 55075 57699 55141 57700
rect 54891 57628 54957 57629
rect 54891 57564 54892 57628
rect 54956 57564 54957 57628
rect 54891 57563 54957 57564
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 53603 56540 53669 56541
rect 53603 56476 53604 56540
rect 53668 56476 53669 56540
rect 53603 56475 53669 56476
rect 52131 56268 52197 56269
rect 52131 56204 52132 56268
rect 52196 56204 52197 56268
rect 52131 56203 52197 56204
rect 50843 54908 50909 54909
rect 50843 54844 50844 54908
rect 50908 54844 50909 54908
rect 50843 54843 50909 54844
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 21454 56414 56898
rect 57470 54773 57530 140795
rect 57654 57221 57714 145827
rect 57651 57220 57717 57221
rect 57651 57156 57652 57220
rect 57716 57156 57717 57220
rect 57651 57155 57717 57156
rect 57838 56133 57898 163235
rect 58574 57357 58634 465563
rect 58571 57356 58637 57357
rect 58571 57292 58572 57356
rect 58636 57292 58637 57356
rect 58571 57291 58637 57292
rect 58758 57085 58818 467059
rect 58942 57493 59002 469779
rect 59126 58989 59186 490179
rect 59123 58988 59189 58989
rect 59123 58924 59124 58988
rect 59188 58924 59189 58988
rect 59123 58923 59189 58924
rect 59310 58445 59370 490315
rect 59514 476114 60134 491000
rect 59514 475878 59546 476114
rect 59782 475878 59866 476114
rect 60102 475878 60134 476114
rect 59514 475794 60134 475878
rect 59514 475558 59546 475794
rect 59782 475558 59866 475794
rect 60102 475558 60134 475794
rect 59514 466308 60134 475558
rect 60230 465490 60290 491131
rect 63234 479834 63854 491000
rect 63234 479598 63266 479834
rect 63502 479598 63586 479834
rect 63822 479598 63854 479834
rect 63234 479514 63854 479598
rect 63234 479278 63266 479514
rect 63502 479278 63586 479514
rect 63822 479278 63854 479514
rect 63234 466308 63854 479278
rect 66954 481674 67574 491000
rect 66954 481438 66986 481674
rect 67222 481438 67306 481674
rect 67542 481438 67574 481674
rect 66954 481354 67574 481438
rect 66954 481118 66986 481354
rect 67222 481118 67306 481354
rect 67542 481118 67574 481354
rect 66954 466308 67574 481118
rect 73794 471454 74414 491000
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 466308 74414 470898
rect 77514 475174 78134 491000
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 466308 78134 474618
rect 81234 478894 81854 491000
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 466308 81854 478338
rect 84954 482614 85574 491000
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 466308 85574 482058
rect 91794 489454 92414 491000
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 466308 92414 488898
rect 95514 476114 96134 491000
rect 95514 475878 95546 476114
rect 95782 475878 95866 476114
rect 96102 475878 96134 476114
rect 95514 475794 96134 475878
rect 95514 475558 95546 475794
rect 95782 475558 95866 475794
rect 96102 475558 96134 475794
rect 95514 466308 96134 475558
rect 99234 479834 99854 491000
rect 99234 479598 99266 479834
rect 99502 479598 99586 479834
rect 99822 479598 99854 479834
rect 99234 479514 99854 479598
rect 99234 479278 99266 479514
rect 99502 479278 99586 479514
rect 99822 479278 99854 479514
rect 99234 466308 99854 479278
rect 102954 481674 103574 491000
rect 102954 481438 102986 481674
rect 103222 481438 103306 481674
rect 103542 481438 103574 481674
rect 102954 481354 103574 481438
rect 102954 481118 102986 481354
rect 103222 481118 103306 481354
rect 103542 481118 103574 481354
rect 102954 466308 103574 481118
rect 109794 471454 110414 491000
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109794 466308 110414 470898
rect 113514 475174 114134 491000
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 113514 466308 114134 474618
rect 117234 478894 117854 491000
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 117234 466308 117854 478338
rect 120954 482614 121574 491000
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120954 466308 121574 482058
rect 127794 489454 128414 491000
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 466308 128414 488898
rect 131514 476114 132134 491000
rect 131514 475878 131546 476114
rect 131782 475878 131866 476114
rect 132102 475878 132134 476114
rect 131514 475794 132134 475878
rect 131514 475558 131546 475794
rect 131782 475558 131866 475794
rect 132102 475558 132134 475794
rect 131514 466308 132134 475558
rect 135234 479834 135854 491000
rect 135234 479598 135266 479834
rect 135502 479598 135586 479834
rect 135822 479598 135854 479834
rect 135234 479514 135854 479598
rect 135234 479278 135266 479514
rect 135502 479278 135586 479514
rect 135822 479278 135854 479514
rect 135234 466308 135854 479278
rect 138954 481674 139574 491000
rect 138954 481438 138986 481674
rect 139222 481438 139306 481674
rect 139542 481438 139574 481674
rect 138954 481354 139574 481438
rect 138954 481118 138986 481354
rect 139222 481118 139306 481354
rect 139542 481118 139574 481354
rect 138954 466308 139574 481118
rect 145794 471454 146414 491000
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 466308 146414 470898
rect 149514 475174 150134 491000
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 466308 150134 474618
rect 153234 478894 153854 491000
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 466308 153854 478338
rect 156954 482614 157574 491000
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 466308 157574 482058
rect 163794 489454 164414 491000
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 466308 164414 488898
rect 167514 476114 168134 491000
rect 167514 475878 167546 476114
rect 167782 475878 167866 476114
rect 168102 475878 168134 476114
rect 167514 475794 168134 475878
rect 167514 475558 167546 475794
rect 167782 475558 167866 475794
rect 168102 475558 168134 475794
rect 167514 466308 168134 475558
rect 171234 479834 171854 491000
rect 171234 479598 171266 479834
rect 171502 479598 171586 479834
rect 171822 479598 171854 479834
rect 171234 479514 171854 479598
rect 171234 479278 171266 479514
rect 171502 479278 171586 479514
rect 171822 479278 171854 479514
rect 171234 466308 171854 479278
rect 174954 481674 175574 491000
rect 174954 481438 174986 481674
rect 175222 481438 175306 481674
rect 175542 481438 175574 481674
rect 174954 481354 175574 481438
rect 174954 481118 174986 481354
rect 175222 481118 175306 481354
rect 175542 481118 175574 481354
rect 174954 466308 175574 481118
rect 181794 471454 182414 491000
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 178355 466580 178421 466581
rect 178355 466516 178356 466580
rect 178420 466516 178421 466580
rect 178355 466515 178421 466516
rect 179643 466580 179709 466581
rect 179643 466516 179644 466580
rect 179708 466516 179709 466580
rect 179643 466515 179709 466516
rect 59862 465430 60290 465490
rect 59862 379810 59922 465430
rect 178358 464810 178418 466515
rect 179646 464810 179706 466515
rect 181794 466308 182414 470898
rect 185514 475174 186134 491000
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 466308 186134 474618
rect 189234 478894 189854 491000
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 466308 189854 478338
rect 192954 482614 193574 491000
rect 196571 490924 196637 490925
rect 196571 490860 196572 490924
rect 196636 490860 196637 490924
rect 196571 490859 196637 490860
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 190867 466580 190933 466581
rect 190867 466516 190868 466580
rect 190932 466516 190933 466580
rect 190867 466515 190933 466516
rect 190870 464810 190930 466515
rect 192954 466308 193574 482058
rect 178358 464750 178524 464810
rect 179646 464750 179748 464810
rect 178464 464202 178524 464750
rect 179688 464202 179748 464750
rect 190840 464750 190930 464810
rect 190840 464202 190900 464750
rect 60272 453454 60620 453486
rect 60272 453218 60328 453454
rect 60564 453218 60620 453454
rect 60272 453134 60620 453218
rect 60272 452898 60328 453134
rect 60564 452898 60620 453134
rect 60272 452866 60620 452898
rect 196000 453454 196348 453486
rect 196000 453218 196056 453454
rect 196292 453218 196348 453454
rect 196000 453134 196348 453218
rect 196000 452898 196056 453134
rect 196292 452898 196348 453134
rect 196000 452866 196348 452898
rect 60952 435454 61300 435486
rect 60952 435218 61008 435454
rect 61244 435218 61300 435454
rect 60952 435134 61300 435218
rect 60952 434898 61008 435134
rect 61244 434898 61300 435134
rect 60952 434866 61300 434898
rect 195320 435454 195668 435486
rect 195320 435218 195376 435454
rect 195612 435218 195668 435454
rect 195320 435134 195668 435218
rect 195320 434898 195376 435134
rect 195612 434898 195668 435134
rect 195320 434866 195668 434898
rect 60272 417454 60620 417486
rect 60272 417218 60328 417454
rect 60564 417218 60620 417454
rect 60272 417134 60620 417218
rect 60272 416898 60328 417134
rect 60564 416898 60620 417134
rect 60272 416866 60620 416898
rect 196000 417454 196348 417486
rect 196000 417218 196056 417454
rect 196292 417218 196348 417454
rect 196000 417134 196348 417218
rect 196000 416898 196056 417134
rect 196292 416898 196348 417134
rect 196000 416866 196348 416898
rect 60952 399454 61300 399486
rect 60952 399218 61008 399454
rect 61244 399218 61300 399454
rect 60952 399134 61300 399218
rect 60952 398898 61008 399134
rect 61244 398898 61300 399134
rect 60952 398866 61300 398898
rect 195320 399454 195668 399486
rect 195320 399218 195376 399454
rect 195612 399218 195668 399454
rect 195320 399134 195668 399218
rect 195320 398898 195376 399134
rect 195612 398898 195668 399134
rect 195320 398866 195668 398898
rect 76056 380490 76116 381106
rect 76054 380430 76116 380490
rect 77144 380490 77204 381106
rect 78232 380490 78292 381106
rect 79592 380490 79652 381106
rect 80544 380898 80604 381106
rect 77144 380430 77218 380490
rect 78232 380430 78322 380490
rect 59862 379750 60290 379810
rect 59514 368114 60134 379000
rect 59514 367878 59546 368114
rect 59782 367878 59866 368114
rect 60102 367878 60134 368114
rect 59514 367794 60134 367878
rect 59514 367558 59546 367794
rect 59782 367558 59866 367794
rect 60102 367558 60134 367794
rect 59514 359308 60134 367558
rect 60230 358730 60290 379750
rect 63234 369954 63854 379000
rect 63234 369718 63266 369954
rect 63502 369718 63586 369954
rect 63822 369718 63854 369954
rect 63234 369634 63854 369718
rect 63234 369398 63266 369634
rect 63502 369398 63586 369634
rect 63822 369398 63854 369634
rect 63234 359308 63854 369398
rect 66954 373674 67574 379000
rect 66954 373438 66986 373674
rect 67222 373438 67306 373674
rect 67542 373438 67574 373674
rect 66954 373354 67574 373438
rect 66954 373118 66986 373354
rect 67222 373118 67306 373354
rect 67542 373118 67574 373354
rect 66954 359308 67574 373118
rect 73794 363454 74414 379000
rect 76054 378589 76114 380430
rect 77158 379405 77218 380430
rect 77155 379404 77221 379405
rect 77155 379340 77156 379404
rect 77220 379340 77221 379404
rect 77155 379339 77221 379340
rect 78262 379269 78322 380430
rect 79550 380430 79652 380490
rect 80470 380838 80604 380898
rect 78259 379268 78325 379269
rect 78259 379204 78260 379268
rect 78324 379204 78325 379268
rect 78259 379203 78325 379204
rect 76051 378588 76117 378589
rect 76051 378524 76052 378588
rect 76116 378524 76117 378588
rect 76051 378523 76117 378524
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 359308 74414 362898
rect 77514 367174 78134 379000
rect 78262 378997 78322 379203
rect 78259 378996 78325 378997
rect 78259 378932 78260 378996
rect 78324 378932 78325 378996
rect 78259 378931 78325 378932
rect 79550 378861 79610 380430
rect 80470 379405 80530 380838
rect 81768 380490 81828 381106
rect 83128 380765 83188 381106
rect 84216 380901 84276 381106
rect 84213 380900 84279 380901
rect 84213 380836 84214 380900
rect 84278 380836 84279 380900
rect 84213 380835 84279 380836
rect 83125 380764 83191 380765
rect 83125 380700 83126 380764
rect 83190 380700 83191 380764
rect 83125 380699 83191 380700
rect 85440 380490 85500 381106
rect 81758 380430 81828 380490
rect 85438 380430 85500 380490
rect 86528 380490 86588 381106
rect 87616 380490 87676 381106
rect 88296 380490 88356 381106
rect 88704 380490 88764 381106
rect 90064 380490 90124 381106
rect 86528 380430 86602 380490
rect 87616 380430 87706 380490
rect 88296 380430 88442 380490
rect 88704 380430 88810 380490
rect 80467 379404 80533 379405
rect 80467 379340 80468 379404
rect 80532 379340 80533 379404
rect 80467 379339 80533 379340
rect 81758 379269 81818 380430
rect 85438 379405 85498 380430
rect 86542 379405 86602 380430
rect 85435 379404 85501 379405
rect 85435 379340 85436 379404
rect 85500 379340 85501 379404
rect 85435 379339 85501 379340
rect 86539 379404 86605 379405
rect 86539 379340 86540 379404
rect 86604 379340 86605 379404
rect 86539 379339 86605 379340
rect 81755 379268 81821 379269
rect 81755 379204 81756 379268
rect 81820 379204 81821 379268
rect 81755 379203 81821 379204
rect 79547 378860 79613 378861
rect 79547 378796 79548 378860
rect 79612 378796 79613 378860
rect 79547 378795 79613 378796
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 359308 78134 366618
rect 81234 370894 81854 379000
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 359308 81854 370338
rect 84954 374614 85574 379000
rect 87646 378181 87706 380430
rect 88382 379405 88442 380430
rect 88750 379405 88810 380430
rect 90038 380430 90124 380490
rect 90744 380490 90804 381106
rect 91288 380490 91348 381106
rect 92376 380490 92436 381106
rect 93464 380490 93524 381106
rect 90744 380430 90834 380490
rect 91288 380430 91386 380490
rect 92376 380430 92490 380490
rect 88379 379404 88445 379405
rect 88379 379340 88380 379404
rect 88444 379340 88445 379404
rect 88379 379339 88445 379340
rect 88747 379404 88813 379405
rect 88747 379340 88748 379404
rect 88812 379340 88813 379404
rect 88747 379339 88813 379340
rect 90038 379269 90098 380430
rect 90774 379405 90834 380430
rect 91326 379405 91386 380430
rect 92430 379405 92490 380430
rect 93350 380430 93524 380490
rect 93600 380490 93660 381106
rect 94552 380629 94612 381106
rect 94549 380628 94615 380629
rect 94549 380564 94550 380628
rect 94614 380564 94615 380628
rect 94549 380563 94615 380564
rect 95912 380490 95972 381106
rect 96048 380490 96108 381106
rect 97000 380490 97060 381106
rect 98088 380490 98148 381106
rect 98496 380490 98556 381106
rect 99448 380490 99508 381106
rect 93600 380430 93778 380490
rect 95912 380430 95986 380490
rect 96048 380430 96170 380490
rect 97000 380430 97090 380490
rect 98088 380430 98194 380490
rect 98496 380430 98562 380490
rect 93350 379405 93410 380430
rect 90771 379404 90837 379405
rect 90771 379340 90772 379404
rect 90836 379340 90837 379404
rect 90771 379339 90837 379340
rect 91323 379404 91389 379405
rect 91323 379340 91324 379404
rect 91388 379340 91389 379404
rect 91323 379339 91389 379340
rect 92427 379404 92493 379405
rect 92427 379340 92428 379404
rect 92492 379340 92493 379404
rect 92427 379339 92493 379340
rect 93347 379404 93413 379405
rect 93347 379340 93348 379404
rect 93412 379340 93413 379404
rect 93347 379339 93413 379340
rect 93718 379269 93778 380430
rect 95926 380357 95986 380430
rect 95923 380356 95989 380357
rect 95923 380292 95924 380356
rect 95988 380292 95989 380356
rect 95923 380291 95989 380292
rect 96110 379405 96170 380430
rect 96107 379404 96173 379405
rect 96107 379340 96108 379404
rect 96172 379340 96173 379404
rect 96107 379339 96173 379340
rect 90035 379268 90101 379269
rect 90035 379204 90036 379268
rect 90100 379204 90101 379268
rect 90035 379203 90101 379204
rect 93715 379268 93781 379269
rect 93715 379204 93716 379268
rect 93780 379204 93781 379268
rect 93715 379203 93781 379204
rect 87643 378180 87709 378181
rect 87643 378116 87644 378180
rect 87708 378116 87709 378180
rect 87643 378115 87709 378116
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 359308 85574 374058
rect 91794 364394 92414 379000
rect 91794 364158 91826 364394
rect 92062 364158 92146 364394
rect 92382 364158 92414 364394
rect 91794 364074 92414 364158
rect 91794 363838 91826 364074
rect 92062 363838 92146 364074
rect 92382 363838 92414 364074
rect 91794 359308 92414 363838
rect 95514 368114 96134 379000
rect 97030 378589 97090 380430
rect 98134 378589 98194 380430
rect 98502 379405 98562 380430
rect 99422 380430 99508 380490
rect 100672 380490 100732 381106
rect 101080 380490 101140 381106
rect 100672 380430 100770 380490
rect 98499 379404 98565 379405
rect 98499 379340 98500 379404
rect 98564 379340 98565 379404
rect 98499 379339 98565 379340
rect 99422 379269 99482 380430
rect 99419 379268 99485 379269
rect 99419 379204 99420 379268
rect 99484 379204 99485 379268
rect 99419 379203 99485 379204
rect 97027 378588 97093 378589
rect 97027 378524 97028 378588
rect 97092 378524 97093 378588
rect 97027 378523 97093 378524
rect 98131 378588 98197 378589
rect 98131 378524 98132 378588
rect 98196 378524 98197 378588
rect 98131 378523 98197 378524
rect 95514 367878 95546 368114
rect 95782 367878 95866 368114
rect 96102 367878 96134 368114
rect 95514 367794 96134 367878
rect 95514 367558 95546 367794
rect 95782 367558 95866 367794
rect 96102 367558 96134 367794
rect 95514 359308 96134 367558
rect 99234 369954 99854 379000
rect 100710 378317 100770 380430
rect 101078 380430 101140 380490
rect 101760 380490 101820 381106
rect 102848 380490 102908 381106
rect 103528 380490 103588 381106
rect 101760 380430 101874 380490
rect 102848 380430 102978 380490
rect 101078 379405 101138 380430
rect 101075 379404 101141 379405
rect 101075 379340 101076 379404
rect 101140 379340 101141 379404
rect 101075 379339 101141 379340
rect 101814 378589 101874 380430
rect 102918 379269 102978 380430
rect 103286 380430 103588 380490
rect 103936 380490 103996 381106
rect 105296 380490 105356 381106
rect 105976 380490 106036 381106
rect 103936 380430 104082 380490
rect 105296 380430 105370 380490
rect 103286 379405 103346 380430
rect 103283 379404 103349 379405
rect 103283 379340 103284 379404
rect 103348 379340 103349 379404
rect 103283 379339 103349 379340
rect 104022 379269 104082 380430
rect 102915 379268 102981 379269
rect 102915 379204 102916 379268
rect 102980 379204 102981 379268
rect 102915 379203 102981 379204
rect 104019 379268 104085 379269
rect 104019 379204 104020 379268
rect 104084 379204 104085 379268
rect 104019 379203 104085 379204
rect 101811 378588 101877 378589
rect 101811 378524 101812 378588
rect 101876 378524 101877 378588
rect 101811 378523 101877 378524
rect 100707 378316 100773 378317
rect 100707 378252 100708 378316
rect 100772 378252 100773 378316
rect 100707 378251 100773 378252
rect 99234 369718 99266 369954
rect 99502 369718 99586 369954
rect 99822 369718 99854 369954
rect 99234 369634 99854 369718
rect 99234 369398 99266 369634
rect 99502 369398 99586 369634
rect 99822 369398 99854 369634
rect 99234 359308 99854 369398
rect 102954 373674 103574 379000
rect 105310 378045 105370 380430
rect 105862 380430 106036 380490
rect 106384 380490 106444 381106
rect 107608 380490 107668 381106
rect 108288 380490 108348 381106
rect 106384 380430 106474 380490
rect 105862 379405 105922 380430
rect 105859 379404 105925 379405
rect 105859 379340 105860 379404
rect 105924 379340 105925 379404
rect 105859 379339 105925 379340
rect 105307 378044 105373 378045
rect 105307 377980 105308 378044
rect 105372 377980 105373 378044
rect 105307 377979 105373 377980
rect 106414 377909 106474 380430
rect 107518 380430 107668 380490
rect 108254 380430 108348 380490
rect 108696 380490 108756 381106
rect 109784 380490 109844 381106
rect 108696 380430 108866 380490
rect 107518 378589 107578 380430
rect 108254 379405 108314 380430
rect 108806 379405 108866 380430
rect 109726 380430 109844 380490
rect 111008 380490 111068 381106
rect 111144 380490 111204 381106
rect 112232 380490 112292 381106
rect 113320 380490 113380 381106
rect 113592 380490 113652 381106
rect 111008 380430 111074 380490
rect 111144 380430 111258 380490
rect 112232 380430 112362 380490
rect 113320 380430 113466 380490
rect 109726 379405 109786 380430
rect 111014 380357 111074 380430
rect 111011 380356 111077 380357
rect 111011 380292 111012 380356
rect 111076 380292 111077 380356
rect 111011 380291 111077 380292
rect 111198 379405 111258 380430
rect 112302 379405 112362 380430
rect 113406 379405 113466 380430
rect 113590 380430 113652 380490
rect 114408 380490 114468 381106
rect 115768 380490 115828 381106
rect 116040 380490 116100 381106
rect 114408 380430 114570 380490
rect 115768 380430 115858 380490
rect 113590 380357 113650 380430
rect 113587 380356 113653 380357
rect 113587 380292 113588 380356
rect 113652 380292 113653 380356
rect 113587 380291 113653 380292
rect 114510 379405 114570 380430
rect 115798 379405 115858 380430
rect 115982 380430 116100 380490
rect 116992 380490 117052 381106
rect 118080 380490 118140 381106
rect 118488 380490 118548 381106
rect 119168 380490 119228 381106
rect 116992 380430 117146 380490
rect 118080 380430 118250 380490
rect 115982 380357 116042 380430
rect 115979 380356 116045 380357
rect 115979 380292 115980 380356
rect 116044 380292 116045 380356
rect 115979 380291 116045 380292
rect 117086 379405 117146 380430
rect 108251 379404 108317 379405
rect 108251 379340 108252 379404
rect 108316 379340 108317 379404
rect 108251 379339 108317 379340
rect 108803 379404 108869 379405
rect 108803 379340 108804 379404
rect 108868 379340 108869 379404
rect 108803 379339 108869 379340
rect 109723 379404 109789 379405
rect 109723 379340 109724 379404
rect 109788 379340 109789 379404
rect 109723 379339 109789 379340
rect 111195 379404 111261 379405
rect 111195 379340 111196 379404
rect 111260 379340 111261 379404
rect 111195 379339 111261 379340
rect 112299 379404 112365 379405
rect 112299 379340 112300 379404
rect 112364 379340 112365 379404
rect 112299 379339 112365 379340
rect 113403 379404 113469 379405
rect 113403 379340 113404 379404
rect 113468 379340 113469 379404
rect 113403 379339 113469 379340
rect 114507 379404 114573 379405
rect 114507 379340 114508 379404
rect 114572 379340 114573 379404
rect 114507 379339 114573 379340
rect 115795 379404 115861 379405
rect 115795 379340 115796 379404
rect 115860 379340 115861 379404
rect 115795 379339 115861 379340
rect 117083 379404 117149 379405
rect 117083 379340 117084 379404
rect 117148 379340 117149 379404
rect 117083 379339 117149 379340
rect 118190 379269 118250 380430
rect 118374 380430 118548 380490
rect 119110 380430 119228 380490
rect 120936 380490 120996 381106
rect 123520 380490 123580 381106
rect 125968 380490 126028 381106
rect 120936 380430 121010 380490
rect 123520 380430 123586 380490
rect 118374 380357 118434 380430
rect 118371 380356 118437 380357
rect 118371 380292 118372 380356
rect 118436 380292 118437 380356
rect 118371 380291 118437 380292
rect 118187 379268 118253 379269
rect 118187 379204 118188 379268
rect 118252 379204 118253 379268
rect 118187 379203 118253 379204
rect 107515 378588 107581 378589
rect 107515 378524 107516 378588
rect 107580 378524 107581 378588
rect 107515 378523 107581 378524
rect 106411 377908 106477 377909
rect 106411 377844 106412 377908
rect 106476 377844 106477 377908
rect 106411 377843 106477 377844
rect 102954 373438 102986 373674
rect 103222 373438 103306 373674
rect 103542 373438 103574 373674
rect 102954 373354 103574 373438
rect 102954 373118 102986 373354
rect 103222 373118 103306 373354
rect 103542 373118 103574 373354
rect 102954 359308 103574 373118
rect 109794 363454 110414 379000
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 359308 110414 362898
rect 113514 367174 114134 379000
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 359308 114134 366618
rect 117234 370894 117854 379000
rect 119110 378589 119170 380430
rect 120950 380357 121010 380430
rect 123526 380357 123586 380430
rect 125918 380430 126028 380490
rect 128280 380490 128340 381106
rect 131000 380490 131060 381106
rect 133448 380490 133508 381106
rect 135896 380490 135956 381106
rect 138480 380490 138540 381106
rect 128280 380430 128370 380490
rect 131000 380430 131130 380490
rect 133448 380430 133522 380490
rect 120947 380356 121013 380357
rect 120947 380292 120948 380356
rect 121012 380292 121013 380356
rect 120947 380291 121013 380292
rect 123523 380356 123589 380357
rect 123523 380292 123524 380356
rect 123588 380292 123589 380356
rect 123523 380291 123589 380292
rect 119107 378588 119173 378589
rect 119107 378524 119108 378588
rect 119172 378524 119173 378588
rect 119107 378523 119173 378524
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 359308 117854 370338
rect 120954 374614 121574 379000
rect 125918 378453 125978 380430
rect 128310 380357 128370 380430
rect 128307 380356 128373 380357
rect 128307 380292 128308 380356
rect 128372 380292 128373 380356
rect 128307 380291 128373 380292
rect 125915 378452 125981 378453
rect 125915 378388 125916 378452
rect 125980 378388 125981 378452
rect 125915 378387 125981 378388
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 359308 121574 374058
rect 127794 364394 128414 379000
rect 131070 378453 131130 380430
rect 131067 378452 131133 378453
rect 131067 378388 131068 378452
rect 131132 378388 131133 378452
rect 131067 378387 131133 378388
rect 127794 364158 127826 364394
rect 128062 364158 128146 364394
rect 128382 364158 128414 364394
rect 127794 364074 128414 364158
rect 127794 363838 127826 364074
rect 128062 363838 128146 364074
rect 128382 363838 128414 364074
rect 127794 359308 128414 363838
rect 131514 368114 132134 379000
rect 133462 378453 133522 380430
rect 135854 380430 135956 380490
rect 138430 380430 138540 380490
rect 140928 380490 140988 381106
rect 143512 380490 143572 381106
rect 145960 380490 146020 381106
rect 148544 380490 148604 381106
rect 150992 380490 151052 381106
rect 140928 380430 141066 380490
rect 143512 380430 143642 380490
rect 145960 380430 146034 380490
rect 148544 380430 148610 380490
rect 135854 380357 135914 380430
rect 135851 380356 135917 380357
rect 135851 380292 135852 380356
rect 135916 380292 135917 380356
rect 135851 380291 135917 380292
rect 133459 378452 133525 378453
rect 133459 378388 133460 378452
rect 133524 378388 133525 378452
rect 133459 378387 133525 378388
rect 131514 367878 131546 368114
rect 131782 367878 131866 368114
rect 132102 367878 132134 368114
rect 131514 367794 132134 367878
rect 131514 367558 131546 367794
rect 131782 367558 131866 367794
rect 132102 367558 132134 367794
rect 131514 359308 132134 367558
rect 135234 369954 135854 379000
rect 138430 378453 138490 380430
rect 141006 379405 141066 380430
rect 143582 380357 143642 380430
rect 143579 380356 143645 380357
rect 143579 380292 143580 380356
rect 143644 380292 143645 380356
rect 143579 380291 143645 380292
rect 145974 379405 146034 380430
rect 148550 380357 148610 380430
rect 150942 380430 151052 380490
rect 153440 380490 153500 381106
rect 155888 380490 155948 381106
rect 158472 380490 158532 381106
rect 160920 380490 160980 381106
rect 153440 380430 153578 380490
rect 155888 380430 155970 380490
rect 158472 380430 158546 380490
rect 148547 380356 148613 380357
rect 148547 380292 148548 380356
rect 148612 380292 148613 380356
rect 148547 380291 148613 380292
rect 150942 379405 151002 380430
rect 153518 379405 153578 380430
rect 155910 380357 155970 380430
rect 158486 380357 158546 380430
rect 160878 380430 160980 380490
rect 163368 380490 163428 381106
rect 165952 380490 166012 381106
rect 183224 380490 183284 381106
rect 163368 380430 163514 380490
rect 165952 380430 166090 380490
rect 160878 380357 160938 380430
rect 163454 380357 163514 380430
rect 166030 380357 166090 380430
rect 183142 380430 183284 380490
rect 183360 380490 183420 381106
rect 183360 380430 183570 380490
rect 155907 380356 155973 380357
rect 155907 380292 155908 380356
rect 155972 380292 155973 380356
rect 155907 380291 155973 380292
rect 158483 380356 158549 380357
rect 158483 380292 158484 380356
rect 158548 380292 158549 380356
rect 158483 380291 158549 380292
rect 160875 380356 160941 380357
rect 160875 380292 160876 380356
rect 160940 380292 160941 380356
rect 160875 380291 160941 380292
rect 163451 380356 163517 380357
rect 163451 380292 163452 380356
rect 163516 380292 163517 380356
rect 163451 380291 163517 380292
rect 166027 380356 166093 380357
rect 166027 380292 166028 380356
rect 166092 380292 166093 380356
rect 166027 380291 166093 380292
rect 141003 379404 141069 379405
rect 141003 379340 141004 379404
rect 141068 379340 141069 379404
rect 141003 379339 141069 379340
rect 145971 379404 146037 379405
rect 145971 379340 145972 379404
rect 146036 379340 146037 379404
rect 145971 379339 146037 379340
rect 150939 379404 151005 379405
rect 150939 379340 150940 379404
rect 151004 379340 151005 379404
rect 150939 379339 151005 379340
rect 153515 379404 153581 379405
rect 153515 379340 153516 379404
rect 153580 379340 153581 379404
rect 153515 379339 153581 379340
rect 138427 378452 138493 378453
rect 138427 378388 138428 378452
rect 138492 378388 138493 378452
rect 138427 378387 138493 378388
rect 135234 369718 135266 369954
rect 135502 369718 135586 369954
rect 135822 369718 135854 369954
rect 135234 369634 135854 369718
rect 135234 369398 135266 369634
rect 135502 369398 135586 369634
rect 135822 369398 135854 369634
rect 135234 359308 135854 369398
rect 138954 373674 139574 379000
rect 138954 373438 138986 373674
rect 139222 373438 139306 373674
rect 139542 373438 139574 373674
rect 138954 373354 139574 373438
rect 138954 373118 138986 373354
rect 139222 373118 139306 373354
rect 139542 373118 139574 373354
rect 138954 359308 139574 373118
rect 145794 363454 146414 379000
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 359308 146414 362898
rect 149514 367174 150134 379000
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 359308 150134 366618
rect 153234 370894 153854 379000
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 359308 153854 370338
rect 156954 374614 157574 379000
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 359308 157574 374058
rect 163794 364394 164414 379000
rect 163794 364158 163826 364394
rect 164062 364158 164146 364394
rect 164382 364158 164414 364394
rect 163794 364074 164414 364158
rect 163794 363838 163826 364074
rect 164062 363838 164146 364074
rect 164382 363838 164414 364074
rect 163794 359308 164414 363838
rect 167514 368114 168134 379000
rect 167514 367878 167546 368114
rect 167782 367878 167866 368114
rect 168102 367878 168134 368114
rect 167514 367794 168134 367878
rect 167514 367558 167546 367794
rect 167782 367558 167866 367794
rect 168102 367558 168134 367794
rect 167514 359308 168134 367558
rect 171234 369954 171854 379000
rect 171234 369718 171266 369954
rect 171502 369718 171586 369954
rect 171822 369718 171854 369954
rect 171234 369634 171854 369718
rect 171234 369398 171266 369634
rect 171502 369398 171586 369634
rect 171822 369398 171854 369634
rect 171234 359308 171854 369398
rect 174954 373674 175574 379000
rect 174954 373438 174986 373674
rect 175222 373438 175306 373674
rect 175542 373438 175574 373674
rect 174954 373354 175574 373438
rect 174954 373118 174986 373354
rect 175222 373118 175306 373354
rect 175542 373118 175574 373354
rect 174954 359308 175574 373118
rect 181794 363454 182414 379000
rect 183142 378317 183202 380430
rect 183510 378453 183570 380430
rect 183507 378452 183573 378453
rect 183507 378388 183508 378452
rect 183572 378388 183573 378452
rect 183507 378387 183573 378388
rect 183139 378316 183205 378317
rect 183139 378252 183140 378316
rect 183204 378252 183205 378316
rect 183139 378251 183205 378252
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 359308 182414 362898
rect 185514 367174 186134 379000
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 359308 186134 366618
rect 189234 370894 189854 379000
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 359308 189854 370338
rect 192954 374614 193574 379000
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 359308 193574 374058
rect 178539 358868 178605 358869
rect 178539 358804 178540 358868
rect 178604 358804 178605 358868
rect 178539 358803 178605 358804
rect 179643 358868 179709 358869
rect 179643 358804 179644 358868
rect 179708 358804 179709 358868
rect 179643 358803 179709 358804
rect 190867 358868 190933 358869
rect 190867 358804 190868 358868
rect 190932 358804 190933 358868
rect 190867 358803 190933 358804
rect 59862 358670 60290 358730
rect 59862 272370 59922 358670
rect 178542 358050 178602 358803
rect 178464 357990 178602 358050
rect 179646 358050 179706 358803
rect 190870 358050 190930 358803
rect 179646 357990 179748 358050
rect 178464 357202 178524 357990
rect 179688 357202 179748 357990
rect 190840 357990 190930 358050
rect 190840 357202 190900 357990
rect 60272 345454 60620 345486
rect 60272 345218 60328 345454
rect 60564 345218 60620 345454
rect 60272 345134 60620 345218
rect 60272 344898 60328 345134
rect 60564 344898 60620 345134
rect 60272 344866 60620 344898
rect 196000 345454 196348 345486
rect 196000 345218 196056 345454
rect 196292 345218 196348 345454
rect 196000 345134 196348 345218
rect 196000 344898 196056 345134
rect 196292 344898 196348 345134
rect 196000 344866 196348 344898
rect 60952 327454 61300 327486
rect 60952 327218 61008 327454
rect 61244 327218 61300 327454
rect 60952 327134 61300 327218
rect 60952 326898 61008 327134
rect 61244 326898 61300 327134
rect 60952 326866 61300 326898
rect 195320 327454 195668 327486
rect 195320 327218 195376 327454
rect 195612 327218 195668 327454
rect 195320 327134 195668 327218
rect 195320 326898 195376 327134
rect 195612 326898 195668 327134
rect 195320 326866 195668 326898
rect 60272 309454 60620 309486
rect 60272 309218 60328 309454
rect 60564 309218 60620 309454
rect 60272 309134 60620 309218
rect 60272 308898 60328 309134
rect 60564 308898 60620 309134
rect 60272 308866 60620 308898
rect 196000 309454 196348 309486
rect 196000 309218 196056 309454
rect 196292 309218 196348 309454
rect 196000 309134 196348 309218
rect 196000 308898 196056 309134
rect 196292 308898 196348 309134
rect 196000 308866 196348 308898
rect 60952 291454 61300 291486
rect 60952 291218 61008 291454
rect 61244 291218 61300 291454
rect 60952 291134 61300 291218
rect 60952 290898 61008 291134
rect 61244 290898 61300 291134
rect 60952 290866 61300 290898
rect 195320 291454 195668 291486
rect 195320 291218 195376 291454
rect 195612 291218 195668 291454
rect 195320 291134 195668 291218
rect 195320 290898 195376 291134
rect 195612 290898 195668 291134
rect 195320 290866 195668 290898
rect 76056 273730 76116 274040
rect 76054 273670 76116 273730
rect 77144 273730 77204 274040
rect 78232 273730 78292 274040
rect 79592 273730 79652 274040
rect 80544 273730 80604 274040
rect 77144 273670 77218 273730
rect 78232 273670 78322 273730
rect 59862 272310 60290 272370
rect 59514 260114 60134 272000
rect 59514 259878 59546 260114
rect 59782 259878 59866 260114
rect 60102 259878 60134 260114
rect 59514 259794 60134 259878
rect 59514 259558 59546 259794
rect 59782 259558 59866 259794
rect 60102 259558 60134 259794
rect 59514 252308 60134 259558
rect 60230 251970 60290 272310
rect 63234 261954 63854 272000
rect 63234 261718 63266 261954
rect 63502 261718 63586 261954
rect 63822 261718 63854 261954
rect 63234 261634 63854 261718
rect 63234 261398 63266 261634
rect 63502 261398 63586 261634
rect 63822 261398 63854 261634
rect 63234 252308 63854 261398
rect 66954 265674 67574 272000
rect 66954 265438 66986 265674
rect 67222 265438 67306 265674
rect 67542 265438 67574 265674
rect 66954 265354 67574 265438
rect 66954 265118 66986 265354
rect 67222 265118 67306 265354
rect 67542 265118 67574 265354
rect 66954 252308 67574 265118
rect 73794 255454 74414 272000
rect 76054 271829 76114 273670
rect 77158 273189 77218 273670
rect 77155 273188 77221 273189
rect 77155 273124 77156 273188
rect 77220 273124 77221 273188
rect 77155 273123 77221 273124
rect 76051 271828 76117 271829
rect 76051 271764 76052 271828
rect 76116 271764 76117 271828
rect 76051 271763 76117 271764
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 252308 74414 254898
rect 77514 259174 78134 272000
rect 78262 271421 78322 273670
rect 79550 273670 79652 273730
rect 80470 273670 80604 273730
rect 81768 273730 81828 274040
rect 83128 273730 83188 274040
rect 84216 273730 84276 274040
rect 85440 273730 85500 274040
rect 81768 273670 82002 273730
rect 78259 271420 78325 271421
rect 78259 271356 78260 271420
rect 78324 271356 78325 271420
rect 78259 271355 78325 271356
rect 79550 271013 79610 273670
rect 80470 271693 80530 273670
rect 80467 271692 80533 271693
rect 80467 271628 80468 271692
rect 80532 271628 80533 271692
rect 80467 271627 80533 271628
rect 79547 271012 79613 271013
rect 79547 270948 79548 271012
rect 79612 270948 79613 271012
rect 79547 270947 79613 270948
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 252308 78134 258618
rect 81234 262894 81854 272000
rect 81942 271285 82002 273670
rect 83046 273670 83188 273730
rect 83966 273670 84276 273730
rect 85438 273670 85500 273730
rect 86528 273730 86588 274040
rect 87616 273730 87676 274040
rect 88296 273730 88356 274040
rect 88704 273730 88764 274040
rect 90064 273730 90124 274040
rect 86528 273670 86602 273730
rect 87616 273670 87706 273730
rect 88296 273670 88442 273730
rect 88704 273670 88810 273730
rect 83046 272373 83106 273670
rect 83043 272372 83109 272373
rect 83043 272308 83044 272372
rect 83108 272308 83109 272372
rect 83043 272307 83109 272308
rect 83966 271829 84026 273670
rect 85438 272237 85498 273670
rect 85435 272236 85501 272237
rect 85435 272172 85436 272236
rect 85500 272172 85501 272236
rect 85435 272171 85501 272172
rect 83963 271828 84029 271829
rect 83963 271764 83964 271828
rect 84028 271764 84029 271828
rect 83963 271763 84029 271764
rect 81939 271284 82005 271285
rect 81939 271220 81940 271284
rect 82004 271220 82005 271284
rect 81939 271219 82005 271220
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 252308 81854 262338
rect 84954 266614 85574 272000
rect 86542 270741 86602 273670
rect 86539 270740 86605 270741
rect 86539 270676 86540 270740
rect 86604 270676 86605 270740
rect 86539 270675 86605 270676
rect 87646 270605 87706 273670
rect 88382 273189 88442 273670
rect 88379 273188 88445 273189
rect 88379 273124 88380 273188
rect 88444 273124 88445 273188
rect 88379 273123 88445 273124
rect 88750 271829 88810 273670
rect 90038 273670 90124 273730
rect 90744 273730 90804 274040
rect 91288 273730 91348 274040
rect 92376 273730 92436 274040
rect 93464 273730 93524 274040
rect 90744 273670 90834 273730
rect 91288 273670 91386 273730
rect 88747 271828 88813 271829
rect 88747 271764 88748 271828
rect 88812 271764 88813 271828
rect 88747 271763 88813 271764
rect 90038 270741 90098 273670
rect 90774 273189 90834 273670
rect 90771 273188 90837 273189
rect 90771 273124 90772 273188
rect 90836 273124 90837 273188
rect 90771 273123 90837 273124
rect 90035 270740 90101 270741
rect 90035 270676 90036 270740
rect 90100 270676 90101 270740
rect 90035 270675 90101 270676
rect 91326 270605 91386 273670
rect 91510 273670 92436 273730
rect 93350 273670 93524 273730
rect 93600 273730 93660 274040
rect 94552 273730 94612 274040
rect 95912 273869 95972 274040
rect 95909 273868 95975 273869
rect 95909 273804 95910 273868
rect 95974 273804 95975 273868
rect 95909 273803 95975 273804
rect 96048 273730 96108 274040
rect 93600 273670 93778 273730
rect 91510 271421 91570 273670
rect 91507 271420 91573 271421
rect 91507 271356 91508 271420
rect 91572 271356 91573 271420
rect 91507 271355 91573 271356
rect 87643 270604 87709 270605
rect 87643 270540 87644 270604
rect 87708 270540 87709 270604
rect 87643 270539 87709 270540
rect 91323 270604 91389 270605
rect 91323 270540 91324 270604
rect 91388 270540 91389 270604
rect 91323 270539 91389 270540
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 252308 85574 266058
rect 91794 256394 92414 272000
rect 93350 270741 93410 273670
rect 93718 273189 93778 273670
rect 94454 273670 94612 273730
rect 95926 273670 96108 273730
rect 97000 273730 97060 274040
rect 98088 273730 98148 274040
rect 98496 273730 98556 274040
rect 99448 273730 99508 274040
rect 97000 273670 97090 273730
rect 98088 273670 98194 273730
rect 98496 273670 98562 273730
rect 93715 273188 93781 273189
rect 93715 273124 93716 273188
rect 93780 273124 93781 273188
rect 93715 273123 93781 273124
rect 94454 271829 94514 273670
rect 95926 272781 95986 273670
rect 95923 272780 95989 272781
rect 95923 272716 95924 272780
rect 95988 272716 95989 272780
rect 95923 272715 95989 272716
rect 94451 271828 94517 271829
rect 94451 271764 94452 271828
rect 94516 271764 94517 271828
rect 94451 271763 94517 271764
rect 93347 270740 93413 270741
rect 93347 270676 93348 270740
rect 93412 270676 93413 270740
rect 93347 270675 93413 270676
rect 91794 256158 91826 256394
rect 92062 256158 92146 256394
rect 92382 256158 92414 256394
rect 91794 256074 92414 256158
rect 91794 255838 91826 256074
rect 92062 255838 92146 256074
rect 92382 255838 92414 256074
rect 91794 252308 92414 255838
rect 95514 260114 96134 272000
rect 97030 270877 97090 273670
rect 98134 273189 98194 273670
rect 98131 273188 98197 273189
rect 98131 273124 98132 273188
rect 98196 273124 98197 273188
rect 98131 273123 98197 273124
rect 98502 272917 98562 273670
rect 99422 273670 99508 273730
rect 100672 273730 100732 274040
rect 101080 273730 101140 274040
rect 100672 273670 100770 273730
rect 99422 272917 99482 273670
rect 98499 272916 98565 272917
rect 98499 272852 98500 272916
rect 98564 272852 98565 272916
rect 98499 272851 98565 272852
rect 99419 272916 99485 272917
rect 99419 272852 99420 272916
rect 99484 272852 99485 272916
rect 99419 272851 99485 272852
rect 100710 272781 100770 273670
rect 101078 273670 101140 273730
rect 101760 273730 101820 274040
rect 102848 273730 102908 274040
rect 101760 273670 101874 273730
rect 100707 272780 100773 272781
rect 100707 272716 100708 272780
rect 100772 272716 100773 272780
rect 100707 272715 100773 272716
rect 97027 270876 97093 270877
rect 97027 270812 97028 270876
rect 97092 270812 97093 270876
rect 97027 270811 97093 270812
rect 95514 259878 95546 260114
rect 95782 259878 95866 260114
rect 96102 259878 96134 260114
rect 95514 259794 96134 259878
rect 95514 259558 95546 259794
rect 95782 259558 95866 259794
rect 96102 259558 96134 259794
rect 95514 252308 96134 259558
rect 99234 261954 99854 272000
rect 101078 271557 101138 273670
rect 101814 273189 101874 273670
rect 102734 273670 102908 273730
rect 103528 273730 103588 274040
rect 103936 273730 103996 274040
rect 105296 273730 105356 274040
rect 105976 273730 106036 274040
rect 103528 273670 103714 273730
rect 103936 273670 104082 273730
rect 105296 273670 105370 273730
rect 101811 273188 101877 273189
rect 101811 273124 101812 273188
rect 101876 273124 101877 273188
rect 101811 273123 101877 273124
rect 101814 272373 101874 273123
rect 101811 272372 101877 272373
rect 101811 272308 101812 272372
rect 101876 272308 101877 272372
rect 101811 272307 101877 272308
rect 102734 271829 102794 273670
rect 102731 271828 102797 271829
rect 102731 271764 102732 271828
rect 102796 271764 102797 271828
rect 102731 271763 102797 271764
rect 101075 271556 101141 271557
rect 101075 271492 101076 271556
rect 101140 271492 101141 271556
rect 101075 271491 101141 271492
rect 99234 261718 99266 261954
rect 99502 261718 99586 261954
rect 99822 261718 99854 261954
rect 99234 261634 99854 261718
rect 99234 261398 99266 261634
rect 99502 261398 99586 261634
rect 99822 261398 99854 261634
rect 99234 252308 99854 261398
rect 102954 265674 103574 272000
rect 103654 271690 103714 273670
rect 103835 271692 103901 271693
rect 103835 271690 103836 271692
rect 103654 271630 103836 271690
rect 103835 271628 103836 271630
rect 103900 271628 103901 271692
rect 103835 271627 103901 271628
rect 104022 270605 104082 273670
rect 105310 271013 105370 273670
rect 105862 273670 106036 273730
rect 106384 273730 106444 274040
rect 107608 273730 107668 274040
rect 108288 273730 108348 274040
rect 108696 273730 108756 274040
rect 109784 273730 109844 274040
rect 106384 273670 106474 273730
rect 105862 271421 105922 273670
rect 105859 271420 105925 271421
rect 105859 271356 105860 271420
rect 105924 271356 105925 271420
rect 105859 271355 105925 271356
rect 105307 271012 105373 271013
rect 105307 270948 105308 271012
rect 105372 270948 105373 271012
rect 105307 270947 105373 270948
rect 106414 270605 106474 273670
rect 107518 273670 107668 273730
rect 108254 273670 108348 273730
rect 108622 273670 108756 273730
rect 109542 273670 109844 273730
rect 111008 273730 111068 274040
rect 111144 273730 111204 274040
rect 112232 273730 112292 274040
rect 113320 273730 113380 274040
rect 113592 273730 113652 274040
rect 111008 273670 111074 273730
rect 111144 273670 111258 273730
rect 107518 271285 107578 273670
rect 108254 271829 108314 273670
rect 108251 271828 108317 271829
rect 108251 271764 108252 271828
rect 108316 271764 108317 271828
rect 108251 271763 108317 271764
rect 107515 271284 107581 271285
rect 107515 271220 107516 271284
rect 107580 271220 107581 271284
rect 107515 271219 107581 271220
rect 108622 270605 108682 273670
rect 109542 271149 109602 273670
rect 109539 271148 109605 271149
rect 109539 271084 109540 271148
rect 109604 271084 109605 271148
rect 109539 271083 109605 271084
rect 104019 270604 104085 270605
rect 104019 270540 104020 270604
rect 104084 270540 104085 270604
rect 104019 270539 104085 270540
rect 106411 270604 106477 270605
rect 106411 270540 106412 270604
rect 106476 270540 106477 270604
rect 106411 270539 106477 270540
rect 108619 270604 108685 270605
rect 108619 270540 108620 270604
rect 108684 270540 108685 270604
rect 108619 270539 108685 270540
rect 102954 265438 102986 265674
rect 103222 265438 103306 265674
rect 103542 265438 103574 265674
rect 102954 265354 103574 265438
rect 102954 265118 102986 265354
rect 103222 265118 103306 265354
rect 103542 265118 103574 265354
rect 102954 252308 103574 265118
rect 109794 255454 110414 272000
rect 111014 271693 111074 273670
rect 111011 271692 111077 271693
rect 111011 271628 111012 271692
rect 111076 271628 111077 271692
rect 111011 271627 111077 271628
rect 111198 270605 111258 273670
rect 112118 273670 112292 273730
rect 113222 273670 113380 273730
rect 113590 273670 113652 273730
rect 114408 273730 114468 274040
rect 115768 273730 115828 274040
rect 116040 273730 116100 274040
rect 116992 273730 117052 274040
rect 118080 273730 118140 274040
rect 118488 273730 118548 274040
rect 119168 273730 119228 274040
rect 120936 273730 120996 274040
rect 114408 273670 114570 273730
rect 115768 273670 115858 273730
rect 112118 273053 112178 273670
rect 112115 273052 112181 273053
rect 112115 272988 112116 273052
rect 112180 272988 112181 273052
rect 112115 272987 112181 272988
rect 113222 270605 113282 273670
rect 113590 272237 113650 273670
rect 113587 272236 113653 272237
rect 113587 272172 113588 272236
rect 113652 272172 113653 272236
rect 113587 272171 113653 272172
rect 111195 270604 111261 270605
rect 111195 270540 111196 270604
rect 111260 270540 111261 270604
rect 111195 270539 111261 270540
rect 113219 270604 113285 270605
rect 113219 270540 113220 270604
rect 113284 270540 113285 270604
rect 113219 270539 113285 270540
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 252308 110414 254898
rect 113514 259174 114134 272000
rect 114510 270605 114570 273670
rect 115798 270605 115858 273670
rect 115982 273670 116100 273730
rect 116902 273670 117052 273730
rect 118006 273670 118140 273730
rect 118374 273670 118548 273730
rect 119110 273670 119228 273730
rect 120766 273670 120996 273730
rect 123520 273730 123580 274040
rect 125968 273730 126028 274040
rect 123520 273670 123586 273730
rect 115982 271557 116042 273670
rect 115979 271556 116045 271557
rect 115979 271492 115980 271556
rect 116044 271492 116045 271556
rect 115979 271491 116045 271492
rect 116902 270877 116962 273670
rect 118006 272645 118066 273670
rect 118003 272644 118069 272645
rect 118003 272580 118004 272644
rect 118068 272580 118069 272644
rect 118003 272579 118069 272580
rect 116899 270876 116965 270877
rect 116899 270812 116900 270876
rect 116964 270812 116965 270876
rect 116899 270811 116965 270812
rect 114507 270604 114573 270605
rect 114507 270540 114508 270604
rect 114572 270540 114573 270604
rect 114507 270539 114573 270540
rect 115795 270604 115861 270605
rect 115795 270540 115796 270604
rect 115860 270540 115861 270604
rect 115795 270539 115861 270540
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 252308 114134 258618
rect 117234 262894 117854 272000
rect 118374 271557 118434 273670
rect 119110 272509 119170 273670
rect 119107 272508 119173 272509
rect 119107 272444 119108 272508
rect 119172 272444 119173 272508
rect 119107 272443 119173 272444
rect 120766 271693 120826 273670
rect 120763 271692 120829 271693
rect 120763 271628 120764 271692
rect 120828 271628 120829 271692
rect 120763 271627 120829 271628
rect 118371 271556 118437 271557
rect 118371 271492 118372 271556
rect 118436 271492 118437 271556
rect 118371 271491 118437 271492
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 252308 117854 262338
rect 120954 266614 121574 272000
rect 123526 271693 123586 273670
rect 125918 273670 126028 273730
rect 128280 273730 128340 274040
rect 131000 273733 131060 274040
rect 130997 273732 131063 273733
rect 128280 273670 128738 273730
rect 125918 271829 125978 273670
rect 125915 271828 125981 271829
rect 125915 271764 125916 271828
rect 125980 271764 125981 271828
rect 125915 271763 125981 271764
rect 123523 271692 123589 271693
rect 123523 271628 123524 271692
rect 123588 271628 123589 271692
rect 123523 271627 123589 271628
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 252308 121574 266058
rect 127794 256394 128414 272000
rect 128678 271149 128738 273670
rect 130997 273668 130998 273732
rect 131062 273668 131063 273732
rect 130997 273667 131063 273668
rect 133448 273597 133508 274040
rect 135896 273597 135956 274040
rect 138480 273597 138540 274040
rect 140928 273597 140988 274040
rect 143512 273730 143572 274040
rect 145960 273733 146020 274040
rect 145957 273732 146023 273733
rect 143512 273670 143642 273730
rect 133445 273596 133511 273597
rect 133445 273532 133446 273596
rect 133510 273532 133511 273596
rect 133445 273531 133511 273532
rect 135893 273596 135959 273597
rect 135893 273532 135894 273596
rect 135958 273532 135959 273596
rect 135893 273531 135959 273532
rect 138477 273596 138543 273597
rect 138477 273532 138478 273596
rect 138542 273532 138543 273596
rect 138477 273531 138543 273532
rect 140925 273596 140991 273597
rect 140925 273532 140926 273596
rect 140990 273532 140991 273596
rect 140925 273531 140991 273532
rect 128675 271148 128741 271149
rect 128675 271084 128676 271148
rect 128740 271084 128741 271148
rect 128675 271083 128741 271084
rect 127794 256158 127826 256394
rect 128062 256158 128146 256394
rect 128382 256158 128414 256394
rect 127794 256074 128414 256158
rect 127794 255838 127826 256074
rect 128062 255838 128146 256074
rect 128382 255838 128414 256074
rect 127794 252308 128414 255838
rect 131514 260114 132134 272000
rect 131514 259878 131546 260114
rect 131782 259878 131866 260114
rect 132102 259878 132134 260114
rect 131514 259794 132134 259878
rect 131514 259558 131546 259794
rect 131782 259558 131866 259794
rect 132102 259558 132134 259794
rect 131514 252308 132134 259558
rect 135234 261954 135854 272000
rect 135234 261718 135266 261954
rect 135502 261718 135586 261954
rect 135822 261718 135854 261954
rect 135234 261634 135854 261718
rect 135234 261398 135266 261634
rect 135502 261398 135586 261634
rect 135822 261398 135854 261634
rect 135234 252308 135854 261398
rect 138954 265674 139574 272000
rect 143582 271829 143642 273670
rect 145957 273668 145958 273732
rect 146022 273668 146023 273732
rect 148544 273730 148604 274040
rect 150992 273730 151052 274040
rect 148544 273670 148610 273730
rect 145957 273667 146023 273668
rect 143579 271828 143645 271829
rect 143579 271764 143580 271828
rect 143644 271764 143645 271828
rect 143579 271763 143645 271764
rect 138954 265438 138986 265674
rect 139222 265438 139306 265674
rect 139542 265438 139574 265674
rect 138954 265354 139574 265438
rect 138954 265118 138986 265354
rect 139222 265118 139306 265354
rect 139542 265118 139574 265354
rect 138954 252308 139574 265118
rect 145794 255454 146414 272000
rect 148550 270877 148610 273670
rect 150942 273670 151052 273730
rect 153440 273730 153500 274040
rect 155888 273730 155948 274040
rect 158472 273730 158532 274040
rect 160920 273730 160980 274040
rect 153440 273670 154130 273730
rect 155888 273670 155970 273730
rect 158472 273670 158546 273730
rect 148547 270876 148613 270877
rect 148547 270812 148548 270876
rect 148612 270812 148613 270876
rect 148547 270811 148613 270812
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 252308 146414 254898
rect 149514 259174 150134 272000
rect 150942 271557 151002 273670
rect 150939 271556 151005 271557
rect 150939 271492 150940 271556
rect 151004 271492 151005 271556
rect 150939 271491 151005 271492
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 252308 150134 258618
rect 153234 262894 153854 272000
rect 154070 271829 154130 273670
rect 155910 271829 155970 273670
rect 154067 271828 154133 271829
rect 154067 271764 154068 271828
rect 154132 271764 154133 271828
rect 154067 271763 154133 271764
rect 155907 271828 155973 271829
rect 155907 271764 155908 271828
rect 155972 271764 155973 271828
rect 155907 271763 155973 271764
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 252308 153854 262338
rect 156954 266614 157574 272000
rect 158486 271829 158546 273670
rect 160878 273670 160980 273730
rect 163368 273730 163428 274040
rect 165952 273730 166012 274040
rect 183224 273730 183284 274040
rect 163368 273670 163514 273730
rect 165952 273670 166090 273730
rect 158483 271828 158549 271829
rect 158483 271764 158484 271828
rect 158548 271764 158549 271828
rect 158483 271763 158549 271764
rect 160878 271693 160938 273670
rect 163454 271693 163514 273670
rect 160875 271692 160941 271693
rect 160875 271628 160876 271692
rect 160940 271628 160941 271692
rect 160875 271627 160941 271628
rect 163451 271692 163517 271693
rect 163451 271628 163452 271692
rect 163516 271628 163517 271692
rect 163451 271627 163517 271628
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 252308 157574 266058
rect 163794 256394 164414 272000
rect 166030 271693 166090 273670
rect 183142 273670 183284 273730
rect 183360 273730 183420 274040
rect 183360 273670 183570 273730
rect 166027 271692 166093 271693
rect 166027 271628 166028 271692
rect 166092 271628 166093 271692
rect 166027 271627 166093 271628
rect 163794 256158 163826 256394
rect 164062 256158 164146 256394
rect 164382 256158 164414 256394
rect 163794 256074 164414 256158
rect 163794 255838 163826 256074
rect 164062 255838 164146 256074
rect 164382 255838 164414 256074
rect 163794 252308 164414 255838
rect 167514 260114 168134 272000
rect 167514 259878 167546 260114
rect 167782 259878 167866 260114
rect 168102 259878 168134 260114
rect 167514 259794 168134 259878
rect 167514 259558 167546 259794
rect 167782 259558 167866 259794
rect 168102 259558 168134 259794
rect 167514 252308 168134 259558
rect 171234 261954 171854 272000
rect 171234 261718 171266 261954
rect 171502 261718 171586 261954
rect 171822 261718 171854 261954
rect 171234 261634 171854 261718
rect 171234 261398 171266 261634
rect 171502 261398 171586 261634
rect 171822 261398 171854 261634
rect 171234 252308 171854 261398
rect 174954 265674 175574 272000
rect 174954 265438 174986 265674
rect 175222 265438 175306 265674
rect 175542 265438 175574 265674
rect 174954 265354 175574 265438
rect 174954 265118 174986 265354
rect 175222 265118 175306 265354
rect 175542 265118 175574 265354
rect 174954 252308 175574 265118
rect 181794 255454 182414 272000
rect 183142 271421 183202 273670
rect 183139 271420 183205 271421
rect 183139 271356 183140 271420
rect 183204 271356 183205 271420
rect 183139 271355 183205 271356
rect 183510 271149 183570 273670
rect 196574 272645 196634 490859
rect 197859 490788 197925 490789
rect 197859 490724 197860 490788
rect 197924 490724 197925 490788
rect 197859 490723 197925 490724
rect 196755 474060 196821 474061
rect 196755 473996 196756 474060
rect 196820 473996 196821 474060
rect 196755 473995 196821 473996
rect 196758 273189 196818 473995
rect 196755 273188 196821 273189
rect 196755 273124 196756 273188
rect 196820 273124 196821 273188
rect 196755 273123 196821 273124
rect 196571 272644 196637 272645
rect 196571 272580 196572 272644
rect 196636 272580 196637 272644
rect 196571 272579 196637 272580
rect 183507 271148 183573 271149
rect 183507 271084 183508 271148
rect 183572 271084 183573 271148
rect 183507 271083 183573 271084
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 179643 253332 179709 253333
rect 179643 253268 179644 253332
rect 179708 253268 179709 253332
rect 179643 253267 179709 253268
rect 178539 253196 178605 253197
rect 178539 253132 178540 253196
rect 178604 253132 178605 253196
rect 178539 253131 178605 253132
rect 59862 251910 60290 251970
rect 59862 166290 59922 251910
rect 178542 250610 178602 253131
rect 178464 250550 178602 250610
rect 179646 250610 179706 253267
rect 181794 252308 182414 254898
rect 185514 259174 186134 272000
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 252308 186134 258618
rect 189234 262894 189854 272000
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 252308 189854 262338
rect 192954 266614 193574 272000
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 190867 252652 190933 252653
rect 190867 252588 190868 252652
rect 190932 252588 190933 252652
rect 190867 252587 190933 252588
rect 190870 250610 190930 252587
rect 192954 252308 193574 266058
rect 179646 250550 179748 250610
rect 178464 250240 178524 250550
rect 179688 250240 179748 250550
rect 190840 250550 190930 250610
rect 190840 250240 190900 250550
rect 60272 237454 60620 237486
rect 60272 237218 60328 237454
rect 60564 237218 60620 237454
rect 60272 237134 60620 237218
rect 60272 236898 60328 237134
rect 60564 236898 60620 237134
rect 60272 236866 60620 236898
rect 196000 237454 196348 237486
rect 196000 237218 196056 237454
rect 196292 237218 196348 237454
rect 196000 237134 196348 237218
rect 196000 236898 196056 237134
rect 196292 236898 196348 237134
rect 196000 236866 196348 236898
rect 60952 219454 61300 219486
rect 60952 219218 61008 219454
rect 61244 219218 61300 219454
rect 60952 219134 61300 219218
rect 60952 218898 61008 219134
rect 61244 218898 61300 219134
rect 60952 218866 61300 218898
rect 195320 219454 195668 219486
rect 195320 219218 195376 219454
rect 195612 219218 195668 219454
rect 195320 219134 195668 219218
rect 195320 218898 195376 219134
rect 195612 218898 195668 219134
rect 195320 218866 195668 218898
rect 60272 201454 60620 201486
rect 60272 201218 60328 201454
rect 60564 201218 60620 201454
rect 60272 201134 60620 201218
rect 60272 200898 60328 201134
rect 60564 200898 60620 201134
rect 60272 200866 60620 200898
rect 196000 201454 196348 201486
rect 196000 201218 196056 201454
rect 196292 201218 196348 201454
rect 196000 201134 196348 201218
rect 196000 200898 196056 201134
rect 196292 200898 196348 201134
rect 196000 200866 196348 200898
rect 60952 183454 61300 183486
rect 60952 183218 61008 183454
rect 61244 183218 61300 183454
rect 60952 183134 61300 183218
rect 60952 182898 61008 183134
rect 61244 182898 61300 183134
rect 60952 182866 61300 182898
rect 195320 183454 195668 183486
rect 195320 183218 195376 183454
rect 195612 183218 195668 183454
rect 195320 183134 195668 183218
rect 195320 182898 195376 183134
rect 195612 182898 195668 183134
rect 195320 182866 195668 182898
rect 76056 166290 76116 167106
rect 59862 166230 60290 166290
rect 59514 152114 60134 165000
rect 59514 151878 59546 152114
rect 59782 151878 59866 152114
rect 60102 151878 60134 152114
rect 59514 151794 60134 151878
rect 59514 151558 59546 151794
rect 59782 151558 59866 151794
rect 60102 151558 60134 151794
rect 59514 145308 60134 151558
rect 60230 145210 60290 166230
rect 76054 166230 76116 166290
rect 77144 166290 77204 167106
rect 78232 166290 78292 167106
rect 79592 166290 79652 167106
rect 80544 167010 80604 167106
rect 81768 167010 81828 167106
rect 83128 167010 83188 167106
rect 84216 167010 84276 167106
rect 85440 167010 85500 167106
rect 77144 166230 77218 166290
rect 78232 166230 78322 166290
rect 63234 155834 63854 165000
rect 63234 155598 63266 155834
rect 63502 155598 63586 155834
rect 63822 155598 63854 155834
rect 63234 155514 63854 155598
rect 63234 155278 63266 155514
rect 63502 155278 63586 155514
rect 63822 155278 63854 155514
rect 63234 145308 63854 155278
rect 66954 157674 67574 165000
rect 66954 157438 66986 157674
rect 67222 157438 67306 157674
rect 67542 157438 67574 157674
rect 66954 157354 67574 157438
rect 66954 157118 66986 157354
rect 67222 157118 67306 157354
rect 67542 157118 67574 157354
rect 66954 145308 67574 157118
rect 73794 147454 74414 165000
rect 76054 164253 76114 166230
rect 77158 164389 77218 166230
rect 77155 164388 77221 164389
rect 77155 164324 77156 164388
rect 77220 164324 77221 164388
rect 77155 164323 77221 164324
rect 76051 164252 76117 164253
rect 76051 164188 76052 164252
rect 76116 164188 76117 164252
rect 76051 164187 76117 164188
rect 73794 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 74414 147454
rect 73794 147134 74414 147218
rect 73794 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 74414 147134
rect 73794 145308 74414 146898
rect 77514 151174 78134 165000
rect 78262 164253 78322 166230
rect 79550 166230 79652 166290
rect 80470 166950 80604 167010
rect 81758 166950 81828 167010
rect 83046 166950 83188 167010
rect 84150 166950 84276 167010
rect 85438 166950 85500 167010
rect 86528 167010 86588 167106
rect 87616 167010 87676 167106
rect 88296 167010 88356 167106
rect 88704 167010 88764 167106
rect 90064 167010 90124 167106
rect 86528 166950 86602 167010
rect 87616 166950 87706 167010
rect 88296 166950 88442 167010
rect 88704 166950 88810 167010
rect 79550 164253 79610 166230
rect 80470 164253 80530 166950
rect 81758 165613 81818 166950
rect 81755 165612 81821 165613
rect 81755 165548 81756 165612
rect 81820 165548 81821 165612
rect 81755 165547 81821 165548
rect 78259 164252 78325 164253
rect 78259 164188 78260 164252
rect 78324 164188 78325 164252
rect 78259 164187 78325 164188
rect 79547 164252 79613 164253
rect 79547 164188 79548 164252
rect 79612 164188 79613 164252
rect 79547 164187 79613 164188
rect 80467 164252 80533 164253
rect 80467 164188 80468 164252
rect 80532 164188 80533 164252
rect 80467 164187 80533 164188
rect 77514 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 78134 151174
rect 77514 150854 78134 150938
rect 77514 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 78134 150854
rect 77514 145308 78134 150618
rect 81234 154894 81854 165000
rect 83046 164253 83106 166950
rect 84150 164253 84210 166950
rect 85438 165613 85498 166950
rect 85435 165612 85501 165613
rect 85435 165548 85436 165612
rect 85500 165548 85501 165612
rect 85435 165547 85501 165548
rect 83043 164252 83109 164253
rect 83043 164188 83044 164252
rect 83108 164188 83109 164252
rect 83043 164187 83109 164188
rect 84147 164252 84213 164253
rect 84147 164188 84148 164252
rect 84212 164188 84213 164252
rect 84147 164187 84213 164188
rect 81234 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 81854 154894
rect 81234 154574 81854 154658
rect 81234 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 81854 154574
rect 81234 145308 81854 154338
rect 84954 158614 85574 165000
rect 86542 164253 86602 166950
rect 87646 164253 87706 166950
rect 88382 164797 88442 166950
rect 88379 164796 88445 164797
rect 88379 164732 88380 164796
rect 88444 164732 88445 164796
rect 88379 164731 88445 164732
rect 88750 164253 88810 166950
rect 90038 166950 90124 167010
rect 90744 167010 90804 167106
rect 91288 167010 91348 167106
rect 92376 167010 92436 167106
rect 93464 167010 93524 167106
rect 90744 166950 90834 167010
rect 91288 166950 91386 167010
rect 92376 166950 92490 167010
rect 90038 164253 90098 166950
rect 90774 165613 90834 166950
rect 90771 165612 90837 165613
rect 90771 165548 90772 165612
rect 90836 165548 90837 165612
rect 90771 165547 90837 165548
rect 91326 164253 91386 166950
rect 92430 165613 92490 166950
rect 93350 166950 93524 167010
rect 93600 167010 93660 167106
rect 94552 167010 94612 167106
rect 95912 167010 95972 167106
rect 93600 166950 93778 167010
rect 92427 165612 92493 165613
rect 92427 165548 92428 165612
rect 92492 165548 92493 165612
rect 92427 165547 92493 165548
rect 86539 164252 86605 164253
rect 86539 164188 86540 164252
rect 86604 164188 86605 164252
rect 86539 164187 86605 164188
rect 87643 164252 87709 164253
rect 87643 164188 87644 164252
rect 87708 164188 87709 164252
rect 87643 164187 87709 164188
rect 88747 164252 88813 164253
rect 88747 164188 88748 164252
rect 88812 164188 88813 164252
rect 88747 164187 88813 164188
rect 90035 164252 90101 164253
rect 90035 164188 90036 164252
rect 90100 164188 90101 164252
rect 90035 164187 90101 164188
rect 91323 164252 91389 164253
rect 91323 164188 91324 164252
rect 91388 164188 91389 164252
rect 91323 164187 91389 164188
rect 84954 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 85574 158614
rect 84954 158294 85574 158378
rect 84954 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 85574 158294
rect 84954 145308 85574 158058
rect 91794 148394 92414 165000
rect 93350 164253 93410 166950
rect 93718 165069 93778 166950
rect 94454 166950 94612 167010
rect 95742 166950 95972 167010
rect 96048 167010 96108 167106
rect 97000 167010 97060 167106
rect 98088 167010 98148 167106
rect 98496 167010 98556 167106
rect 99448 167010 99508 167106
rect 96048 166950 96170 167010
rect 97000 166950 97090 167010
rect 98088 166950 98194 167010
rect 98496 166950 98562 167010
rect 93715 165068 93781 165069
rect 93715 165004 93716 165068
rect 93780 165004 93781 165068
rect 93715 165003 93781 165004
rect 94454 164253 94514 166950
rect 95742 165613 95802 166950
rect 96110 166293 96170 166950
rect 96107 166292 96173 166293
rect 96107 166228 96108 166292
rect 96172 166228 96173 166292
rect 96107 166227 96173 166228
rect 95739 165612 95805 165613
rect 95739 165548 95740 165612
rect 95804 165548 95805 165612
rect 95739 165547 95805 165548
rect 93347 164252 93413 164253
rect 93347 164188 93348 164252
rect 93412 164188 93413 164252
rect 93347 164187 93413 164188
rect 94451 164252 94517 164253
rect 94451 164188 94452 164252
rect 94516 164188 94517 164252
rect 94451 164187 94517 164188
rect 91794 148158 91826 148394
rect 92062 148158 92146 148394
rect 92382 148158 92414 148394
rect 91794 148074 92414 148158
rect 91794 147838 91826 148074
rect 92062 147838 92146 148074
rect 92382 147838 92414 148074
rect 91794 145308 92414 147838
rect 95514 152114 96134 165000
rect 97030 164253 97090 166950
rect 98134 164253 98194 166950
rect 98502 166701 98562 166950
rect 99422 166950 99508 167010
rect 100672 167010 100732 167106
rect 101080 167010 101140 167106
rect 100672 166950 100770 167010
rect 98499 166700 98565 166701
rect 98499 166636 98500 166700
rect 98564 166636 98565 166700
rect 98499 166635 98565 166636
rect 99422 165613 99482 166950
rect 99419 165612 99485 165613
rect 99419 165548 99420 165612
rect 99484 165548 99485 165612
rect 99419 165547 99485 165548
rect 97027 164252 97093 164253
rect 97027 164188 97028 164252
rect 97092 164188 97093 164252
rect 97027 164187 97093 164188
rect 98131 164252 98197 164253
rect 98131 164188 98132 164252
rect 98196 164188 98197 164252
rect 98131 164187 98197 164188
rect 95514 151878 95546 152114
rect 95782 151878 95866 152114
rect 96102 151878 96134 152114
rect 95514 151794 96134 151878
rect 95514 151558 95546 151794
rect 95782 151558 95866 151794
rect 96102 151558 96134 151794
rect 95514 145308 96134 151558
rect 99234 155834 99854 165000
rect 100710 164525 100770 166950
rect 101078 166950 101140 167010
rect 101760 167010 101820 167106
rect 102848 167010 102908 167106
rect 103528 167010 103588 167106
rect 103936 167010 103996 167106
rect 101760 166950 101874 167010
rect 101078 166701 101138 166950
rect 101075 166700 101141 166701
rect 101075 166636 101076 166700
rect 101140 166636 101141 166700
rect 101075 166635 101141 166636
rect 100707 164524 100773 164525
rect 100707 164460 100708 164524
rect 100772 164460 100773 164524
rect 100707 164459 100773 164460
rect 101814 164253 101874 166950
rect 102734 166950 102908 167010
rect 103470 166950 103588 167010
rect 103838 166950 103996 167010
rect 105296 167010 105356 167106
rect 105976 167010 106036 167106
rect 105296 166950 105370 167010
rect 102734 164253 102794 166950
rect 103470 165613 103530 166950
rect 103467 165612 103533 165613
rect 103467 165548 103468 165612
rect 103532 165548 103533 165612
rect 103467 165547 103533 165548
rect 101811 164252 101877 164253
rect 101811 164188 101812 164252
rect 101876 164188 101877 164252
rect 101811 164187 101877 164188
rect 102731 164252 102797 164253
rect 102731 164188 102732 164252
rect 102796 164188 102797 164252
rect 102731 164187 102797 164188
rect 99234 155598 99266 155834
rect 99502 155598 99586 155834
rect 99822 155598 99854 155834
rect 99234 155514 99854 155598
rect 99234 155278 99266 155514
rect 99502 155278 99586 155514
rect 99822 155278 99854 155514
rect 99234 145308 99854 155278
rect 102954 157674 103574 165000
rect 103838 164253 103898 166950
rect 105310 164933 105370 166950
rect 105862 166950 106036 167010
rect 106384 167010 106444 167106
rect 107608 167010 107668 167106
rect 108288 167010 108348 167106
rect 108696 167010 108756 167106
rect 106384 166950 106474 167010
rect 105862 166701 105922 166950
rect 105859 166700 105925 166701
rect 105859 166636 105860 166700
rect 105924 166636 105925 166700
rect 105859 166635 105925 166636
rect 106414 164933 106474 166950
rect 107518 166950 107668 167010
rect 108254 166950 108348 167010
rect 108622 166950 108756 167010
rect 105307 164932 105373 164933
rect 105307 164868 105308 164932
rect 105372 164868 105373 164932
rect 105307 164867 105373 164868
rect 106411 164932 106477 164933
rect 106411 164868 106412 164932
rect 106476 164868 106477 164932
rect 106411 164867 106477 164868
rect 107518 164797 107578 166950
rect 108254 166701 108314 166950
rect 108251 166700 108317 166701
rect 108251 166636 108252 166700
rect 108316 166636 108317 166700
rect 108251 166635 108317 166636
rect 107515 164796 107581 164797
rect 107515 164732 107516 164796
rect 107580 164732 107581 164796
rect 107515 164731 107581 164732
rect 108622 164525 108682 166950
rect 109784 166562 109844 167106
rect 109726 166502 109844 166562
rect 111008 166562 111068 167106
rect 111144 166562 111204 167106
rect 112232 166562 112292 167106
rect 113320 166565 113380 167106
rect 111008 166502 111074 166562
rect 111144 166502 111258 166562
rect 109726 165613 109786 166502
rect 111014 165613 111074 166502
rect 111198 165613 111258 166502
rect 112118 166502 112292 166562
rect 113317 166564 113383 166565
rect 112118 165613 112178 166502
rect 113317 166500 113318 166564
rect 113382 166500 113383 166564
rect 113317 166499 113383 166500
rect 113592 166290 113652 167106
rect 113590 166230 113652 166290
rect 114408 166290 114468 167106
rect 115768 166290 115828 167106
rect 116040 166290 116100 167106
rect 116992 166290 117052 167106
rect 118080 166290 118140 167106
rect 118488 166290 118548 167106
rect 119168 166290 119228 167106
rect 114408 166230 114570 166290
rect 115768 166230 115858 166290
rect 113590 165613 113650 166230
rect 109723 165612 109789 165613
rect 109723 165548 109724 165612
rect 109788 165548 109789 165612
rect 109723 165547 109789 165548
rect 111011 165612 111077 165613
rect 111011 165548 111012 165612
rect 111076 165548 111077 165612
rect 111011 165547 111077 165548
rect 111195 165612 111261 165613
rect 111195 165548 111196 165612
rect 111260 165548 111261 165612
rect 111195 165547 111261 165548
rect 112115 165612 112181 165613
rect 112115 165548 112116 165612
rect 112180 165548 112181 165612
rect 112115 165547 112181 165548
rect 113587 165612 113653 165613
rect 113587 165548 113588 165612
rect 113652 165548 113653 165612
rect 113587 165547 113653 165548
rect 108619 164524 108685 164525
rect 108619 164460 108620 164524
rect 108684 164460 108685 164524
rect 108619 164459 108685 164460
rect 103835 164252 103901 164253
rect 103835 164188 103836 164252
rect 103900 164188 103901 164252
rect 103835 164187 103901 164188
rect 102954 157438 102986 157674
rect 103222 157438 103306 157674
rect 103542 157438 103574 157674
rect 102954 157354 103574 157438
rect 102954 157118 102986 157354
rect 103222 157118 103306 157354
rect 103542 157118 103574 157354
rect 102954 145308 103574 157118
rect 109794 147454 110414 165000
rect 109794 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 110414 147454
rect 109794 147134 110414 147218
rect 109794 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 110414 147134
rect 109794 145308 110414 146898
rect 113514 151174 114134 165000
rect 114510 164933 114570 166230
rect 114507 164932 114573 164933
rect 114507 164868 114508 164932
rect 114572 164868 114573 164932
rect 114507 164867 114573 164868
rect 115798 164525 115858 166230
rect 115982 166230 116100 166290
rect 116902 166230 117052 166290
rect 118006 166230 118140 166290
rect 118374 166230 118548 166290
rect 119110 166230 119228 166290
rect 120936 166290 120996 167106
rect 123520 166290 123580 167106
rect 125968 166290 126028 167106
rect 128280 167010 128340 167106
rect 131000 167010 131060 167106
rect 128280 166950 128554 167010
rect 128280 166910 128370 166950
rect 120936 166230 121010 166290
rect 123520 166230 123586 166290
rect 115982 165613 116042 166230
rect 116902 165613 116962 166230
rect 118006 165613 118066 166230
rect 118374 165613 118434 166230
rect 115979 165612 116045 165613
rect 115979 165548 115980 165612
rect 116044 165548 116045 165612
rect 115979 165547 116045 165548
rect 116899 165612 116965 165613
rect 116899 165548 116900 165612
rect 116964 165548 116965 165612
rect 116899 165547 116965 165548
rect 118003 165612 118069 165613
rect 118003 165548 118004 165612
rect 118068 165548 118069 165612
rect 118003 165547 118069 165548
rect 118371 165612 118437 165613
rect 118371 165548 118372 165612
rect 118436 165548 118437 165612
rect 118371 165547 118437 165548
rect 119110 165069 119170 166230
rect 120950 165613 121010 166230
rect 123526 165613 123586 166230
rect 125918 166230 126028 166290
rect 125918 165613 125978 166230
rect 128494 165613 128554 166950
rect 130886 166950 131060 167010
rect 133448 167010 133508 167106
rect 135896 167010 135956 167106
rect 133448 166950 133522 167010
rect 130886 165613 130946 166950
rect 133462 165613 133522 166950
rect 135854 166950 135956 167010
rect 120947 165612 121013 165613
rect 120947 165548 120948 165612
rect 121012 165548 121013 165612
rect 120947 165547 121013 165548
rect 123523 165612 123589 165613
rect 123523 165548 123524 165612
rect 123588 165548 123589 165612
rect 123523 165547 123589 165548
rect 125915 165612 125981 165613
rect 125915 165548 125916 165612
rect 125980 165548 125981 165612
rect 125915 165547 125981 165548
rect 128491 165612 128557 165613
rect 128491 165548 128492 165612
rect 128556 165548 128557 165612
rect 128491 165547 128557 165548
rect 130883 165612 130949 165613
rect 130883 165548 130884 165612
rect 130948 165548 130949 165612
rect 130883 165547 130949 165548
rect 133459 165612 133525 165613
rect 133459 165548 133460 165612
rect 133524 165548 133525 165612
rect 133459 165547 133525 165548
rect 135854 165205 135914 166950
rect 138480 166837 138540 167106
rect 138477 166836 138543 166837
rect 138477 166772 138478 166836
rect 138542 166772 138543 166836
rect 138477 166771 138543 166772
rect 140928 166701 140988 167106
rect 143512 166837 143572 167106
rect 145960 166837 146020 167106
rect 148544 167010 148604 167106
rect 150992 167010 151052 167106
rect 153440 167010 153500 167106
rect 148366 166973 148604 167010
rect 148363 166972 148604 166973
rect 148363 166908 148364 166972
rect 148428 166950 148604 166972
rect 150942 166950 151052 167010
rect 153334 166950 153500 167010
rect 155888 167010 155948 167106
rect 155888 166950 155970 167010
rect 148428 166908 148429 166950
rect 148363 166907 148429 166908
rect 143509 166836 143575 166837
rect 143509 166772 143510 166836
rect 143574 166772 143575 166836
rect 143509 166771 143575 166772
rect 145957 166836 146023 166837
rect 145957 166772 145958 166836
rect 146022 166772 146023 166836
rect 145957 166771 146023 166772
rect 140925 166700 140991 166701
rect 140925 166636 140926 166700
rect 140990 166636 140991 166700
rect 140925 166635 140991 166636
rect 150942 166565 151002 166950
rect 153334 166565 153394 166950
rect 150939 166564 151005 166565
rect 150939 166500 150940 166564
rect 151004 166500 151005 166564
rect 150939 166499 151005 166500
rect 153331 166564 153397 166565
rect 153331 166500 153332 166564
rect 153396 166500 153397 166564
rect 153331 166499 153397 166500
rect 155910 165477 155970 166950
rect 158472 166290 158532 167106
rect 160920 166290 160980 167106
rect 163368 166701 163428 167106
rect 165952 166701 166012 167106
rect 183224 167010 183284 167106
rect 183142 166950 183284 167010
rect 183360 167010 183420 167106
rect 183360 166950 183570 167010
rect 163365 166700 163431 166701
rect 163365 166636 163366 166700
rect 163430 166636 163431 166700
rect 163365 166635 163431 166636
rect 165949 166700 166015 166701
rect 165949 166636 165950 166700
rect 166014 166636 166015 166700
rect 165949 166635 166015 166636
rect 158472 166230 158546 166290
rect 155907 165476 155973 165477
rect 155907 165412 155908 165476
rect 155972 165412 155973 165476
rect 155907 165411 155973 165412
rect 158486 165341 158546 166230
rect 160878 166230 160980 166290
rect 158483 165340 158549 165341
rect 158483 165276 158484 165340
rect 158548 165276 158549 165340
rect 158483 165275 158549 165276
rect 135851 165204 135917 165205
rect 135851 165140 135852 165204
rect 135916 165140 135917 165204
rect 135851 165139 135917 165140
rect 119107 165068 119173 165069
rect 119107 165004 119108 165068
rect 119172 165004 119173 165068
rect 119107 165003 119173 165004
rect 115795 164524 115861 164525
rect 115795 164460 115796 164524
rect 115860 164460 115861 164524
rect 115795 164459 115861 164460
rect 113514 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 114134 151174
rect 113514 150854 114134 150938
rect 113514 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 114134 150854
rect 113514 145308 114134 150618
rect 117234 154894 117854 165000
rect 117234 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 117854 154894
rect 117234 154574 117854 154658
rect 117234 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 117854 154574
rect 117234 145308 117854 154338
rect 120954 158614 121574 165000
rect 120954 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 121574 158614
rect 120954 158294 121574 158378
rect 120954 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 121574 158294
rect 120954 145308 121574 158058
rect 127794 148394 128414 165000
rect 127794 148158 127826 148394
rect 128062 148158 128146 148394
rect 128382 148158 128414 148394
rect 127794 148074 128414 148158
rect 127794 147838 127826 148074
rect 128062 147838 128146 148074
rect 128382 147838 128414 148074
rect 127794 145308 128414 147838
rect 131514 152114 132134 165000
rect 131514 151878 131546 152114
rect 131782 151878 131866 152114
rect 132102 151878 132134 152114
rect 131514 151794 132134 151878
rect 131514 151558 131546 151794
rect 131782 151558 131866 151794
rect 132102 151558 132134 151794
rect 131514 145308 132134 151558
rect 135234 155834 135854 165000
rect 135234 155598 135266 155834
rect 135502 155598 135586 155834
rect 135822 155598 135854 155834
rect 135234 155514 135854 155598
rect 135234 155278 135266 155514
rect 135502 155278 135586 155514
rect 135822 155278 135854 155514
rect 135234 145308 135854 155278
rect 138954 157674 139574 165000
rect 138954 157438 138986 157674
rect 139222 157438 139306 157674
rect 139542 157438 139574 157674
rect 138954 157354 139574 157438
rect 138954 157118 138986 157354
rect 139222 157118 139306 157354
rect 139542 157118 139574 157354
rect 138954 145308 139574 157118
rect 145794 147454 146414 165000
rect 145794 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 146414 147454
rect 145794 147134 146414 147218
rect 145794 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 146414 147134
rect 145794 145308 146414 146898
rect 149514 151174 150134 165000
rect 149514 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 150134 151174
rect 149514 150854 150134 150938
rect 149514 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 150134 150854
rect 149514 145308 150134 150618
rect 153234 154894 153854 165000
rect 153234 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 153854 154894
rect 153234 154574 153854 154658
rect 153234 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 153854 154574
rect 153234 145308 153854 154338
rect 156954 158614 157574 165000
rect 160878 164661 160938 166230
rect 183142 165613 183202 166950
rect 183139 165612 183205 165613
rect 183139 165548 183140 165612
rect 183204 165548 183205 165612
rect 183139 165547 183205 165548
rect 183510 165069 183570 166950
rect 183507 165068 183573 165069
rect 183507 165004 183508 165068
rect 183572 165004 183573 165068
rect 183507 165003 183573 165004
rect 160875 164660 160941 164661
rect 160875 164596 160876 164660
rect 160940 164596 160941 164660
rect 160875 164595 160941 164596
rect 156954 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 157574 158614
rect 156954 158294 157574 158378
rect 156954 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 157574 158294
rect 156954 145308 157574 158058
rect 163794 148394 164414 165000
rect 163794 148158 163826 148394
rect 164062 148158 164146 148394
rect 164382 148158 164414 148394
rect 163794 148074 164414 148158
rect 163794 147838 163826 148074
rect 164062 147838 164146 148074
rect 164382 147838 164414 148074
rect 163794 145308 164414 147838
rect 167514 152114 168134 165000
rect 167514 151878 167546 152114
rect 167782 151878 167866 152114
rect 168102 151878 168134 152114
rect 167514 151794 168134 151878
rect 167514 151558 167546 151794
rect 167782 151558 167866 151794
rect 168102 151558 168134 151794
rect 167514 145308 168134 151558
rect 171234 155834 171854 165000
rect 171234 155598 171266 155834
rect 171502 155598 171586 155834
rect 171822 155598 171854 155834
rect 171234 155514 171854 155598
rect 171234 155278 171266 155514
rect 171502 155278 171586 155514
rect 171822 155278 171854 155514
rect 171234 145308 171854 155278
rect 174954 157674 175574 165000
rect 174954 157438 174986 157674
rect 175222 157438 175306 157674
rect 175542 157438 175574 157674
rect 174954 157354 175574 157438
rect 174954 157118 174986 157354
rect 175222 157118 175306 157354
rect 175542 157118 175574 157354
rect 174954 145308 175574 157118
rect 181794 147454 182414 165000
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 145308 182414 146898
rect 185514 151174 186134 165000
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 145308 186134 150618
rect 189234 154894 189854 165000
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 145308 189854 154338
rect 192954 158614 193574 165000
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 190867 145484 190933 145485
rect 190867 145420 190868 145484
rect 190932 145420 190933 145484
rect 190867 145419 190933 145420
rect 59862 145150 60290 145210
rect 59862 58581 59922 145150
rect 178539 144940 178605 144941
rect 178539 144876 178540 144940
rect 178604 144876 178605 144940
rect 178539 144875 178605 144876
rect 179643 144940 179709 144941
rect 179643 144876 179644 144940
rect 179708 144876 179709 144940
rect 179643 144875 179709 144876
rect 178542 143850 178602 144875
rect 178464 143790 178602 143850
rect 179646 143850 179706 144875
rect 190870 143850 190930 145419
rect 192954 145308 193574 158058
rect 179646 143790 179748 143850
rect 178464 143202 178524 143790
rect 179688 143202 179748 143790
rect 190840 143790 190930 143850
rect 190840 143202 190900 143790
rect 60272 129454 60620 129486
rect 60272 129218 60328 129454
rect 60564 129218 60620 129454
rect 60272 129134 60620 129218
rect 60272 128898 60328 129134
rect 60564 128898 60620 129134
rect 60272 128866 60620 128898
rect 196000 129454 196348 129486
rect 196000 129218 196056 129454
rect 196292 129218 196348 129454
rect 196000 129134 196348 129218
rect 196000 128898 196056 129134
rect 196292 128898 196348 129134
rect 196000 128866 196348 128898
rect 60952 111454 61300 111486
rect 60952 111218 61008 111454
rect 61244 111218 61300 111454
rect 60952 111134 61300 111218
rect 60952 110898 61008 111134
rect 61244 110898 61300 111134
rect 60952 110866 61300 110898
rect 195320 111454 195668 111486
rect 195320 111218 195376 111454
rect 195612 111218 195668 111454
rect 195320 111134 195668 111218
rect 195320 110898 195376 111134
rect 195612 110898 195668 111134
rect 195320 110866 195668 110898
rect 60272 93454 60620 93486
rect 60272 93218 60328 93454
rect 60564 93218 60620 93454
rect 60272 93134 60620 93218
rect 60272 92898 60328 93134
rect 60564 92898 60620 93134
rect 60272 92866 60620 92898
rect 196000 93454 196348 93486
rect 196000 93218 196056 93454
rect 196292 93218 196348 93454
rect 196000 93134 196348 93218
rect 196000 92898 196056 93134
rect 196292 92898 196348 93134
rect 196000 92866 196348 92898
rect 60952 75454 61300 75486
rect 60952 75218 61008 75454
rect 61244 75218 61300 75454
rect 60952 75134 61300 75218
rect 60952 74898 61008 75134
rect 61244 74898 61300 75134
rect 60952 74866 61300 74898
rect 195320 75454 195668 75486
rect 195320 75218 195376 75454
rect 195612 75218 195668 75454
rect 195320 75134 195668 75218
rect 195320 74898 195376 75134
rect 195612 74898 195668 75134
rect 195320 74866 195668 74898
rect 76056 59530 76116 60106
rect 77144 59805 77204 60106
rect 77141 59804 77207 59805
rect 77141 59740 77142 59804
rect 77206 59740 77207 59804
rect 77141 59739 77207 59740
rect 76054 59470 76116 59530
rect 78232 59530 78292 60106
rect 79592 59530 79652 60106
rect 80544 59802 80604 60106
rect 78232 59470 78322 59530
rect 59859 58580 59925 58581
rect 59859 58516 59860 58580
rect 59924 58516 59925 58580
rect 59859 58515 59925 58516
rect 59307 58444 59373 58445
rect 59307 58380 59308 58444
rect 59372 58380 59373 58444
rect 59307 58379 59373 58380
rect 58939 57492 59005 57493
rect 58939 57428 58940 57492
rect 59004 57428 59005 57492
rect 58939 57427 59005 57428
rect 58755 57084 58821 57085
rect 58755 57020 58756 57084
rect 58820 57020 58821 57084
rect 58755 57019 58821 57020
rect 57835 56132 57901 56133
rect 57835 56068 57836 56132
rect 57900 56068 57901 56132
rect 57835 56067 57901 56068
rect 57467 54772 57533 54773
rect 57467 54708 57468 54772
rect 57532 54708 57533 54772
rect 57467 54707 57533 54708
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 25174 60134 58000
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 28894 63854 58000
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 32614 67574 58000
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 39454 74414 58000
rect 76054 57901 76114 59470
rect 76051 57900 76117 57901
rect 76051 57836 76052 57900
rect 76116 57836 76117 57900
rect 76051 57835 76117 57836
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 43174 78134 58000
rect 78262 57901 78322 59470
rect 79550 59470 79652 59530
rect 80470 59742 80604 59802
rect 79550 57901 79610 59470
rect 80470 57901 80530 59742
rect 81768 59530 81828 60106
rect 83128 59805 83188 60106
rect 84216 59805 84276 60106
rect 83125 59804 83191 59805
rect 83125 59740 83126 59804
rect 83190 59740 83191 59804
rect 83125 59739 83191 59740
rect 84213 59804 84279 59805
rect 84213 59740 84214 59804
rect 84278 59740 84279 59804
rect 84213 59739 84279 59740
rect 85440 59530 85500 60106
rect 81768 59470 82002 59530
rect 78259 57900 78325 57901
rect 78259 57836 78260 57900
rect 78324 57836 78325 57900
rect 78259 57835 78325 57836
rect 79547 57900 79613 57901
rect 79547 57836 79548 57900
rect 79612 57836 79613 57900
rect 79547 57835 79613 57836
rect 80467 57900 80533 57901
rect 80467 57836 80468 57900
rect 80532 57836 80533 57900
rect 80467 57835 80533 57836
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 46894 81854 58000
rect 81942 57901 82002 59470
rect 85438 59470 85500 59530
rect 86528 59530 86588 60106
rect 87616 59530 87676 60106
rect 88296 59530 88356 60106
rect 88704 59530 88764 60106
rect 90064 59530 90124 60106
rect 86528 59470 86602 59530
rect 87616 59470 87706 59530
rect 88296 59470 88442 59530
rect 88704 59470 88810 59530
rect 85438 59397 85498 59470
rect 85435 59396 85501 59397
rect 85435 59332 85436 59396
rect 85500 59332 85501 59396
rect 85435 59331 85501 59332
rect 81939 57900 82005 57901
rect 81939 57836 81940 57900
rect 82004 57836 82005 57900
rect 81939 57835 82005 57836
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 50614 85574 58000
rect 86542 57901 86602 59470
rect 87646 57901 87706 59470
rect 86539 57900 86605 57901
rect 86539 57836 86540 57900
rect 86604 57836 86605 57900
rect 86539 57835 86605 57836
rect 87643 57900 87709 57901
rect 87643 57836 87644 57900
rect 87708 57836 87709 57900
rect 87643 57835 87709 57836
rect 88382 57085 88442 59470
rect 88750 57901 88810 59470
rect 90038 59470 90124 59530
rect 90744 59530 90804 60106
rect 91288 59530 91348 60106
rect 92376 59530 92436 60106
rect 93464 59530 93524 60106
rect 90744 59470 90834 59530
rect 91288 59470 91386 59530
rect 90038 57901 90098 59470
rect 90774 57901 90834 59470
rect 91326 57901 91386 59470
rect 92246 59470 92436 59530
rect 93350 59470 93524 59530
rect 93600 59530 93660 60106
rect 94552 59666 94612 60106
rect 94454 59606 94612 59666
rect 95912 59666 95972 60106
rect 95912 59606 95986 59666
rect 93600 59470 93778 59530
rect 92246 58173 92306 59470
rect 92243 58172 92309 58173
rect 92243 58108 92244 58172
rect 92308 58108 92309 58172
rect 92243 58107 92309 58108
rect 88747 57900 88813 57901
rect 88747 57836 88748 57900
rect 88812 57836 88813 57900
rect 88747 57835 88813 57836
rect 90035 57900 90101 57901
rect 90035 57836 90036 57900
rect 90100 57836 90101 57900
rect 90035 57835 90101 57836
rect 90771 57900 90837 57901
rect 90771 57836 90772 57900
rect 90836 57836 90837 57900
rect 90771 57835 90837 57836
rect 91323 57900 91389 57901
rect 91323 57836 91324 57900
rect 91388 57836 91389 57900
rect 91323 57835 91389 57836
rect 91794 57454 92414 58000
rect 93350 57901 93410 59470
rect 93718 57901 93778 59470
rect 94454 57901 94514 59606
rect 95926 59397 95986 59606
rect 96048 59530 96108 60106
rect 97000 59530 97060 60106
rect 98088 59666 98148 60106
rect 98088 59606 98194 59666
rect 96048 59470 96354 59530
rect 97000 59470 97090 59530
rect 95923 59396 95989 59397
rect 95923 59332 95924 59396
rect 95988 59332 95989 59396
rect 95923 59331 95989 59332
rect 93347 57900 93413 57901
rect 93347 57836 93348 57900
rect 93412 57836 93413 57900
rect 93347 57835 93413 57836
rect 93715 57900 93781 57901
rect 93715 57836 93716 57900
rect 93780 57836 93781 57900
rect 93715 57835 93781 57836
rect 94451 57900 94517 57901
rect 94451 57836 94452 57900
rect 94516 57836 94517 57900
rect 94451 57835 94517 57836
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 88379 57084 88445 57085
rect 88379 57020 88380 57084
rect 88444 57020 88445 57084
rect 88379 57019 88445 57020
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 25174 96134 58000
rect 96294 56949 96354 59470
rect 97030 57085 97090 59470
rect 98134 59397 98194 59606
rect 98496 59530 98556 60106
rect 99448 59805 99508 60106
rect 99445 59804 99511 59805
rect 99445 59740 99446 59804
rect 99510 59740 99511 59804
rect 99445 59739 99511 59740
rect 100672 59669 100732 60106
rect 100672 59668 100773 59669
rect 100672 59606 100708 59668
rect 100707 59604 100708 59606
rect 100772 59604 100773 59668
rect 100707 59603 100773 59604
rect 101080 59530 101140 60106
rect 98496 59470 98562 59530
rect 98131 59396 98197 59397
rect 98131 59332 98132 59396
rect 98196 59332 98197 59396
rect 98131 59331 98197 59332
rect 98502 57901 98562 59470
rect 101078 59470 101140 59530
rect 101760 59530 101820 60106
rect 102848 59805 102908 60106
rect 102845 59804 102911 59805
rect 102845 59740 102846 59804
rect 102910 59740 102911 59804
rect 102845 59739 102911 59740
rect 103528 59530 103588 60106
rect 103936 59669 103996 60106
rect 103933 59668 103999 59669
rect 103933 59604 103934 59668
rect 103998 59604 103999 59668
rect 103933 59603 103999 59604
rect 105296 59530 105356 60106
rect 105976 59530 106036 60106
rect 101760 59470 101874 59530
rect 103528 59470 103898 59530
rect 105296 59470 105370 59530
rect 101078 58445 101138 59470
rect 101075 58444 101141 58445
rect 101075 58380 101076 58444
rect 101140 58380 101141 58444
rect 101075 58379 101141 58380
rect 98499 57900 98565 57901
rect 98499 57836 98500 57900
rect 98564 57836 98565 57900
rect 98499 57835 98565 57836
rect 97027 57084 97093 57085
rect 97027 57020 97028 57084
rect 97092 57020 97093 57084
rect 97027 57019 97093 57020
rect 96291 56948 96357 56949
rect 96291 56884 96292 56948
rect 96356 56884 96357 56948
rect 96291 56883 96357 56884
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 28894 99854 58000
rect 101814 57901 101874 59470
rect 101811 57900 101877 57901
rect 101811 57836 101812 57900
rect 101876 57836 101877 57900
rect 101811 57835 101877 57836
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 32614 103574 58000
rect 103838 57357 103898 59470
rect 105310 59397 105370 59470
rect 105862 59470 106036 59530
rect 106384 59530 106444 60106
rect 107608 59805 107668 60106
rect 107605 59804 107671 59805
rect 107605 59740 107606 59804
rect 107670 59740 107671 59804
rect 107605 59739 107671 59740
rect 108288 59530 108348 60106
rect 108696 59530 108756 60106
rect 109784 59530 109844 60106
rect 106384 59470 106474 59530
rect 105307 59396 105373 59397
rect 105307 59332 105308 59396
rect 105372 59332 105373 59396
rect 105307 59331 105373 59332
rect 103835 57356 103901 57357
rect 103835 57292 103836 57356
rect 103900 57292 103901 57356
rect 103835 57291 103901 57292
rect 105862 57221 105922 59470
rect 106414 59397 106474 59470
rect 108254 59470 108348 59530
rect 108622 59470 108756 59530
rect 109542 59470 109844 59530
rect 111008 59530 111068 60106
rect 111144 59530 111204 60106
rect 112232 59530 112292 60106
rect 113320 59530 113380 60106
rect 113592 59530 113652 60106
rect 114408 59669 114468 60106
rect 114405 59668 114471 59669
rect 114405 59604 114406 59668
rect 114470 59604 114471 59668
rect 114405 59603 114471 59604
rect 111008 59470 111074 59530
rect 111144 59470 111258 59530
rect 106411 59396 106477 59397
rect 106411 59332 106412 59396
rect 106476 59332 106477 59396
rect 106411 59331 106477 59332
rect 108254 58717 108314 59470
rect 108251 58716 108317 58717
rect 108251 58652 108252 58716
rect 108316 58652 108317 58716
rect 108251 58651 108317 58652
rect 108622 57901 108682 59470
rect 109542 57901 109602 59470
rect 111014 58853 111074 59470
rect 111011 58852 111077 58853
rect 111011 58788 111012 58852
rect 111076 58788 111077 58852
rect 111011 58787 111077 58788
rect 108619 57900 108685 57901
rect 108619 57836 108620 57900
rect 108684 57836 108685 57900
rect 108619 57835 108685 57836
rect 109539 57900 109605 57901
rect 109539 57836 109540 57900
rect 109604 57836 109605 57900
rect 109539 57835 109605 57836
rect 105859 57220 105925 57221
rect 105859 57156 105860 57220
rect 105924 57156 105925 57220
rect 105859 57155 105925 57156
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 39454 110414 58000
rect 111198 57901 111258 59470
rect 112118 59470 112292 59530
rect 113222 59470 113380 59530
rect 113590 59470 113652 59530
rect 115768 59530 115828 60106
rect 116040 59530 116100 60106
rect 116992 59530 117052 60106
rect 118080 59530 118140 60106
rect 118488 59530 118548 60106
rect 119168 59530 119228 60106
rect 120936 59530 120996 60106
rect 115768 59470 115858 59530
rect 111195 57900 111261 57901
rect 111195 57836 111196 57900
rect 111260 57836 111261 57900
rect 111195 57835 111261 57836
rect 112118 57493 112178 59470
rect 113222 57493 113282 59470
rect 113590 58173 113650 59470
rect 113587 58172 113653 58173
rect 113587 58108 113588 58172
rect 113652 58108 113653 58172
rect 113587 58107 113653 58108
rect 112115 57492 112181 57493
rect 112115 57428 112116 57492
rect 112180 57428 112181 57492
rect 112115 57427 112181 57428
rect 113219 57492 113285 57493
rect 113219 57428 113220 57492
rect 113284 57428 113285 57492
rect 113219 57427 113285 57428
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 43174 114134 58000
rect 115798 57629 115858 59470
rect 115982 59470 116100 59530
rect 116902 59470 117052 59530
rect 118006 59470 118140 59530
rect 118374 59470 118548 59530
rect 119110 59470 119228 59530
rect 120766 59470 120996 59530
rect 123520 59530 123580 60106
rect 125968 59530 126028 60106
rect 123520 59470 123586 59530
rect 115982 58581 116042 59470
rect 115979 58580 116045 58581
rect 115979 58516 115980 58580
rect 116044 58516 116045 58580
rect 115979 58515 116045 58516
rect 116902 57901 116962 59470
rect 116899 57900 116965 57901
rect 116899 57836 116900 57900
rect 116964 57836 116965 57900
rect 116899 57835 116965 57836
rect 115795 57628 115861 57629
rect 115795 57564 115796 57628
rect 115860 57564 115861 57628
rect 115795 57563 115861 57564
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 46894 117854 58000
rect 118006 57901 118066 59470
rect 118003 57900 118069 57901
rect 118003 57836 118004 57900
rect 118068 57836 118069 57900
rect 118003 57835 118069 57836
rect 118374 57493 118434 59470
rect 119110 57629 119170 59470
rect 120766 57901 120826 59470
rect 120763 57900 120829 57901
rect 120763 57836 120764 57900
rect 120828 57836 120829 57900
rect 120763 57835 120829 57836
rect 119107 57628 119173 57629
rect 119107 57564 119108 57628
rect 119172 57564 119173 57628
rect 119107 57563 119173 57564
rect 118371 57492 118437 57493
rect 118371 57428 118372 57492
rect 118436 57428 118437 57492
rect 118371 57427 118437 57428
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 50614 121574 58000
rect 123526 57901 123586 59470
rect 125918 59470 126028 59530
rect 128280 59530 128340 60106
rect 131000 59530 131060 60106
rect 128280 59470 128370 59530
rect 125918 58989 125978 59470
rect 125915 58988 125981 58989
rect 125915 58924 125916 58988
rect 125980 58924 125981 58988
rect 125915 58923 125981 58924
rect 128310 58173 128370 59470
rect 130886 59470 131060 59530
rect 133448 59530 133508 60106
rect 135896 59530 135956 60106
rect 138480 59530 138540 60106
rect 140928 59530 140988 60106
rect 143512 59669 143572 60106
rect 143509 59668 143575 59669
rect 143509 59604 143510 59668
rect 143574 59604 143575 59668
rect 143509 59603 143575 59604
rect 145960 59530 146020 60106
rect 133448 59470 133522 59530
rect 128307 58172 128373 58173
rect 128307 58108 128308 58172
rect 128372 58108 128373 58172
rect 128307 58107 128373 58108
rect 123523 57900 123589 57901
rect 123523 57836 123524 57900
rect 123588 57836 123589 57900
rect 123523 57835 123589 57836
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 58000
rect 130886 57901 130946 59470
rect 130883 57900 130949 57901
rect 130883 57836 130884 57900
rect 130948 57836 130949 57900
rect 130883 57835 130949 57836
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 25174 132134 58000
rect 133462 56677 133522 59470
rect 135854 59470 135956 59530
rect 138430 59470 138540 59530
rect 140822 59470 140988 59530
rect 145606 59470 146020 59530
rect 148544 59530 148604 60106
rect 150992 59530 151052 60106
rect 153440 59530 153500 60106
rect 148544 59470 148610 59530
rect 135854 59125 135914 59470
rect 138430 59125 138490 59470
rect 140822 59261 140882 59470
rect 140819 59260 140885 59261
rect 140819 59196 140820 59260
rect 140884 59196 140885 59260
rect 140819 59195 140885 59196
rect 135851 59124 135917 59125
rect 135851 59060 135852 59124
rect 135916 59060 135917 59124
rect 135851 59059 135917 59060
rect 138427 59124 138493 59125
rect 138427 59060 138428 59124
rect 138492 59060 138493 59124
rect 138427 59059 138493 59060
rect 133459 56676 133525 56677
rect 133459 56612 133460 56676
rect 133524 56612 133525 56676
rect 133459 56611 133525 56612
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 28894 135854 58000
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 32614 139574 58000
rect 145606 57901 145666 59470
rect 148550 59261 148610 59470
rect 150942 59470 151052 59530
rect 153334 59470 153500 59530
rect 155888 59530 155948 60106
rect 158472 59530 158532 60106
rect 160920 59530 160980 60106
rect 163368 59530 163428 60106
rect 165952 59530 166012 60106
rect 183224 59530 183284 60106
rect 155888 59470 155970 59530
rect 158472 59470 158546 59530
rect 150942 59261 151002 59470
rect 148547 59260 148613 59261
rect 148547 59196 148548 59260
rect 148612 59196 148613 59260
rect 148547 59195 148613 59196
rect 150939 59260 151005 59261
rect 150939 59196 150940 59260
rect 151004 59196 151005 59260
rect 150939 59195 151005 59196
rect 153334 58173 153394 59470
rect 153331 58172 153397 58173
rect 153331 58108 153332 58172
rect 153396 58108 153397 58172
rect 153331 58107 153397 58108
rect 145603 57900 145669 57901
rect 145603 57836 145604 57900
rect 145668 57836 145669 57900
rect 145603 57835 145669 57836
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 39454 146414 58000
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 43174 150134 58000
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 46894 153854 58000
rect 155910 57629 155970 59470
rect 155907 57628 155973 57629
rect 155907 57564 155908 57628
rect 155972 57564 155973 57628
rect 155907 57563 155973 57564
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 50614 157574 58000
rect 158486 56405 158546 59470
rect 160878 59470 160980 59530
rect 163270 59470 163428 59530
rect 165846 59470 166012 59530
rect 183142 59470 183284 59530
rect 183360 59530 183420 60106
rect 183360 59470 183570 59530
rect 160878 57629 160938 59470
rect 160875 57628 160941 57629
rect 160875 57564 160876 57628
rect 160940 57564 160941 57628
rect 160875 57563 160941 57564
rect 163270 56677 163330 59470
rect 163794 57454 164414 58000
rect 165846 57629 165906 59470
rect 165843 57628 165909 57629
rect 165843 57564 165844 57628
rect 165908 57564 165909 57628
rect 165843 57563 165909 57564
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163267 56676 163333 56677
rect 163267 56612 163268 56676
rect 163332 56612 163333 56676
rect 163267 56611 163333 56612
rect 158483 56404 158549 56405
rect 158483 56340 158484 56404
rect 158548 56340 158549 56404
rect 158483 56339 158549 56340
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 25174 168134 58000
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 28894 171854 58000
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 32614 175574 58000
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 39454 182414 58000
rect 183142 57765 183202 59470
rect 183510 57901 183570 59470
rect 183507 57900 183573 57901
rect 183507 57836 183508 57900
rect 183572 57836 183573 57900
rect 183507 57835 183573 57836
rect 183139 57764 183205 57765
rect 183139 57700 183140 57764
rect 183204 57700 183205 57764
rect 183139 57699 183205 57700
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 43174 186134 58000
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 46894 189854 58000
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 50614 193574 58000
rect 197862 56133 197922 490723
rect 198043 490380 198109 490381
rect 198043 490316 198044 490380
rect 198108 490316 198109 490380
rect 198043 490315 198109 490316
rect 198046 273189 198106 490315
rect 198043 273188 198109 273189
rect 198043 273124 198044 273188
rect 198108 273124 198109 273188
rect 198043 273123 198109 273124
rect 198230 273053 198290 491131
rect 199331 491060 199397 491061
rect 199331 490996 199332 491060
rect 199396 490996 199397 491060
rect 202643 491060 202709 491061
rect 199331 490995 199397 490996
rect 198411 490244 198477 490245
rect 198411 490180 198412 490244
rect 198476 490180 198477 490244
rect 198411 490179 198477 490180
rect 198414 381037 198474 490179
rect 198963 466172 199029 466173
rect 198963 466108 198964 466172
rect 199028 466108 199029 466172
rect 198963 466107 199029 466108
rect 198779 465764 198845 465765
rect 198779 465700 198780 465764
rect 198844 465700 198845 465764
rect 198779 465699 198845 465700
rect 198411 381036 198477 381037
rect 198411 380972 198412 381036
rect 198476 380972 198477 381036
rect 198411 380971 198477 380972
rect 198227 273052 198293 273053
rect 198227 272988 198228 273052
rect 198292 272988 198293 273052
rect 198227 272987 198293 272988
rect 198782 271557 198842 465699
rect 198966 271693 199026 466107
rect 199334 272917 199394 490995
rect 199794 489454 200414 491000
rect 202643 490996 202644 491060
rect 202708 490996 202709 491060
rect 206691 491060 206757 491061
rect 202643 490995 202709 490996
rect 201355 490924 201421 490925
rect 201355 490860 201356 490924
rect 201420 490860 201421 490924
rect 201355 490859 201421 490860
rect 200619 490652 200685 490653
rect 200619 490588 200620 490652
rect 200684 490588 200685 490652
rect 200619 490587 200685 490588
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199515 469028 199581 469029
rect 199515 468964 199516 469028
rect 199580 468964 199581 469028
rect 199515 468963 199581 468964
rect 199331 272916 199397 272917
rect 199331 272852 199332 272916
rect 199396 272852 199397 272916
rect 199331 272851 199397 272852
rect 199518 272781 199578 468963
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 364394 200414 380898
rect 199794 364158 199826 364394
rect 200062 364158 200146 364394
rect 200382 364158 200414 364394
rect 199794 364074 200414 364158
rect 199794 363838 199826 364074
rect 200062 363838 200146 364074
rect 200382 363838 200414 364074
rect 199794 345454 200414 363838
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199515 272780 199581 272781
rect 199515 272716 199516 272780
rect 199580 272716 199581 272780
rect 199515 272715 199581 272716
rect 198963 271692 199029 271693
rect 198963 271628 198964 271692
rect 199028 271628 199029 271692
rect 198963 271627 199029 271628
rect 198779 271556 198845 271557
rect 198779 271492 198780 271556
rect 198844 271492 198845 271556
rect 198779 271491 198845 271492
rect 199794 256394 200414 272898
rect 199794 256158 199826 256394
rect 200062 256158 200146 256394
rect 200382 256158 200414 256394
rect 199794 256074 200414 256158
rect 199794 255838 199826 256074
rect 200062 255838 200146 256074
rect 200382 255838 200414 256074
rect 199794 237454 200414 255838
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 148394 200414 164898
rect 199794 148158 199826 148394
rect 200062 148158 200146 148394
rect 200382 148158 200414 148394
rect 199794 148074 200414 148158
rect 199794 147838 199826 148074
rect 200062 147838 200146 148074
rect 200382 147838 200414 148074
rect 199794 129454 200414 147838
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 200622 59397 200682 490587
rect 200987 490380 201053 490381
rect 200987 490316 200988 490380
rect 201052 490316 201053 490380
rect 200987 490315 201053 490316
rect 200803 468892 200869 468893
rect 200803 468828 200804 468892
rect 200868 468828 200869 468892
rect 200803 468827 200869 468828
rect 200806 165205 200866 468827
rect 200990 381037 201050 490315
rect 200987 381036 201053 381037
rect 200987 380972 200988 381036
rect 201052 380972 201053 381036
rect 200987 380971 201053 380972
rect 200803 165204 200869 165205
rect 200803 165140 200804 165204
rect 200868 165140 200869 165204
rect 200803 165139 200869 165140
rect 200619 59396 200685 59397
rect 200619 59332 200620 59396
rect 200684 59332 200685 59396
rect 200619 59331 200685 59332
rect 201358 58989 201418 490859
rect 202091 490516 202157 490517
rect 202091 490452 202092 490516
rect 202156 490452 202157 490516
rect 202091 490451 202157 490452
rect 201355 58988 201421 58989
rect 201355 58924 201356 58988
rect 201420 58924 201421 58988
rect 201355 58923 201421 58924
rect 202094 58717 202154 490451
rect 202275 482220 202341 482221
rect 202275 482156 202276 482220
rect 202340 482156 202341 482220
rect 202275 482155 202341 482156
rect 202091 58716 202157 58717
rect 202091 58652 202092 58716
rect 202156 58652 202157 58716
rect 202091 58651 202157 58652
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 202278 57357 202338 482155
rect 202459 472564 202525 472565
rect 202459 472500 202460 472564
rect 202524 472500 202525 472564
rect 202459 472499 202525 472500
rect 202462 164797 202522 472499
rect 202459 164796 202525 164797
rect 202459 164732 202460 164796
rect 202524 164732 202525 164796
rect 202459 164731 202525 164732
rect 202646 58853 202706 490995
rect 203514 476114 204134 491000
rect 206691 490996 206692 491060
rect 206756 490996 206757 491060
rect 206691 490995 206757 490996
rect 205219 490924 205285 490925
rect 205219 490860 205220 490924
rect 205284 490860 205285 490924
rect 205219 490859 205285 490860
rect 204851 480860 204917 480861
rect 204851 480796 204852 480860
rect 204916 480796 204917 480860
rect 204851 480795 204917 480796
rect 203514 475878 203546 476114
rect 203782 475878 203866 476114
rect 204102 475878 204134 476114
rect 203514 475794 204134 475878
rect 203514 475558 203546 475794
rect 203782 475558 203866 475794
rect 204102 475558 204134 475794
rect 203195 474332 203261 474333
rect 203195 474268 203196 474332
rect 203260 474268 203261 474332
rect 203195 474267 203261 474268
rect 203011 471884 203077 471885
rect 203011 471820 203012 471884
rect 203076 471820 203077 471884
rect 203011 471819 203077 471820
rect 203014 164117 203074 471819
rect 203011 164116 203077 164117
rect 203011 164052 203012 164116
rect 203076 164052 203077 164116
rect 203011 164051 203077 164052
rect 202643 58852 202709 58853
rect 202643 58788 202644 58852
rect 202708 58788 202709 58852
rect 202643 58787 202709 58788
rect 202275 57356 202341 57357
rect 202275 57292 202276 57356
rect 202340 57292 202341 57356
rect 202275 57291 202341 57292
rect 203198 57221 203258 474267
rect 203514 457174 204134 475558
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 368114 204134 384618
rect 203514 367878 203546 368114
rect 203782 367878 203866 368114
rect 204102 367878 204134 368114
rect 203514 367794 204134 367878
rect 203514 367558 203546 367794
rect 203782 367558 203866 367794
rect 204102 367558 204134 367794
rect 203514 349174 204134 367558
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 277174 204134 312618
rect 203514 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 204134 277174
rect 203514 276854 204134 276938
rect 203514 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 204134 276854
rect 203514 260114 204134 276618
rect 203514 259878 203546 260114
rect 203782 259878 203866 260114
rect 204102 259878 204134 260114
rect 203514 259794 204134 259878
rect 203514 259558 203546 259794
rect 203782 259558 203866 259794
rect 204102 259558 204134 259794
rect 203514 241174 204134 259558
rect 203514 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 204134 241174
rect 203514 240854 204134 240938
rect 203514 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 204134 240854
rect 203514 205174 204134 240618
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 152114 204134 168618
rect 203514 151878 203546 152114
rect 203782 151878 203866 152114
rect 204102 151878 204134 152114
rect 203514 151794 204134 151878
rect 203514 151558 203546 151794
rect 203782 151558 203866 151794
rect 204102 151558 204134 151794
rect 203514 133174 204134 151558
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 199794 57134 200414 57218
rect 203195 57220 203261 57221
rect 203195 57156 203196 57220
rect 203260 57156 203261 57220
rect 203195 57155 203261 57156
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 197859 56132 197925 56133
rect 197859 56068 197860 56132
rect 197924 56068 197925 56132
rect 197859 56067 197925 56068
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 204854 3909 204914 480795
rect 205035 471748 205101 471749
rect 205035 471684 205036 471748
rect 205100 471684 205101 471748
rect 205035 471683 205101 471684
rect 205038 163981 205098 471683
rect 205035 163980 205101 163981
rect 205035 163916 205036 163980
rect 205100 163916 205101 163980
rect 205035 163915 205101 163916
rect 205222 59261 205282 490859
rect 205403 490516 205469 490517
rect 205403 490452 205404 490516
rect 205468 490452 205469 490516
rect 205403 490451 205469 490452
rect 205219 59260 205285 59261
rect 205219 59196 205220 59260
rect 205284 59196 205285 59260
rect 205219 59195 205285 59196
rect 205406 56541 205466 490451
rect 206139 476780 206205 476781
rect 206139 476716 206140 476780
rect 206204 476716 206205 476780
rect 206139 476715 206205 476716
rect 206142 57765 206202 476715
rect 206323 467124 206389 467125
rect 206323 467060 206324 467124
rect 206388 467060 206389 467124
rect 206323 467059 206389 467060
rect 206326 166973 206386 467059
rect 206323 166972 206389 166973
rect 206323 166908 206324 166972
rect 206388 166908 206389 166972
rect 206323 166907 206389 166908
rect 206694 59125 206754 490995
rect 206875 490380 206941 490381
rect 206875 490316 206876 490380
rect 206940 490316 206941 490380
rect 206875 490315 206941 490316
rect 206691 59124 206757 59125
rect 206691 59060 206692 59124
rect 206756 59060 206757 59124
rect 206691 59059 206757 59060
rect 206139 57764 206205 57765
rect 206139 57700 206140 57764
rect 206204 57700 206205 57764
rect 206139 57699 206205 57700
rect 205403 56540 205469 56541
rect 205403 56476 205404 56540
rect 205468 56476 205469 56540
rect 205403 56475 205469 56476
rect 206878 56269 206938 490315
rect 207234 479834 207854 491000
rect 207979 483852 208045 483853
rect 207979 483788 207980 483852
rect 208044 483788 208045 483852
rect 207979 483787 208045 483788
rect 207234 479598 207266 479834
rect 207502 479598 207586 479834
rect 207822 479598 207854 479834
rect 207234 479514 207854 479598
rect 207234 479278 207266 479514
rect 207502 479278 207586 479514
rect 207822 479278 207854 479514
rect 207234 460894 207854 479278
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 369954 207854 388338
rect 207234 369718 207266 369954
rect 207502 369718 207586 369954
rect 207822 369718 207854 369954
rect 207234 369634 207854 369718
rect 207234 369398 207266 369634
rect 207502 369398 207586 369634
rect 207822 369398 207854 369634
rect 207234 352894 207854 369398
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 280894 207854 316338
rect 207234 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 207854 280894
rect 207234 280574 207854 280658
rect 207234 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 207854 280574
rect 207234 261954 207854 280338
rect 207234 261718 207266 261954
rect 207502 261718 207586 261954
rect 207822 261718 207854 261954
rect 207234 261634 207854 261718
rect 207234 261398 207266 261634
rect 207502 261398 207586 261634
rect 207822 261398 207854 261634
rect 207234 244894 207854 261398
rect 207234 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 207854 244894
rect 207234 244574 207854 244658
rect 207234 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 207854 244574
rect 207234 208894 207854 244338
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 155834 207854 172338
rect 207234 155598 207266 155834
rect 207502 155598 207586 155834
rect 207822 155598 207854 155834
rect 207234 155514 207854 155598
rect 207234 155278 207266 155514
rect 207502 155278 207586 155514
rect 207822 155278 207854 155514
rect 207234 136894 207854 155278
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 207234 64894 207854 100338
rect 207982 70005 208042 483787
rect 208347 478140 208413 478141
rect 208347 478076 208348 478140
rect 208412 478076 208413 478140
rect 208347 478075 208413 478076
rect 208163 466036 208229 466037
rect 208163 465972 208164 466036
rect 208228 465972 208229 466036
rect 208163 465971 208229 465972
rect 208166 166701 208226 465971
rect 208350 378589 208410 478075
rect 208347 378588 208413 378589
rect 208347 378524 208348 378588
rect 208412 378524 208413 378588
rect 208347 378523 208413 378524
rect 208163 166700 208229 166701
rect 208163 166636 208164 166700
rect 208228 166636 208229 166700
rect 208163 166635 208229 166636
rect 207979 70004 208045 70005
rect 207979 69940 207980 70004
rect 208044 69940 208045 70004
rect 207979 69939 208045 69940
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 206875 56268 206941 56269
rect 206875 56204 206876 56268
rect 206940 56204 206941 56268
rect 206875 56203 206941 56204
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 204851 3908 204917 3909
rect 204851 3844 204852 3908
rect 204916 3844 204917 3908
rect 204851 3843 204917 3844
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 -5146 207854 28338
rect 208902 4045 208962 491811
rect 216627 491196 216693 491197
rect 216627 491132 216628 491196
rect 216692 491132 216693 491196
rect 216627 491131 216693 491132
rect 219939 491196 220005 491197
rect 219939 491132 219940 491196
rect 220004 491132 220005 491196
rect 219939 491131 220005 491132
rect 209635 490380 209701 490381
rect 209635 490316 209636 490380
rect 209700 490316 209701 490380
rect 209635 490315 209701 490316
rect 209638 56405 209698 490315
rect 209819 485076 209885 485077
rect 209819 485012 209820 485076
rect 209884 485012 209885 485076
rect 209819 485011 209885 485012
rect 209822 379541 209882 485011
rect 210371 482220 210437 482221
rect 210371 482156 210372 482220
rect 210436 482156 210437 482220
rect 210371 482155 210437 482156
rect 209819 379540 209885 379541
rect 209819 379476 209820 379540
rect 209884 379476 209885 379540
rect 209819 379475 209885 379476
rect 209635 56404 209701 56405
rect 209635 56340 209636 56404
rect 209700 56340 209701 56404
rect 209635 56339 209701 56340
rect 208899 4044 208965 4045
rect 208899 3980 208900 4044
rect 208964 3980 208965 4044
rect 208899 3979 208965 3980
rect 210374 3773 210434 482155
rect 210954 481674 211574 491000
rect 213315 490652 213381 490653
rect 213315 490588 213316 490652
rect 213380 490588 213381 490652
rect 213315 490587 213381 490588
rect 213131 489156 213197 489157
rect 213131 489092 213132 489156
rect 213196 489092 213197 489156
rect 213131 489091 213197 489092
rect 211659 483716 211725 483717
rect 211659 483652 211660 483716
rect 211724 483652 211725 483716
rect 211659 483651 211725 483652
rect 210954 481438 210986 481674
rect 211222 481438 211306 481674
rect 211542 481438 211574 481674
rect 210954 481354 211574 481438
rect 210954 481118 210986 481354
rect 211222 481118 211306 481354
rect 211542 481118 211574 481354
rect 210555 468756 210621 468757
rect 210555 468692 210556 468756
rect 210620 468692 210621 468756
rect 210555 468691 210621 468692
rect 210558 166837 210618 468691
rect 210954 464614 211574 481118
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 373674 211574 392058
rect 210954 373438 210986 373674
rect 211222 373438 211306 373674
rect 211542 373438 211574 373674
rect 210954 373354 211574 373438
rect 210954 373118 210986 373354
rect 211222 373118 211306 373354
rect 211542 373118 211574 373354
rect 210954 356614 211574 373118
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 284614 211574 320058
rect 210954 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 211574 284614
rect 210954 284294 211574 284378
rect 210954 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 211574 284294
rect 210954 265674 211574 284058
rect 210954 265438 210986 265674
rect 211222 265438 211306 265674
rect 211542 265438 211574 265674
rect 210954 265354 211574 265438
rect 210954 265118 210986 265354
rect 211222 265118 211306 265354
rect 211542 265118 211574 265354
rect 210954 248614 211574 265118
rect 210954 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 211574 248614
rect 210954 248294 211574 248378
rect 210954 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 211574 248294
rect 210954 212614 211574 248058
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210555 166836 210621 166837
rect 210555 166772 210556 166836
rect 210620 166772 210621 166836
rect 210555 166771 210621 166772
rect 210954 157674 211574 176058
rect 210954 157438 210986 157674
rect 211222 157438 211306 157674
rect 211542 157438 211574 157674
rect 210954 157354 211574 157438
rect 210954 157118 210986 157354
rect 211222 157118 211306 157354
rect 211542 157118 211574 157354
rect 210954 140614 211574 157118
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 211662 56677 211722 483651
rect 211843 482492 211909 482493
rect 211843 482428 211844 482492
rect 211908 482428 211909 482492
rect 211843 482427 211909 482428
rect 211846 378045 211906 482427
rect 211843 378044 211909 378045
rect 211843 377980 211844 378044
rect 211908 377980 211909 378044
rect 211843 377979 211909 377980
rect 213134 57493 213194 489091
rect 213318 378045 213378 490587
rect 214051 482356 214117 482357
rect 214051 482292 214052 482356
rect 214116 482292 214117 482356
rect 214051 482291 214117 482292
rect 213867 476916 213933 476917
rect 213867 476852 213868 476916
rect 213932 476852 213933 476916
rect 213867 476851 213933 476852
rect 213315 378044 213381 378045
rect 213315 377980 213316 378044
rect 213380 377980 213381 378044
rect 213315 377979 213381 377980
rect 213870 271829 213930 476851
rect 214054 376549 214114 482291
rect 215891 480996 215957 480997
rect 215891 480932 215892 480996
rect 215956 480932 215957 480996
rect 215891 480931 215957 480932
rect 215339 475420 215405 475421
rect 215339 475356 215340 475420
rect 215404 475356 215405 475420
rect 215339 475355 215405 475356
rect 214235 474196 214301 474197
rect 214235 474132 214236 474196
rect 214300 474132 214301 474196
rect 214235 474131 214301 474132
rect 214238 376685 214298 474131
rect 215342 378045 215402 475355
rect 215339 378044 215405 378045
rect 215339 377980 215340 378044
rect 215404 377980 215405 378044
rect 215339 377979 215405 377980
rect 214235 376684 214301 376685
rect 214235 376620 214236 376684
rect 214300 376620 214301 376684
rect 214235 376619 214301 376620
rect 214051 376548 214117 376549
rect 214051 376484 214052 376548
rect 214116 376484 214117 376548
rect 214051 376483 214117 376484
rect 213867 271828 213933 271829
rect 213867 271764 213868 271828
rect 213932 271764 213933 271828
rect 213867 271763 213933 271764
rect 215894 57629 215954 480931
rect 216075 479500 216141 479501
rect 216075 479436 216076 479500
rect 216140 479436 216141 479500
rect 216075 479435 216141 479436
rect 215891 57628 215957 57629
rect 215891 57564 215892 57628
rect 215956 57564 215957 57628
rect 215891 57563 215957 57564
rect 213131 57492 213197 57493
rect 213131 57428 213132 57492
rect 213196 57428 213197 57492
rect 213131 57427 213197 57428
rect 216078 57085 216138 479435
rect 216259 474468 216325 474469
rect 216259 474404 216260 474468
rect 216324 474404 216325 474468
rect 216259 474403 216325 474404
rect 216262 165341 216322 474403
rect 216630 380221 216690 491131
rect 216811 491060 216877 491061
rect 216811 490996 216812 491060
rect 216876 490996 216877 491060
rect 216811 490995 216877 490996
rect 216814 396677 216874 490995
rect 217547 490516 217613 490517
rect 217547 490452 217548 490516
rect 217612 490452 217613 490516
rect 217547 490451 217613 490452
rect 217179 471612 217245 471613
rect 217179 471548 217180 471612
rect 217244 471548 217245 471612
rect 217179 471547 217245 471548
rect 216811 396676 216877 396677
rect 216811 396612 216812 396676
rect 216876 396612 216877 396676
rect 216811 396611 216877 396612
rect 216627 380220 216693 380221
rect 216627 380156 216628 380220
rect 216692 380156 216693 380220
rect 216627 380155 216693 380156
rect 216627 374644 216693 374645
rect 216627 374580 216628 374644
rect 216692 374580 216693 374644
rect 216627 374579 216693 374580
rect 216630 252517 216690 374579
rect 217182 272509 217242 471547
rect 217550 380765 217610 490451
rect 217794 471454 218414 491000
rect 219019 490788 219085 490789
rect 219019 490724 219020 490788
rect 219084 490724 219085 490788
rect 219019 490723 219085 490724
rect 218835 490652 218901 490653
rect 218835 490588 218836 490652
rect 218900 490588 218901 490652
rect 218835 490587 218901 490588
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 466308 218414 470898
rect 217547 380764 217613 380765
rect 217547 380700 217548 380764
rect 217612 380700 217613 380764
rect 217547 380699 217613 380700
rect 217363 379676 217429 379677
rect 217363 379612 217364 379676
rect 217428 379612 217429 379676
rect 217363 379611 217429 379612
rect 217179 272508 217245 272509
rect 217179 272444 217180 272508
rect 217244 272444 217245 272508
rect 217179 272443 217245 272444
rect 217366 270061 217426 379611
rect 218838 379541 218898 490587
rect 218835 379540 218901 379541
rect 218835 379476 218836 379540
rect 218900 379476 218901 379540
rect 218835 379475 218901 379476
rect 217547 375732 217613 375733
rect 217547 375668 217548 375732
rect 217612 375668 217613 375732
rect 217547 375667 217613 375668
rect 217363 270060 217429 270061
rect 217363 269996 217364 270060
rect 217428 269996 217429 270060
rect 217363 269995 217429 269996
rect 217550 268429 217610 375667
rect 217794 363454 218414 379000
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 359308 218414 362898
rect 217547 268428 217613 268429
rect 217547 268364 217548 268428
rect 217612 268364 217613 268428
rect 217547 268363 217613 268364
rect 217794 255454 218414 272000
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 216627 252516 216693 252517
rect 216627 252452 216628 252516
rect 216692 252452 216693 252516
rect 216627 252451 216693 252452
rect 217363 252516 217429 252517
rect 217363 252452 217364 252516
rect 217428 252452 217429 252516
rect 217363 252451 217429 252452
rect 216259 165340 216325 165341
rect 216259 165276 216260 165340
rect 216324 165276 216325 165340
rect 216259 165275 216325 165276
rect 217366 163573 217426 252451
rect 217794 252308 218414 254898
rect 217547 251836 217613 251837
rect 217547 251772 217548 251836
rect 217612 251772 217613 251836
rect 217547 251771 217613 251772
rect 217363 163572 217429 163573
rect 217363 163508 217364 163572
rect 217428 163508 217429 163572
rect 217363 163507 217429 163508
rect 217550 162757 217610 251771
rect 217547 162756 217613 162757
rect 217547 162692 217548 162756
rect 217612 162692 217613 162756
rect 217547 162691 217613 162692
rect 217547 162620 217613 162621
rect 217547 162556 217548 162620
rect 217612 162556 217613 162620
rect 217547 162555 217613 162556
rect 217363 148340 217429 148341
rect 217363 148276 217364 148340
rect 217428 148276 217429 148340
rect 217363 148275 217429 148276
rect 217179 144940 217245 144941
rect 217179 144876 217180 144940
rect 217244 144876 217245 144940
rect 217179 144875 217245 144876
rect 217182 58309 217242 144875
rect 217179 58308 217245 58309
rect 217179 58244 217180 58308
rect 217244 58244 217245 58308
rect 217179 58243 217245 58244
rect 216075 57084 216141 57085
rect 216075 57020 216076 57084
rect 216140 57020 216141 57084
rect 216075 57019 216141 57020
rect 211659 56676 211725 56677
rect 211659 56612 211660 56676
rect 211724 56612 211725 56676
rect 211659 56611 211725 56612
rect 217366 55045 217426 148275
rect 217550 58445 217610 162555
rect 217794 147454 218414 165000
rect 217794 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 218414 147454
rect 217794 147134 218414 147218
rect 217794 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 218414 147134
rect 217794 145308 218414 146898
rect 219022 59533 219082 490723
rect 219203 490516 219269 490517
rect 219203 490452 219204 490516
rect 219268 490452 219269 490516
rect 219203 490451 219269 490452
rect 219019 59532 219085 59533
rect 219019 59468 219020 59532
rect 219084 59468 219085 59532
rect 219019 59467 219085 59468
rect 219206 58581 219266 490451
rect 219942 167109 220002 491131
rect 221514 475174 222134 491000
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 466308 222134 474618
rect 225234 478894 225854 491000
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 466308 225854 478338
rect 228954 482614 229574 491000
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 466308 229574 482058
rect 235794 489454 236414 491000
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 466308 236414 488898
rect 239514 476114 240134 491000
rect 239514 475878 239546 476114
rect 239782 475878 239866 476114
rect 240102 475878 240134 476114
rect 239514 475794 240134 475878
rect 239514 475558 239546 475794
rect 239782 475558 239866 475794
rect 240102 475558 240134 475794
rect 239514 466308 240134 475558
rect 243234 479834 243854 491000
rect 243234 479598 243266 479834
rect 243502 479598 243586 479834
rect 243822 479598 243854 479834
rect 243234 479514 243854 479598
rect 243234 479278 243266 479514
rect 243502 479278 243586 479514
rect 243822 479278 243854 479514
rect 243234 466308 243854 479278
rect 246954 481674 247574 491000
rect 246954 481438 246986 481674
rect 247222 481438 247306 481674
rect 247542 481438 247574 481674
rect 246954 481354 247574 481438
rect 246954 481118 246986 481354
rect 247222 481118 247306 481354
rect 247542 481118 247574 481354
rect 246954 466308 247574 481118
rect 253794 471454 254414 491000
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 466308 254414 470898
rect 257514 475174 258134 491000
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 466308 258134 474618
rect 261234 478894 261854 491000
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 466308 261854 478338
rect 264954 482614 265574 491000
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 466308 265574 482058
rect 271794 489454 272414 491000
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 466308 272414 488898
rect 275514 476114 276134 491000
rect 275514 475878 275546 476114
rect 275782 475878 275866 476114
rect 276102 475878 276134 476114
rect 275514 475794 276134 475878
rect 275514 475558 275546 475794
rect 275782 475558 275866 475794
rect 276102 475558 276134 475794
rect 275514 466308 276134 475558
rect 279234 479834 279854 491000
rect 279234 479598 279266 479834
rect 279502 479598 279586 479834
rect 279822 479598 279854 479834
rect 279234 479514 279854 479598
rect 279234 479278 279266 479514
rect 279502 479278 279586 479514
rect 279822 479278 279854 479514
rect 279234 466308 279854 479278
rect 282954 481674 283574 491000
rect 282954 481438 282986 481674
rect 283222 481438 283306 481674
rect 283542 481438 283574 481674
rect 282954 481354 283574 481438
rect 282954 481118 282986 481354
rect 283222 481118 283306 481354
rect 283542 481118 283574 481354
rect 282954 466308 283574 481118
rect 289794 471454 290414 491000
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 466308 290414 470898
rect 293514 475174 294134 491000
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 466308 294134 474618
rect 297234 478894 297854 491000
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 466308 297854 478338
rect 300954 482614 301574 491000
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 466308 301574 482058
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 466308 308414 488898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 466308 312134 492618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 466308 315854 496338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 647033 326414 650898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 647033 330134 654618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 647033 333854 658338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 647033 337574 662058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 647033 344414 668898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 647033 348134 672618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 647033 351854 676338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 647033 355574 680058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 647033 362414 650898
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 647033 366134 654618
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 647033 369854 658338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 647033 373574 662058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 647033 380414 668898
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 647033 384134 672618
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 647033 387854 676338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 647033 391574 680058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 647033 398414 650898
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 647033 402134 654618
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 647033 405854 658338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 647033 409574 662058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 647033 416414 668898
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 647033 420134 672618
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 647033 423854 676338
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 647033 427574 680058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 647033 434414 650898
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 344568 633454 344888 633486
rect 344568 633218 344610 633454
rect 344846 633218 344888 633454
rect 344568 633134 344888 633218
rect 344568 632898 344610 633134
rect 344846 632898 344888 633134
rect 344568 632866 344888 632898
rect 375288 633454 375608 633486
rect 375288 633218 375330 633454
rect 375566 633218 375608 633454
rect 375288 633134 375608 633218
rect 375288 632898 375330 633134
rect 375566 632898 375608 633134
rect 375288 632866 375608 632898
rect 406008 633454 406328 633486
rect 406008 633218 406050 633454
rect 406286 633218 406328 633454
rect 406008 633134 406328 633218
rect 406008 632898 406050 633134
rect 406286 632898 406328 633134
rect 406008 632866 406328 632898
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 329208 615454 329528 615486
rect 329208 615218 329250 615454
rect 329486 615218 329528 615454
rect 329208 615134 329528 615218
rect 329208 614898 329250 615134
rect 329486 614898 329528 615134
rect 329208 614866 329528 614898
rect 359928 615454 360248 615486
rect 359928 615218 359970 615454
rect 360206 615218 360248 615454
rect 359928 615134 360248 615218
rect 359928 614898 359970 615134
rect 360206 614898 360248 615134
rect 359928 614866 360248 614898
rect 390648 615454 390968 615486
rect 390648 615218 390690 615454
rect 390926 615218 390968 615454
rect 390648 615134 390968 615218
rect 390648 614898 390690 615134
rect 390926 614898 390968 615134
rect 390648 614866 390968 614898
rect 421368 615454 421688 615486
rect 421368 615218 421410 615454
rect 421646 615218 421688 615454
rect 421368 615134 421688 615218
rect 421368 614898 421410 615134
rect 421646 614898 421688 615134
rect 421368 614866 421688 614898
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 436139 606388 436205 606389
rect 436139 606324 436140 606388
rect 436204 606324 436205 606388
rect 436139 606323 436205 606324
rect 344568 597454 344888 597486
rect 344568 597218 344610 597454
rect 344846 597218 344888 597454
rect 344568 597134 344888 597218
rect 344568 596898 344610 597134
rect 344846 596898 344888 597134
rect 344568 596866 344888 596898
rect 375288 597454 375608 597486
rect 375288 597218 375330 597454
rect 375566 597218 375608 597454
rect 375288 597134 375608 597218
rect 375288 596898 375330 597134
rect 375566 596898 375608 597134
rect 375288 596866 375608 596898
rect 406008 597454 406328 597486
rect 406008 597218 406050 597454
rect 406286 597218 406328 597454
rect 406008 597134 406328 597218
rect 406008 596898 406050 597134
rect 406286 596898 406328 597134
rect 406008 596866 406328 596898
rect 329208 579454 329528 579486
rect 329208 579218 329250 579454
rect 329486 579218 329528 579454
rect 329208 579134 329528 579218
rect 329208 578898 329250 579134
rect 329486 578898 329528 579134
rect 329208 578866 329528 578898
rect 359928 579454 360248 579486
rect 359928 579218 359970 579454
rect 360206 579218 360248 579454
rect 359928 579134 360248 579218
rect 359928 578898 359970 579134
rect 360206 578898 360248 579134
rect 359928 578866 360248 578898
rect 390648 579454 390968 579486
rect 390648 579218 390690 579454
rect 390926 579218 390968 579454
rect 390648 579134 390968 579218
rect 390648 578898 390690 579134
rect 390926 578898 390968 579134
rect 390648 578866 390968 578898
rect 421368 579454 421688 579486
rect 421368 579218 421410 579454
rect 421646 579218 421688 579454
rect 421368 579134 421688 579218
rect 421368 578898 421410 579134
rect 421646 578898 421688 579134
rect 421368 578866 421688 578898
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 344568 561454 344888 561486
rect 344568 561218 344610 561454
rect 344846 561218 344888 561454
rect 344568 561134 344888 561218
rect 344568 560898 344610 561134
rect 344846 560898 344888 561134
rect 344568 560866 344888 560898
rect 375288 561454 375608 561486
rect 375288 561218 375330 561454
rect 375566 561218 375608 561454
rect 375288 561134 375608 561218
rect 375288 560898 375330 561134
rect 375566 560898 375608 561134
rect 375288 560866 375608 560898
rect 406008 561454 406328 561486
rect 406008 561218 406050 561454
rect 406286 561218 406328 561454
rect 406008 561134 406328 561218
rect 406008 560898 406050 561134
rect 406286 560898 406328 561134
rect 406008 560866 406328 560898
rect 329208 543454 329528 543486
rect 329208 543218 329250 543454
rect 329486 543218 329528 543454
rect 329208 543134 329528 543218
rect 329208 542898 329250 543134
rect 329486 542898 329528 543134
rect 329208 542866 329528 542898
rect 359928 543454 360248 543486
rect 359928 543218 359970 543454
rect 360206 543218 360248 543454
rect 359928 543134 360248 543218
rect 359928 542898 359970 543134
rect 360206 542898 360248 543134
rect 359928 542866 360248 542898
rect 390648 543454 390968 543486
rect 390648 543218 390690 543454
rect 390926 543218 390968 543454
rect 390648 543134 390968 543218
rect 390648 542898 390690 543134
rect 390926 542898 390968 543134
rect 390648 542866 390968 542898
rect 421368 543454 421688 543486
rect 421368 543218 421410 543454
rect 421646 543218 421688 543454
rect 421368 543134 421688 543218
rect 421368 542898 421410 543134
rect 421646 542898 421688 543134
rect 421368 542866 421688 542898
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 436142 534581 436202 606323
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 436139 534580 436205 534581
rect 436139 534516 436140 534580
rect 436204 534516 436205 534580
rect 436139 534515 436205 534516
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 466308 319574 500058
rect 325794 507454 326414 532000
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 466308 326414 470898
rect 329514 511174 330134 532000
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 466308 330134 474618
rect 333234 514894 333854 532000
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 466308 333854 478338
rect 336954 518614 337574 532000
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 466308 337574 482058
rect 343794 525454 344414 532000
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 338435 466580 338501 466581
rect 338435 466516 338436 466580
rect 338500 466516 338501 466580
rect 338435 466515 338501 466516
rect 339723 466580 339789 466581
rect 339723 466516 339724 466580
rect 339788 466516 339789 466580
rect 339723 466515 339789 466516
rect 338438 464810 338498 466515
rect 339726 464810 339786 466515
rect 343794 466308 344414 488898
rect 347514 529174 348134 532000
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 466308 348134 492618
rect 351234 496894 351854 532000
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 350947 466580 351013 466581
rect 350947 466516 350948 466580
rect 351012 466516 351013 466580
rect 350947 466515 351013 466516
rect 350950 464810 351010 466515
rect 351234 466308 351854 496338
rect 354954 500614 355574 532000
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 466308 355574 500058
rect 361794 507454 362414 532000
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 357939 491196 358005 491197
rect 357939 491132 357940 491196
rect 358004 491132 358005 491196
rect 357939 491131 358005 491132
rect 338438 464750 338524 464810
rect 338464 464202 338524 464750
rect 339688 464750 339786 464810
rect 350840 464750 351010 464810
rect 339688 464202 339748 464750
rect 350840 464202 350900 464750
rect 220272 453454 220620 453486
rect 220272 453218 220328 453454
rect 220564 453218 220620 453454
rect 220272 453134 220620 453218
rect 220272 452898 220328 453134
rect 220564 452898 220620 453134
rect 220272 452866 220620 452898
rect 356000 453454 356348 453486
rect 356000 453218 356056 453454
rect 356292 453218 356348 453454
rect 356000 453134 356348 453218
rect 356000 452898 356056 453134
rect 356292 452898 356348 453134
rect 356000 452866 356348 452898
rect 220952 435454 221300 435486
rect 220952 435218 221008 435454
rect 221244 435218 221300 435454
rect 220952 435134 221300 435218
rect 220952 434898 221008 435134
rect 221244 434898 221300 435134
rect 220952 434866 221300 434898
rect 355320 435454 355668 435486
rect 355320 435218 355376 435454
rect 355612 435218 355668 435454
rect 355320 435134 355668 435218
rect 355320 434898 355376 435134
rect 355612 434898 355668 435134
rect 355320 434866 355668 434898
rect 220272 417454 220620 417486
rect 220272 417218 220328 417454
rect 220564 417218 220620 417454
rect 220272 417134 220620 417218
rect 220272 416898 220328 417134
rect 220564 416898 220620 417134
rect 220272 416866 220620 416898
rect 356000 417454 356348 417486
rect 356000 417218 356056 417454
rect 356292 417218 356348 417454
rect 356000 417134 356348 417218
rect 356000 416898 356056 417134
rect 356292 416898 356348 417134
rect 356000 416866 356348 416898
rect 220952 399454 221300 399486
rect 220952 399218 221008 399454
rect 221244 399218 221300 399454
rect 220952 399134 221300 399218
rect 220952 398898 221008 399134
rect 221244 398898 221300 399134
rect 220952 398866 221300 398898
rect 355320 399454 355668 399486
rect 355320 399218 355376 399454
rect 355612 399218 355668 399454
rect 355320 399134 355668 399218
rect 355320 398898 355376 399134
rect 355612 398898 355668 399134
rect 355320 398866 355668 398898
rect 236056 380765 236116 381106
rect 237144 380765 237204 381106
rect 236053 380764 236119 380765
rect 236053 380700 236054 380764
rect 236118 380700 236119 380764
rect 236053 380699 236119 380700
rect 237141 380764 237207 380765
rect 237141 380700 237142 380764
rect 237206 380700 237207 380764
rect 237141 380699 237207 380700
rect 238232 380490 238292 381106
rect 238158 380430 238292 380490
rect 239592 380490 239652 381106
rect 240544 380490 240604 381106
rect 241768 380490 241828 381106
rect 243128 380765 243188 381106
rect 243125 380764 243191 380765
rect 243125 380700 243126 380764
rect 243190 380700 243191 380764
rect 243125 380699 243191 380700
rect 244216 380493 244276 381106
rect 244216 380492 244293 380493
rect 239592 380430 239690 380490
rect 240544 380430 240610 380490
rect 241768 380430 241898 380490
rect 244216 380430 244228 380492
rect 238158 379269 238218 380430
rect 239630 379405 239690 380430
rect 239627 379404 239693 379405
rect 239627 379340 239628 379404
rect 239692 379340 239693 379404
rect 239627 379339 239693 379340
rect 238155 379268 238221 379269
rect 238155 379204 238156 379268
rect 238220 379204 238221 379268
rect 238155 379203 238221 379204
rect 221514 367174 222134 379000
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 359308 222134 366618
rect 225234 370894 225854 379000
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 359308 225854 370338
rect 228954 374614 229574 379000
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 359308 229574 374058
rect 235794 364394 236414 379000
rect 235794 364158 235826 364394
rect 236062 364158 236146 364394
rect 236382 364158 236414 364394
rect 235794 364074 236414 364158
rect 235794 363838 235826 364074
rect 236062 363838 236146 364074
rect 236382 363838 236414 364074
rect 235794 359308 236414 363838
rect 239514 368114 240134 379000
rect 240550 378725 240610 380430
rect 240547 378724 240613 378725
rect 240547 378660 240548 378724
rect 240612 378660 240613 378724
rect 240547 378659 240613 378660
rect 241838 378453 241898 380430
rect 244227 380428 244228 380430
rect 244292 380428 244293 380492
rect 245440 380490 245500 381106
rect 246528 380490 246588 381106
rect 247616 380490 247676 381106
rect 248296 380765 248356 381106
rect 248293 380764 248359 380765
rect 248293 380700 248294 380764
rect 248358 380700 248359 380764
rect 248293 380699 248359 380700
rect 248704 380490 248764 381106
rect 244227 380427 244293 380428
rect 245334 380430 245500 380490
rect 246438 380430 246588 380490
rect 247542 380430 247676 380490
rect 248646 380430 248764 380490
rect 250064 380490 250124 381106
rect 250744 380762 250804 381106
rect 251288 380762 251348 381106
rect 250670 380702 250804 380762
rect 251222 380702 251348 380762
rect 250064 380430 250178 380490
rect 245334 379405 245394 380430
rect 246438 379405 246498 380430
rect 247542 380357 247602 380430
rect 247539 380356 247605 380357
rect 247539 380292 247540 380356
rect 247604 380292 247605 380356
rect 247539 380291 247605 380292
rect 248646 379405 248706 380430
rect 250118 379405 250178 380430
rect 245331 379404 245397 379405
rect 245331 379340 245332 379404
rect 245396 379340 245397 379404
rect 245331 379339 245397 379340
rect 246435 379404 246501 379405
rect 246435 379340 246436 379404
rect 246500 379340 246501 379404
rect 246435 379339 246501 379340
rect 248643 379404 248709 379405
rect 248643 379340 248644 379404
rect 248708 379340 248709 379404
rect 248643 379339 248709 379340
rect 250115 379404 250181 379405
rect 250115 379340 250116 379404
rect 250180 379340 250181 379404
rect 250115 379339 250181 379340
rect 241835 378452 241901 378453
rect 241835 378388 241836 378452
rect 241900 378388 241901 378452
rect 241835 378387 241901 378388
rect 239514 367878 239546 368114
rect 239782 367878 239866 368114
rect 240102 367878 240134 368114
rect 239514 367794 240134 367878
rect 239514 367558 239546 367794
rect 239782 367558 239866 367794
rect 240102 367558 240134 367794
rect 239514 359308 240134 367558
rect 243234 369954 243854 379000
rect 243234 369718 243266 369954
rect 243502 369718 243586 369954
rect 243822 369718 243854 369954
rect 243234 369634 243854 369718
rect 243234 369398 243266 369634
rect 243502 369398 243586 369634
rect 243822 369398 243854 369634
rect 243234 359308 243854 369398
rect 246954 373674 247574 379000
rect 250670 378861 250730 380702
rect 251222 379405 251282 380702
rect 252376 380490 252436 381106
rect 253464 380490 253524 381106
rect 252326 380430 252436 380490
rect 253430 380430 253524 380490
rect 253600 380490 253660 381106
rect 254552 380765 254612 381106
rect 255912 380765 255972 381106
rect 254549 380764 254615 380765
rect 254549 380700 254550 380764
rect 254614 380700 254615 380764
rect 254549 380699 254615 380700
rect 255909 380764 255975 380765
rect 255909 380700 255910 380764
rect 255974 380700 255975 380764
rect 255909 380699 255975 380700
rect 256048 380490 256108 381106
rect 257000 380629 257060 381106
rect 258088 380629 258148 381106
rect 256997 380628 257063 380629
rect 256997 380564 256998 380628
rect 257062 380564 257063 380628
rect 256997 380563 257063 380564
rect 258085 380628 258151 380629
rect 258085 380564 258086 380628
rect 258150 380564 258151 380628
rect 258085 380563 258151 380564
rect 258496 380490 258556 381106
rect 253600 380430 253674 380490
rect 252326 379405 252386 380430
rect 253430 379405 253490 380430
rect 251219 379404 251285 379405
rect 251219 379340 251220 379404
rect 251284 379340 251285 379404
rect 251219 379339 251285 379340
rect 252323 379404 252389 379405
rect 252323 379340 252324 379404
rect 252388 379340 252389 379404
rect 252323 379339 252389 379340
rect 253427 379404 253493 379405
rect 253427 379340 253428 379404
rect 253492 379340 253493 379404
rect 253427 379339 253493 379340
rect 250667 378860 250733 378861
rect 250667 378796 250668 378860
rect 250732 378796 250733 378860
rect 250667 378795 250733 378796
rect 253614 378453 253674 380430
rect 256006 380430 256108 380490
rect 258398 380430 258556 380490
rect 259448 380490 259508 381106
rect 260672 380490 260732 381106
rect 261080 380490 261140 381106
rect 261760 380629 261820 381106
rect 261757 380628 261823 380629
rect 261757 380564 261758 380628
rect 261822 380564 261823 380628
rect 261757 380563 261823 380564
rect 262848 380490 262908 381106
rect 259448 380430 259562 380490
rect 253611 378452 253677 378453
rect 253611 378388 253612 378452
rect 253676 378388 253677 378452
rect 253611 378387 253677 378388
rect 246954 373438 246986 373674
rect 247222 373438 247306 373674
rect 247542 373438 247574 373674
rect 246954 373354 247574 373438
rect 246954 373118 246986 373354
rect 247222 373118 247306 373354
rect 247542 373118 247574 373354
rect 246954 359308 247574 373118
rect 253794 363454 254414 379000
rect 256006 378453 256066 380430
rect 256003 378452 256069 378453
rect 256003 378388 256004 378452
rect 256068 378388 256069 378452
rect 256003 378387 256069 378388
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 359308 254414 362898
rect 257514 367174 258134 379000
rect 258398 378589 258458 380430
rect 259502 380085 259562 380430
rect 260606 380430 260732 380490
rect 260974 380430 261140 380490
rect 262814 380430 262908 380490
rect 263528 380490 263588 381106
rect 263936 380490 263996 381106
rect 265296 380490 265356 381106
rect 265976 380490 266036 381106
rect 266384 380490 266444 381106
rect 267608 380490 267668 381106
rect 263528 380430 263610 380490
rect 259499 380084 259565 380085
rect 259499 380020 259500 380084
rect 259564 380020 259565 380084
rect 259499 380019 259565 380020
rect 260606 378589 260666 380430
rect 260974 378589 261034 380430
rect 258395 378588 258461 378589
rect 258395 378524 258396 378588
rect 258460 378524 258461 378588
rect 258395 378523 258461 378524
rect 260603 378588 260669 378589
rect 260603 378524 260604 378588
rect 260668 378524 260669 378588
rect 260603 378523 260669 378524
rect 260971 378588 261037 378589
rect 260971 378524 260972 378588
rect 261036 378524 261037 378588
rect 260971 378523 261037 378524
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 359308 258134 366618
rect 261234 370894 261854 379000
rect 262814 378589 262874 380430
rect 263550 378589 263610 380430
rect 263918 380430 263996 380490
rect 265206 380430 265356 380490
rect 265942 380430 266036 380490
rect 266310 380430 266444 380490
rect 267598 380430 267668 380490
rect 268288 380490 268348 381106
rect 268696 380490 268756 381106
rect 269784 380490 269844 381106
rect 271008 380629 271068 381106
rect 271005 380628 271071 380629
rect 271005 380564 271006 380628
rect 271070 380564 271071 380628
rect 271005 380563 271071 380564
rect 271144 380490 271204 381106
rect 272232 380490 272292 381106
rect 273320 380490 273380 381106
rect 273592 380490 273652 381106
rect 274408 380490 274468 381106
rect 275768 380490 275828 381106
rect 268288 380430 268394 380490
rect 268696 380430 268762 380490
rect 269784 380430 269866 380490
rect 263918 379405 263978 380430
rect 265206 379405 265266 380430
rect 263915 379404 263981 379405
rect 263915 379340 263916 379404
rect 263980 379340 263981 379404
rect 263915 379339 263981 379340
rect 265203 379404 265269 379405
rect 265203 379340 265204 379404
rect 265268 379340 265269 379404
rect 265203 379339 265269 379340
rect 262811 378588 262877 378589
rect 262811 378524 262812 378588
rect 262876 378524 262877 378588
rect 262811 378523 262877 378524
rect 263547 378588 263613 378589
rect 263547 378524 263548 378588
rect 263612 378524 263613 378588
rect 263547 378523 263613 378524
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 359308 261854 370338
rect 264954 374614 265574 379000
rect 265942 378589 266002 380430
rect 266310 378589 266370 380430
rect 267598 378589 267658 380430
rect 268334 378589 268394 380430
rect 268702 379405 268762 380430
rect 269806 379405 269866 380430
rect 271094 380430 271204 380490
rect 272198 380430 272292 380490
rect 273302 380430 273380 380490
rect 273486 380430 273652 380490
rect 274406 380430 274468 380490
rect 275694 380430 275828 380490
rect 276040 380490 276100 381106
rect 276992 380490 277052 381106
rect 276040 380430 276122 380490
rect 271094 379405 271154 380430
rect 272198 379405 272258 380430
rect 273302 379405 273362 380430
rect 268699 379404 268765 379405
rect 268699 379340 268700 379404
rect 268764 379340 268765 379404
rect 268699 379339 268765 379340
rect 269803 379404 269869 379405
rect 269803 379340 269804 379404
rect 269868 379340 269869 379404
rect 269803 379339 269869 379340
rect 271091 379404 271157 379405
rect 271091 379340 271092 379404
rect 271156 379340 271157 379404
rect 271091 379339 271157 379340
rect 272195 379404 272261 379405
rect 272195 379340 272196 379404
rect 272260 379340 272261 379404
rect 272195 379339 272261 379340
rect 273299 379404 273365 379405
rect 273299 379340 273300 379404
rect 273364 379340 273365 379404
rect 273299 379339 273365 379340
rect 265939 378588 266005 378589
rect 265939 378524 265940 378588
rect 266004 378524 266005 378588
rect 265939 378523 266005 378524
rect 266307 378588 266373 378589
rect 266307 378524 266308 378588
rect 266372 378524 266373 378588
rect 266307 378523 266373 378524
rect 267595 378588 267661 378589
rect 267595 378524 267596 378588
rect 267660 378524 267661 378588
rect 267595 378523 267661 378524
rect 268331 378588 268397 378589
rect 268331 378524 268332 378588
rect 268396 378524 268397 378588
rect 268331 378523 268397 378524
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 359308 265574 374058
rect 271794 364394 272414 379000
rect 273486 378997 273546 380430
rect 274406 379269 274466 380430
rect 275694 379405 275754 380430
rect 275691 379404 275757 379405
rect 275691 379340 275692 379404
rect 275756 379340 275757 379404
rect 275691 379339 275757 379340
rect 276062 379269 276122 380430
rect 276982 380430 277052 380490
rect 278080 380490 278140 381106
rect 278488 380490 278548 381106
rect 279168 380490 279228 381106
rect 280936 380490 280996 381106
rect 283520 380490 283580 381106
rect 278080 380430 278146 380490
rect 276982 379269 277042 380430
rect 274403 379268 274469 379269
rect 274403 379204 274404 379268
rect 274468 379204 274469 379268
rect 274403 379203 274469 379204
rect 276059 379268 276125 379269
rect 276059 379204 276060 379268
rect 276124 379204 276125 379268
rect 276059 379203 276125 379204
rect 276979 379268 277045 379269
rect 276979 379204 276980 379268
rect 277044 379204 277045 379268
rect 276979 379203 277045 379204
rect 278086 379133 278146 380430
rect 278454 380430 278548 380490
rect 279006 380430 279228 380490
rect 280846 380430 280996 380490
rect 283422 380430 283580 380490
rect 285968 380490 286028 381106
rect 288280 380490 288340 381106
rect 291000 380490 291060 381106
rect 293448 380490 293508 381106
rect 285968 380430 286058 380490
rect 278454 379269 278514 380430
rect 278451 379268 278517 379269
rect 278451 379204 278452 379268
rect 278516 379204 278517 379268
rect 278451 379203 278517 379204
rect 278083 379132 278149 379133
rect 278083 379068 278084 379132
rect 278148 379068 278149 379132
rect 278083 379067 278149 379068
rect 273483 378996 273549 378997
rect 273483 378932 273484 378996
rect 273548 378932 273549 378996
rect 273483 378931 273549 378932
rect 271794 364158 271826 364394
rect 272062 364158 272146 364394
rect 272382 364158 272414 364394
rect 271794 364074 272414 364158
rect 271794 363838 271826 364074
rect 272062 363838 272146 364074
rect 272382 363838 272414 364074
rect 271794 359308 272414 363838
rect 275514 368114 276134 379000
rect 279006 378181 279066 380430
rect 280846 379269 280906 380430
rect 283422 379269 283482 380430
rect 285998 379405 286058 380430
rect 288206 380430 288340 380490
rect 290966 380430 291060 380490
rect 293358 380430 293508 380490
rect 295896 380490 295956 381106
rect 298480 380490 298540 381106
rect 300928 380490 300988 381106
rect 303512 380490 303572 381106
rect 305960 380490 306020 381106
rect 308544 380490 308604 381106
rect 295896 380430 295994 380490
rect 298480 380430 298570 380490
rect 288206 379405 288266 380430
rect 290966 379405 291026 380430
rect 293358 379405 293418 380430
rect 295934 379405 295994 380430
rect 298510 379405 298570 380430
rect 300902 380430 300988 380490
rect 303478 380430 303572 380490
rect 305870 380430 306020 380490
rect 308446 380430 308604 380490
rect 310992 380490 311052 381106
rect 313440 380765 313500 381106
rect 313437 380764 313503 380765
rect 313437 380700 313438 380764
rect 313502 380700 313503 380764
rect 313437 380699 313503 380700
rect 315888 380629 315948 381106
rect 315885 380628 315951 380629
rect 315885 380564 315886 380628
rect 315950 380564 315951 380628
rect 318472 380626 318532 381106
rect 315885 380563 315951 380564
rect 318382 380566 318532 380626
rect 310992 380430 311082 380490
rect 285995 379404 286061 379405
rect 285995 379340 285996 379404
rect 286060 379340 286061 379404
rect 285995 379339 286061 379340
rect 288203 379404 288269 379405
rect 288203 379340 288204 379404
rect 288268 379340 288269 379404
rect 288203 379339 288269 379340
rect 290963 379404 291029 379405
rect 290963 379340 290964 379404
rect 291028 379340 291029 379404
rect 290963 379339 291029 379340
rect 293355 379404 293421 379405
rect 293355 379340 293356 379404
rect 293420 379340 293421 379404
rect 293355 379339 293421 379340
rect 295931 379404 295997 379405
rect 295931 379340 295932 379404
rect 295996 379340 295997 379404
rect 295931 379339 295997 379340
rect 298507 379404 298573 379405
rect 298507 379340 298508 379404
rect 298572 379340 298573 379404
rect 298507 379339 298573 379340
rect 300902 379269 300962 380430
rect 280843 379268 280909 379269
rect 280843 379204 280844 379268
rect 280908 379204 280909 379268
rect 280843 379203 280909 379204
rect 283419 379268 283485 379269
rect 283419 379204 283420 379268
rect 283484 379204 283485 379268
rect 283419 379203 283485 379204
rect 300899 379268 300965 379269
rect 300899 379204 300900 379268
rect 300964 379204 300965 379268
rect 300899 379203 300965 379204
rect 279003 378180 279069 378181
rect 279003 378116 279004 378180
rect 279068 378116 279069 378180
rect 279003 378115 279069 378116
rect 275514 367878 275546 368114
rect 275782 367878 275866 368114
rect 276102 367878 276134 368114
rect 275514 367794 276134 367878
rect 275514 367558 275546 367794
rect 275782 367558 275866 367794
rect 276102 367558 276134 367794
rect 275514 359308 276134 367558
rect 279234 369954 279854 379000
rect 279234 369718 279266 369954
rect 279502 369718 279586 369954
rect 279822 369718 279854 369954
rect 279234 369634 279854 369718
rect 279234 369398 279266 369634
rect 279502 369398 279586 369634
rect 279822 369398 279854 369634
rect 279234 359308 279854 369398
rect 282954 373674 283574 379000
rect 282954 373438 282986 373674
rect 283222 373438 283306 373674
rect 283542 373438 283574 373674
rect 282954 373354 283574 373438
rect 282954 373118 282986 373354
rect 283222 373118 283306 373354
rect 283542 373118 283574 373354
rect 282954 359308 283574 373118
rect 289794 363454 290414 379000
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 359308 290414 362898
rect 293514 367174 294134 379000
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 359308 294134 366618
rect 297234 370894 297854 379000
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 359308 297854 370338
rect 300954 374614 301574 379000
rect 303478 378997 303538 380430
rect 305870 379405 305930 380430
rect 308446 379405 308506 380430
rect 311022 379405 311082 380430
rect 318382 379405 318442 380566
rect 320920 380490 320980 381106
rect 323368 380901 323428 381106
rect 323365 380900 323431 380901
rect 323365 380836 323366 380900
rect 323430 380836 323431 380900
rect 323365 380835 323431 380836
rect 325952 380490 326012 381106
rect 343224 380490 343284 381106
rect 320920 380430 321018 380490
rect 320958 379405 321018 380430
rect 325926 380430 326012 380490
rect 343222 380430 343284 380490
rect 343360 380490 343420 381106
rect 343360 380430 343466 380490
rect 325926 379405 325986 380430
rect 305867 379404 305933 379405
rect 305867 379340 305868 379404
rect 305932 379340 305933 379404
rect 305867 379339 305933 379340
rect 308443 379404 308509 379405
rect 308443 379340 308444 379404
rect 308508 379340 308509 379404
rect 308443 379339 308509 379340
rect 311019 379404 311085 379405
rect 311019 379340 311020 379404
rect 311084 379340 311085 379404
rect 311019 379339 311085 379340
rect 318379 379404 318445 379405
rect 318379 379340 318380 379404
rect 318444 379340 318445 379404
rect 318379 379339 318445 379340
rect 320955 379404 321021 379405
rect 320955 379340 320956 379404
rect 321020 379340 321021 379404
rect 320955 379339 321021 379340
rect 325923 379404 325989 379405
rect 325923 379340 325924 379404
rect 325988 379340 325989 379404
rect 325923 379339 325989 379340
rect 303475 378996 303541 378997
rect 303475 378932 303476 378996
rect 303540 378932 303541 378996
rect 303475 378931 303541 378932
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 359308 301574 374058
rect 307794 364394 308414 379000
rect 307794 364158 307826 364394
rect 308062 364158 308146 364394
rect 308382 364158 308414 364394
rect 307794 364074 308414 364158
rect 307794 363838 307826 364074
rect 308062 363838 308146 364074
rect 308382 363838 308414 364074
rect 307794 359308 308414 363838
rect 311514 368114 312134 379000
rect 311514 367878 311546 368114
rect 311782 367878 311866 368114
rect 312102 367878 312134 368114
rect 311514 367794 312134 367878
rect 311514 367558 311546 367794
rect 311782 367558 311866 367794
rect 312102 367558 312134 367794
rect 311514 359308 312134 367558
rect 315234 369954 315854 379000
rect 315234 369718 315266 369954
rect 315502 369718 315586 369954
rect 315822 369718 315854 369954
rect 315234 369634 315854 369718
rect 315234 369398 315266 369634
rect 315502 369398 315586 369634
rect 315822 369398 315854 369634
rect 315234 359308 315854 369398
rect 318954 373674 319574 379000
rect 318954 373438 318986 373674
rect 319222 373438 319306 373674
rect 319542 373438 319574 373674
rect 318954 373354 319574 373438
rect 318954 373118 318986 373354
rect 319222 373118 319306 373354
rect 319542 373118 319574 373354
rect 318954 359308 319574 373118
rect 325794 363454 326414 379000
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 359308 326414 362898
rect 329514 367174 330134 379000
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 359308 330134 366618
rect 333234 370894 333854 379000
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 359308 333854 370338
rect 336954 374614 337574 379000
rect 343222 378997 343282 380430
rect 343406 379133 343466 380430
rect 343403 379132 343469 379133
rect 343403 379068 343404 379132
rect 343468 379068 343469 379132
rect 343403 379067 343469 379068
rect 343219 378996 343285 378997
rect 343219 378932 343220 378996
rect 343284 378932 343285 378996
rect 343219 378931 343285 378932
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 359308 337574 374058
rect 343794 364394 344414 379000
rect 343794 364158 343826 364394
rect 344062 364158 344146 364394
rect 344382 364158 344414 364394
rect 343794 364074 344414 364158
rect 343794 363838 343826 364074
rect 344062 363838 344146 364074
rect 344382 363838 344414 364074
rect 343794 359308 344414 363838
rect 347514 368114 348134 379000
rect 347514 367878 347546 368114
rect 347782 367878 347866 368114
rect 348102 367878 348134 368114
rect 347514 367794 348134 367878
rect 347514 367558 347546 367794
rect 347782 367558 347866 367794
rect 348102 367558 348134 367794
rect 347514 359308 348134 367558
rect 351234 369954 351854 379000
rect 351234 369718 351266 369954
rect 351502 369718 351586 369954
rect 351822 369718 351854 369954
rect 351234 369634 351854 369718
rect 351234 369398 351266 369634
rect 351502 369398 351586 369634
rect 351822 369398 351854 369634
rect 351234 359308 351854 369398
rect 354954 373674 355574 379000
rect 354954 373438 354986 373674
rect 355222 373438 355306 373674
rect 355542 373438 355574 373674
rect 354954 373354 355574 373438
rect 354954 373118 354986 373354
rect 355222 373118 355306 373354
rect 355542 373118 355574 373354
rect 354954 359308 355574 373118
rect 338435 358868 338501 358869
rect 338435 358804 338436 358868
rect 338500 358804 338501 358868
rect 338435 358803 338501 358804
rect 339723 358868 339789 358869
rect 339723 358804 339724 358868
rect 339788 358804 339789 358868
rect 339723 358803 339789 358804
rect 350947 358868 351013 358869
rect 350947 358804 350948 358868
rect 351012 358804 351013 358868
rect 350947 358803 351013 358804
rect 338438 358050 338498 358803
rect 339726 358050 339786 358803
rect 350950 358050 351010 358803
rect 338438 357990 338524 358050
rect 338464 357202 338524 357990
rect 339688 357990 339786 358050
rect 350840 357990 351010 358050
rect 339688 357202 339748 357990
rect 350840 357202 350900 357990
rect 220272 345454 220620 345486
rect 220272 345218 220328 345454
rect 220564 345218 220620 345454
rect 220272 345134 220620 345218
rect 220272 344898 220328 345134
rect 220564 344898 220620 345134
rect 220272 344866 220620 344898
rect 356000 345454 356348 345486
rect 356000 345218 356056 345454
rect 356292 345218 356348 345454
rect 356000 345134 356348 345218
rect 356000 344898 356056 345134
rect 356292 344898 356348 345134
rect 356000 344866 356348 344898
rect 220952 327454 221300 327486
rect 220952 327218 221008 327454
rect 221244 327218 221300 327454
rect 220952 327134 221300 327218
rect 220952 326898 221008 327134
rect 221244 326898 221300 327134
rect 220952 326866 221300 326898
rect 355320 327454 355668 327486
rect 355320 327218 355376 327454
rect 355612 327218 355668 327454
rect 355320 327134 355668 327218
rect 355320 326898 355376 327134
rect 355612 326898 355668 327134
rect 355320 326866 355668 326898
rect 220272 309454 220620 309486
rect 220272 309218 220328 309454
rect 220564 309218 220620 309454
rect 220272 309134 220620 309218
rect 220272 308898 220328 309134
rect 220564 308898 220620 309134
rect 220272 308866 220620 308898
rect 356000 309454 356348 309486
rect 356000 309218 356056 309454
rect 356292 309218 356348 309454
rect 356000 309134 356348 309218
rect 356000 308898 356056 309134
rect 356292 308898 356348 309134
rect 356000 308866 356348 308898
rect 220952 291454 221300 291486
rect 220952 291218 221008 291454
rect 221244 291218 221300 291454
rect 220952 291134 221300 291218
rect 220952 290898 221008 291134
rect 221244 290898 221300 291134
rect 220952 290866 221300 290898
rect 355320 291454 355668 291486
rect 355320 291218 355376 291454
rect 355612 291218 355668 291454
rect 355320 291134 355668 291218
rect 355320 290898 355376 291134
rect 355612 290898 355668 291134
rect 355320 290866 355668 290898
rect 236056 273730 236116 274040
rect 237144 273730 237204 274040
rect 238232 273730 238292 274040
rect 239592 273730 239652 274040
rect 235950 273670 236116 273730
rect 237054 273670 237204 273730
rect 238158 273670 238292 273730
rect 239262 273670 239652 273730
rect 240544 273730 240604 274040
rect 241768 273730 241828 274040
rect 243128 273730 243188 274040
rect 240544 273670 240610 273730
rect 235950 272237 236010 273670
rect 235947 272236 236013 272237
rect 235947 272172 235948 272236
rect 236012 272172 236013 272236
rect 235947 272171 236013 272172
rect 221514 259174 222134 272000
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221514 252308 222134 258618
rect 225234 262894 225854 272000
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 225234 252308 225854 262338
rect 228954 266614 229574 272000
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 228954 252308 229574 266058
rect 235794 256394 236414 272000
rect 237054 270605 237114 273670
rect 238158 270605 238218 273670
rect 239262 271149 239322 273670
rect 239259 271148 239325 271149
rect 239259 271084 239260 271148
rect 239324 271084 239325 271148
rect 239259 271083 239325 271084
rect 237051 270604 237117 270605
rect 237051 270540 237052 270604
rect 237116 270540 237117 270604
rect 237051 270539 237117 270540
rect 238155 270604 238221 270605
rect 238155 270540 238156 270604
rect 238220 270540 238221 270604
rect 238155 270539 238221 270540
rect 235794 256158 235826 256394
rect 236062 256158 236146 256394
rect 236382 256158 236414 256394
rect 235794 256074 236414 256158
rect 235794 255838 235826 256074
rect 236062 255838 236146 256074
rect 236382 255838 236414 256074
rect 235794 252308 236414 255838
rect 239514 260114 240134 272000
rect 240550 270197 240610 273670
rect 241654 273670 241828 273730
rect 242942 273670 243188 273730
rect 244216 273730 244276 274040
rect 245440 273730 245500 274040
rect 246528 273730 246588 274040
rect 244216 273670 244290 273730
rect 241654 270333 241714 273670
rect 242942 270605 243002 273670
rect 242939 270604 243005 270605
rect 242939 270540 242940 270604
rect 243004 270540 243005 270604
rect 242939 270539 243005 270540
rect 241651 270332 241717 270333
rect 241651 270268 241652 270332
rect 241716 270268 241717 270332
rect 241651 270267 241717 270268
rect 240547 270196 240613 270197
rect 240547 270132 240548 270196
rect 240612 270132 240613 270196
rect 240547 270131 240613 270132
rect 239514 259878 239546 260114
rect 239782 259878 239866 260114
rect 240102 259878 240134 260114
rect 239514 259794 240134 259878
rect 239514 259558 239546 259794
rect 239782 259558 239866 259794
rect 240102 259558 240134 259794
rect 239514 252308 240134 259558
rect 243234 261954 243854 272000
rect 244230 270605 244290 273670
rect 245334 273670 245500 273730
rect 246438 273670 246588 273730
rect 247616 273730 247676 274040
rect 248296 273730 248356 274040
rect 248704 273730 248764 274040
rect 247616 273670 247786 273730
rect 245334 270741 245394 273670
rect 245331 270740 245397 270741
rect 245331 270676 245332 270740
rect 245396 270676 245397 270740
rect 245331 270675 245397 270676
rect 246438 270605 246498 273670
rect 244227 270604 244293 270605
rect 244227 270540 244228 270604
rect 244292 270540 244293 270604
rect 244227 270539 244293 270540
rect 246435 270604 246501 270605
rect 246435 270540 246436 270604
rect 246500 270540 246501 270604
rect 246435 270539 246501 270540
rect 243234 261718 243266 261954
rect 243502 261718 243586 261954
rect 243822 261718 243854 261954
rect 243234 261634 243854 261718
rect 243234 261398 243266 261634
rect 243502 261398 243586 261634
rect 243822 261398 243854 261634
rect 243234 252308 243854 261398
rect 246954 265674 247574 272000
rect 247726 270605 247786 273670
rect 248278 273670 248356 273730
rect 248646 273670 248764 273730
rect 250064 273730 250124 274040
rect 250064 273670 250178 273730
rect 248278 271149 248338 273670
rect 248275 271148 248341 271149
rect 248275 271084 248276 271148
rect 248340 271084 248341 271148
rect 248275 271083 248341 271084
rect 248646 270605 248706 273670
rect 250118 270605 250178 273670
rect 250744 273597 250804 274040
rect 251288 273730 251348 274040
rect 252376 273730 252436 274040
rect 253464 273730 253524 274040
rect 251222 273670 251348 273730
rect 252326 273670 252436 273730
rect 253430 273670 253524 273730
rect 253600 273730 253660 274040
rect 254552 273730 254612 274040
rect 255912 273730 255972 274040
rect 253600 273670 253674 273730
rect 250741 273596 250807 273597
rect 250741 273532 250742 273596
rect 250806 273532 250807 273596
rect 250741 273531 250807 273532
rect 251222 270605 251282 273670
rect 252326 270741 252386 273670
rect 253430 270877 253490 273670
rect 253614 271149 253674 273670
rect 254534 273670 254612 273730
rect 255822 273670 255972 273730
rect 256048 273730 256108 274040
rect 257000 273730 257060 274040
rect 256048 273670 256250 273730
rect 253611 271148 253677 271149
rect 253611 271084 253612 271148
rect 253676 271084 253677 271148
rect 253611 271083 253677 271084
rect 253427 270876 253493 270877
rect 253427 270812 253428 270876
rect 253492 270812 253493 270876
rect 253427 270811 253493 270812
rect 252323 270740 252389 270741
rect 252323 270676 252324 270740
rect 252388 270676 252389 270740
rect 252323 270675 252389 270676
rect 247723 270604 247789 270605
rect 247723 270540 247724 270604
rect 247788 270540 247789 270604
rect 247723 270539 247789 270540
rect 248643 270604 248709 270605
rect 248643 270540 248644 270604
rect 248708 270540 248709 270604
rect 248643 270539 248709 270540
rect 250115 270604 250181 270605
rect 250115 270540 250116 270604
rect 250180 270540 250181 270604
rect 250115 270539 250181 270540
rect 251219 270604 251285 270605
rect 251219 270540 251220 270604
rect 251284 270540 251285 270604
rect 251219 270539 251285 270540
rect 246954 265438 246986 265674
rect 247222 265438 247306 265674
rect 247542 265438 247574 265674
rect 246954 265354 247574 265438
rect 246954 265118 246986 265354
rect 247222 265118 247306 265354
rect 247542 265118 247574 265354
rect 246954 252308 247574 265118
rect 253794 255454 254414 272000
rect 254534 270605 254594 273670
rect 255822 270605 255882 273670
rect 256190 271829 256250 273670
rect 256926 273670 257060 273730
rect 258088 273730 258148 274040
rect 258496 273730 258556 274040
rect 258088 273670 258274 273730
rect 256187 271828 256253 271829
rect 256187 271764 256188 271828
rect 256252 271764 256253 271828
rect 256187 271763 256253 271764
rect 256926 270605 256986 273670
rect 254531 270604 254597 270605
rect 254531 270540 254532 270604
rect 254596 270540 254597 270604
rect 254531 270539 254597 270540
rect 255819 270604 255885 270605
rect 255819 270540 255820 270604
rect 255884 270540 255885 270604
rect 255819 270539 255885 270540
rect 256923 270604 256989 270605
rect 256923 270540 256924 270604
rect 256988 270540 256989 270604
rect 256923 270539 256989 270540
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 252308 254414 254898
rect 257514 259174 258134 272000
rect 258214 271010 258274 273670
rect 258398 273670 258556 273730
rect 259448 273730 259508 274040
rect 260672 273730 260732 274040
rect 261080 273730 261140 274040
rect 259448 273670 259562 273730
rect 258398 271285 258458 273670
rect 258395 271284 258461 271285
rect 258395 271220 258396 271284
rect 258460 271220 258461 271284
rect 258395 271219 258461 271220
rect 258214 270950 258458 271010
rect 258398 270605 258458 270950
rect 259502 270605 259562 273670
rect 260606 273670 260732 273730
rect 260974 273670 261140 273730
rect 261760 273730 261820 274040
rect 262848 273730 262908 274040
rect 261760 273670 262138 273730
rect 260606 270741 260666 273670
rect 260974 271285 261034 273670
rect 260971 271284 261037 271285
rect 260971 271220 260972 271284
rect 261036 271220 261037 271284
rect 260971 271219 261037 271220
rect 260603 270740 260669 270741
rect 260603 270676 260604 270740
rect 260668 270676 260669 270740
rect 260603 270675 260669 270676
rect 258395 270604 258461 270605
rect 258395 270540 258396 270604
rect 258460 270540 258461 270604
rect 258395 270539 258461 270540
rect 259499 270604 259565 270605
rect 259499 270540 259500 270604
rect 259564 270540 259565 270604
rect 259499 270539 259565 270540
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 252308 258134 258618
rect 261234 262894 261854 272000
rect 262078 271149 262138 273670
rect 262814 273670 262908 273730
rect 263528 273730 263588 274040
rect 263936 273730 263996 274040
rect 263528 273670 263610 273730
rect 262075 271148 262141 271149
rect 262075 271084 262076 271148
rect 262140 271084 262141 271148
rect 262075 271083 262141 271084
rect 262814 270605 262874 273670
rect 263550 271829 263610 273670
rect 263918 273670 263996 273730
rect 265296 273730 265356 274040
rect 265976 273730 266036 274040
rect 266384 273730 266444 274040
rect 267608 273730 267668 274040
rect 265296 273670 265818 273730
rect 263547 271828 263613 271829
rect 263547 271764 263548 271828
rect 263612 271764 263613 271828
rect 263547 271763 263613 271764
rect 263918 270605 263978 273670
rect 262811 270604 262877 270605
rect 262811 270540 262812 270604
rect 262876 270540 262877 270604
rect 262811 270539 262877 270540
rect 263915 270604 263981 270605
rect 263915 270540 263916 270604
rect 263980 270540 263981 270604
rect 263915 270539 263981 270540
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 252308 261854 262338
rect 264954 266614 265574 272000
rect 265758 270877 265818 273670
rect 265942 273670 266036 273730
rect 266310 273670 266444 273730
rect 267598 273670 267668 273730
rect 268288 273730 268348 274040
rect 268696 273730 268756 274040
rect 269784 273730 269844 274040
rect 271008 273730 271068 274040
rect 268288 273670 268394 273730
rect 268696 273670 268762 273730
rect 269784 273670 269866 273730
rect 265942 271829 266002 273670
rect 265939 271828 266005 271829
rect 265939 271764 265940 271828
rect 266004 271764 266005 271828
rect 265939 271763 266005 271764
rect 266310 271149 266370 273670
rect 266307 271148 266373 271149
rect 266307 271084 266308 271148
rect 266372 271084 266373 271148
rect 266307 271083 266373 271084
rect 265755 270876 265821 270877
rect 265755 270812 265756 270876
rect 265820 270812 265821 270876
rect 265755 270811 265821 270812
rect 267598 270741 267658 273670
rect 268334 271829 268394 273670
rect 268331 271828 268397 271829
rect 268331 271764 268332 271828
rect 268396 271764 268397 271828
rect 268331 271763 268397 271764
rect 268702 271149 268762 273670
rect 268699 271148 268765 271149
rect 268699 271084 268700 271148
rect 268764 271084 268765 271148
rect 268699 271083 268765 271084
rect 267595 270740 267661 270741
rect 267595 270676 267596 270740
rect 267660 270676 267661 270740
rect 267595 270675 267661 270676
rect 269806 270605 269866 273670
rect 270910 273670 271068 273730
rect 271144 273730 271204 274040
rect 271144 273670 271338 273730
rect 270910 271829 270970 273670
rect 270907 271828 270973 271829
rect 270907 271764 270908 271828
rect 270972 271764 270973 271828
rect 270907 271763 270973 271764
rect 271278 271149 271338 273670
rect 272232 273597 272292 274040
rect 273320 273730 273380 274040
rect 273592 273730 273652 274040
rect 274408 273730 274468 274040
rect 275768 273730 275828 274040
rect 273302 273670 273380 273730
rect 273486 273670 273652 273730
rect 274406 273670 274468 273730
rect 275326 273670 275828 273730
rect 276040 273730 276100 274040
rect 276992 273730 277052 274040
rect 276040 273670 276306 273730
rect 272229 273596 272295 273597
rect 272229 273532 272230 273596
rect 272294 273532 272295 273596
rect 272229 273531 272295 273532
rect 273302 273461 273362 273670
rect 273299 273460 273365 273461
rect 273299 273396 273300 273460
rect 273364 273396 273365 273460
rect 273299 273395 273365 273396
rect 271275 271148 271341 271149
rect 271275 271084 271276 271148
rect 271340 271084 271341 271148
rect 271275 271083 271341 271084
rect 269803 270604 269869 270605
rect 269803 270540 269804 270604
rect 269868 270540 269869 270604
rect 269803 270539 269869 270540
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 252308 265574 266058
rect 271794 256394 272414 272000
rect 273486 271829 273546 273670
rect 273483 271828 273549 271829
rect 273483 271764 273484 271828
rect 273548 271764 273549 271828
rect 273483 271763 273549 271764
rect 274406 270605 274466 273670
rect 275326 271829 275386 273670
rect 275323 271828 275389 271829
rect 275323 271764 275324 271828
rect 275388 271764 275389 271828
rect 275323 271763 275389 271764
rect 274403 270604 274469 270605
rect 274403 270540 274404 270604
rect 274468 270540 274469 270604
rect 274403 270539 274469 270540
rect 271794 256158 271826 256394
rect 272062 256158 272146 256394
rect 272382 256158 272414 256394
rect 271794 256074 272414 256158
rect 271794 255838 271826 256074
rect 272062 255838 272146 256074
rect 272382 255838 272414 256074
rect 271794 252308 272414 255838
rect 275514 260114 276134 272000
rect 276246 271829 276306 273670
rect 276982 273670 277052 273730
rect 278080 273730 278140 274040
rect 278488 273730 278548 274040
rect 279168 273730 279228 274040
rect 278080 273670 278146 273730
rect 276982 271829 277042 273670
rect 278086 271829 278146 273670
rect 278454 273670 278548 273730
rect 279006 273670 279228 273730
rect 278454 272645 278514 273670
rect 278451 272644 278517 272645
rect 278451 272580 278452 272644
rect 278516 272580 278517 272644
rect 278451 272579 278517 272580
rect 276243 271828 276309 271829
rect 276243 271764 276244 271828
rect 276308 271764 276309 271828
rect 276243 271763 276309 271764
rect 276979 271828 277045 271829
rect 276979 271764 276980 271828
rect 277044 271764 277045 271828
rect 276979 271763 277045 271764
rect 278083 271828 278149 271829
rect 278083 271764 278084 271828
rect 278148 271764 278149 271828
rect 278083 271763 278149 271764
rect 279006 271285 279066 273670
rect 280936 273597 280996 274040
rect 283520 273730 283580 274040
rect 283422 273670 283580 273730
rect 285968 273730 286028 274040
rect 288280 273730 288340 274040
rect 291000 273730 291060 274040
rect 293448 273730 293508 274040
rect 285968 273670 286058 273730
rect 280933 273596 280999 273597
rect 280933 273532 280934 273596
rect 280998 273532 280999 273596
rect 280933 273531 280999 273532
rect 283422 272781 283482 273670
rect 283419 272780 283485 272781
rect 283419 272716 283420 272780
rect 283484 272716 283485 272780
rect 283419 272715 283485 272716
rect 285998 272645 286058 273670
rect 288206 273670 288340 273730
rect 290966 273670 291060 273730
rect 293358 273670 293508 273730
rect 295896 273730 295956 274040
rect 298480 273730 298540 274040
rect 300928 273730 300988 274040
rect 303512 273730 303572 274040
rect 305960 273730 306020 274040
rect 295896 273670 295994 273730
rect 298480 273670 298570 273730
rect 288206 272781 288266 273670
rect 290966 272781 291026 273670
rect 288203 272780 288269 272781
rect 288203 272716 288204 272780
rect 288268 272716 288269 272780
rect 288203 272715 288269 272716
rect 290963 272780 291029 272781
rect 290963 272716 290964 272780
rect 291028 272716 291029 272780
rect 290963 272715 291029 272716
rect 285995 272644 286061 272645
rect 285995 272580 285996 272644
rect 286060 272580 286061 272644
rect 285995 272579 286061 272580
rect 293358 272509 293418 273670
rect 295934 272781 295994 273670
rect 295931 272780 295997 272781
rect 295931 272716 295932 272780
rect 295996 272716 295997 272780
rect 295931 272715 295997 272716
rect 298510 272645 298570 273670
rect 300902 273670 300988 273730
rect 303478 273670 303572 273730
rect 305870 273670 306020 273730
rect 308544 273730 308604 274040
rect 310992 273730 311052 274040
rect 313440 273730 313500 274040
rect 315888 273730 315948 274040
rect 318472 273730 318532 274040
rect 308544 273670 308690 273730
rect 310992 273670 311082 273730
rect 300902 272645 300962 273670
rect 298507 272644 298573 272645
rect 298507 272580 298508 272644
rect 298572 272580 298573 272644
rect 298507 272579 298573 272580
rect 300899 272644 300965 272645
rect 300899 272580 300900 272644
rect 300964 272580 300965 272644
rect 300899 272579 300965 272580
rect 293355 272508 293421 272509
rect 293355 272444 293356 272508
rect 293420 272444 293421 272508
rect 293355 272443 293421 272444
rect 279003 271284 279069 271285
rect 279003 271220 279004 271284
rect 279068 271220 279069 271284
rect 279003 271219 279069 271220
rect 275514 259878 275546 260114
rect 275782 259878 275866 260114
rect 276102 259878 276134 260114
rect 275514 259794 276134 259878
rect 275514 259558 275546 259794
rect 275782 259558 275866 259794
rect 276102 259558 276134 259794
rect 275514 252308 276134 259558
rect 279234 261954 279854 272000
rect 279234 261718 279266 261954
rect 279502 261718 279586 261954
rect 279822 261718 279854 261954
rect 279234 261634 279854 261718
rect 279234 261398 279266 261634
rect 279502 261398 279586 261634
rect 279822 261398 279854 261634
rect 279234 252308 279854 261398
rect 282954 265674 283574 272000
rect 282954 265438 282986 265674
rect 283222 265438 283306 265674
rect 283542 265438 283574 265674
rect 282954 265354 283574 265438
rect 282954 265118 282986 265354
rect 283222 265118 283306 265354
rect 283542 265118 283574 265354
rect 282954 252308 283574 265118
rect 289794 255454 290414 272000
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 252308 290414 254898
rect 293514 259174 294134 272000
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 252308 294134 258618
rect 297234 262894 297854 272000
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 252308 297854 262338
rect 300954 266614 301574 272000
rect 303478 271829 303538 273670
rect 305870 272917 305930 273670
rect 305867 272916 305933 272917
rect 305867 272852 305868 272916
rect 305932 272852 305933 272916
rect 305867 272851 305933 272852
rect 303475 271828 303541 271829
rect 303475 271764 303476 271828
rect 303540 271764 303541 271828
rect 303475 271763 303541 271764
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 252308 301574 266058
rect 307794 256394 308414 272000
rect 308630 271829 308690 273670
rect 311022 273053 311082 273670
rect 313414 273670 313500 273730
rect 315070 273670 315948 273730
rect 318382 273670 318532 273730
rect 320920 273730 320980 274040
rect 323368 273730 323428 274040
rect 325952 273730 326012 274040
rect 343224 273730 343284 274040
rect 320920 273670 321018 273730
rect 311019 273052 311085 273053
rect 311019 272988 311020 273052
rect 311084 272988 311085 273052
rect 311019 272987 311085 272988
rect 308627 271828 308693 271829
rect 308627 271764 308628 271828
rect 308692 271764 308693 271828
rect 308627 271763 308693 271764
rect 307794 256158 307826 256394
rect 308062 256158 308146 256394
rect 308382 256158 308414 256394
rect 307794 256074 308414 256158
rect 307794 255838 307826 256074
rect 308062 255838 308146 256074
rect 308382 255838 308414 256074
rect 307794 252308 308414 255838
rect 311514 260114 312134 272000
rect 313414 271421 313474 273670
rect 315070 271557 315130 273670
rect 318382 273189 318442 273670
rect 318379 273188 318445 273189
rect 318379 273124 318380 273188
rect 318444 273124 318445 273188
rect 318379 273123 318445 273124
rect 315067 271556 315133 271557
rect 315067 271492 315068 271556
rect 315132 271492 315133 271556
rect 315067 271491 315133 271492
rect 313411 271420 313477 271421
rect 313411 271356 313412 271420
rect 313476 271356 313477 271420
rect 313411 271355 313477 271356
rect 311514 259878 311546 260114
rect 311782 259878 311866 260114
rect 312102 259878 312134 260114
rect 311514 259794 312134 259878
rect 311514 259558 311546 259794
rect 311782 259558 311866 259794
rect 312102 259558 312134 259794
rect 311514 252308 312134 259558
rect 315234 261954 315854 272000
rect 315234 261718 315266 261954
rect 315502 261718 315586 261954
rect 315822 261718 315854 261954
rect 315234 261634 315854 261718
rect 315234 261398 315266 261634
rect 315502 261398 315586 261634
rect 315822 261398 315854 261634
rect 315234 252308 315854 261398
rect 318954 265674 319574 272000
rect 320958 271013 321018 273670
rect 323350 273670 323428 273730
rect 325742 273670 326012 273730
rect 343222 273670 343284 273730
rect 343360 273730 343420 274040
rect 343360 273670 343466 273730
rect 320955 271012 321021 271013
rect 320955 270948 320956 271012
rect 321020 270948 321021 271012
rect 320955 270947 321021 270948
rect 323350 270469 323410 273670
rect 325742 272370 325802 273670
rect 325558 272310 325802 272370
rect 325558 271693 325618 272310
rect 325555 271692 325621 271693
rect 325555 271628 325556 271692
rect 325620 271628 325621 271692
rect 325555 271627 325621 271628
rect 323347 270468 323413 270469
rect 323347 270404 323348 270468
rect 323412 270404 323413 270468
rect 323347 270403 323413 270404
rect 318954 265438 318986 265674
rect 319222 265438 319306 265674
rect 319542 265438 319574 265674
rect 318954 265354 319574 265438
rect 318954 265118 318986 265354
rect 319222 265118 319306 265354
rect 319542 265118 319574 265354
rect 318954 252308 319574 265118
rect 325794 255454 326414 272000
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 252308 326414 254898
rect 329514 259174 330134 272000
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 252308 330134 258618
rect 333234 262894 333854 272000
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 252308 333854 262338
rect 336954 266614 337574 272000
rect 343222 271693 343282 273670
rect 343219 271692 343285 271693
rect 343219 271628 343220 271692
rect 343284 271628 343285 271692
rect 343219 271627 343285 271628
rect 343406 271557 343466 273670
rect 343403 271556 343469 271557
rect 343403 271492 343404 271556
rect 343468 271492 343469 271556
rect 343403 271491 343469 271492
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 252308 337574 266058
rect 343794 256394 344414 272000
rect 343794 256158 343826 256394
rect 344062 256158 344146 256394
rect 344382 256158 344414 256394
rect 343794 256074 344414 256158
rect 343794 255838 343826 256074
rect 344062 255838 344146 256074
rect 344382 255838 344414 256074
rect 339723 253468 339789 253469
rect 339723 253404 339724 253468
rect 339788 253404 339789 253468
rect 339723 253403 339789 253404
rect 338435 253060 338501 253061
rect 338435 252996 338436 253060
rect 338500 252996 338501 253060
rect 338435 252995 338501 252996
rect 338438 250610 338498 252995
rect 339726 250610 339786 253403
rect 343794 252308 344414 255838
rect 347514 260114 348134 272000
rect 347514 259878 347546 260114
rect 347782 259878 347866 260114
rect 348102 259878 348134 260114
rect 347514 259794 348134 259878
rect 347514 259558 347546 259794
rect 347782 259558 347866 259794
rect 348102 259558 348134 259794
rect 347514 252308 348134 259558
rect 351234 261954 351854 272000
rect 351234 261718 351266 261954
rect 351502 261718 351586 261954
rect 351822 261718 351854 261954
rect 351234 261634 351854 261718
rect 351234 261398 351266 261634
rect 351502 261398 351586 261634
rect 351822 261398 351854 261634
rect 350947 253196 351013 253197
rect 350947 253132 350948 253196
rect 351012 253132 351013 253196
rect 350947 253131 351013 253132
rect 350950 250610 351010 253131
rect 351234 252308 351854 261398
rect 354954 265674 355574 272000
rect 354954 265438 354986 265674
rect 355222 265438 355306 265674
rect 355542 265438 355574 265674
rect 354954 265354 355574 265438
rect 354954 265118 354986 265354
rect 355222 265118 355306 265354
rect 355542 265118 355574 265354
rect 354954 252308 355574 265118
rect 338438 250550 338524 250610
rect 338464 250240 338524 250550
rect 339688 250550 339786 250610
rect 350840 250550 351010 250610
rect 339688 250240 339748 250550
rect 350840 250240 350900 250550
rect 220272 237454 220620 237486
rect 220272 237218 220328 237454
rect 220564 237218 220620 237454
rect 220272 237134 220620 237218
rect 220272 236898 220328 237134
rect 220564 236898 220620 237134
rect 220272 236866 220620 236898
rect 356000 237454 356348 237486
rect 356000 237218 356056 237454
rect 356292 237218 356348 237454
rect 356000 237134 356348 237218
rect 356000 236898 356056 237134
rect 356292 236898 356348 237134
rect 356000 236866 356348 236898
rect 220952 219454 221300 219486
rect 220952 219218 221008 219454
rect 221244 219218 221300 219454
rect 220952 219134 221300 219218
rect 220952 218898 221008 219134
rect 221244 218898 221300 219134
rect 220952 218866 221300 218898
rect 355320 219454 355668 219486
rect 355320 219218 355376 219454
rect 355612 219218 355668 219454
rect 355320 219134 355668 219218
rect 355320 218898 355376 219134
rect 355612 218898 355668 219134
rect 355320 218866 355668 218898
rect 220272 201454 220620 201486
rect 220272 201218 220328 201454
rect 220564 201218 220620 201454
rect 220272 201134 220620 201218
rect 220272 200898 220328 201134
rect 220564 200898 220620 201134
rect 220272 200866 220620 200898
rect 356000 201454 356348 201486
rect 356000 201218 356056 201454
rect 356292 201218 356348 201454
rect 356000 201134 356348 201218
rect 356000 200898 356056 201134
rect 356292 200898 356348 201134
rect 356000 200866 356348 200898
rect 220952 183454 221300 183486
rect 220952 183218 221008 183454
rect 221244 183218 221300 183454
rect 220952 183134 221300 183218
rect 220952 182898 221008 183134
rect 221244 182898 221300 183134
rect 220952 182866 221300 182898
rect 355320 183454 355668 183486
rect 355320 183218 355376 183454
rect 355612 183218 355668 183454
rect 355320 183134 355668 183218
rect 355320 182898 355376 183134
rect 355612 182898 355668 183134
rect 355320 182866 355668 182898
rect 219939 167108 220005 167109
rect 219939 167044 219940 167108
rect 220004 167044 220005 167108
rect 219939 167043 220005 167044
rect 236056 166290 236116 167106
rect 237144 166290 237204 167106
rect 238232 166290 238292 167106
rect 236056 166230 236194 166290
rect 236134 165613 236194 166230
rect 237054 166230 237204 166290
rect 238158 166230 238292 166290
rect 239592 166290 239652 167106
rect 240544 166290 240604 167106
rect 241768 166290 241828 167106
rect 243128 166290 243188 167106
rect 244216 167010 244276 167106
rect 245440 167010 245500 167106
rect 246528 167010 246588 167106
rect 247616 167010 247676 167106
rect 248296 167010 248356 167106
rect 248704 167010 248764 167106
rect 244216 166950 244474 167010
rect 244216 166910 244290 166950
rect 239592 166230 239690 166290
rect 240544 166230 240610 166290
rect 236131 165612 236197 165613
rect 236131 165548 236132 165612
rect 236196 165548 236197 165612
rect 236131 165547 236197 165548
rect 221514 151174 222134 165000
rect 221514 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 222134 151174
rect 221514 150854 222134 150938
rect 221514 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 222134 150854
rect 221514 145308 222134 150618
rect 225234 154894 225854 165000
rect 225234 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 225854 154894
rect 225234 154574 225854 154658
rect 225234 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 225854 154574
rect 225234 145308 225854 154338
rect 228954 158614 229574 165000
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228954 145308 229574 158058
rect 235794 148394 236414 165000
rect 237054 164253 237114 166230
rect 238158 164253 238218 166230
rect 239630 165613 239690 166230
rect 239627 165612 239693 165613
rect 239627 165548 239628 165612
rect 239692 165548 239693 165612
rect 239627 165547 239693 165548
rect 237051 164252 237117 164253
rect 237051 164188 237052 164252
rect 237116 164188 237117 164252
rect 237051 164187 237117 164188
rect 238155 164252 238221 164253
rect 238155 164188 238156 164252
rect 238220 164188 238221 164252
rect 238155 164187 238221 164188
rect 235794 148158 235826 148394
rect 236062 148158 236146 148394
rect 236382 148158 236414 148394
rect 235794 148074 236414 148158
rect 235794 147838 235826 148074
rect 236062 147838 236146 148074
rect 236382 147838 236414 148074
rect 235794 145308 236414 147838
rect 239514 152114 240134 165000
rect 240550 164253 240610 166230
rect 241654 166230 241828 166290
rect 243126 166230 243188 166290
rect 241654 164253 241714 166230
rect 243126 165613 243186 166230
rect 243123 165612 243189 165613
rect 243123 165548 243124 165612
rect 243188 165548 243189 165612
rect 243123 165547 243189 165548
rect 240547 164252 240613 164253
rect 240547 164188 240548 164252
rect 240612 164188 240613 164252
rect 240547 164187 240613 164188
rect 241651 164252 241717 164253
rect 241651 164188 241652 164252
rect 241716 164188 241717 164252
rect 241651 164187 241717 164188
rect 239514 151878 239546 152114
rect 239782 151878 239866 152114
rect 240102 151878 240134 152114
rect 239514 151794 240134 151878
rect 239514 151558 239546 151794
rect 239782 151558 239866 151794
rect 240102 151558 240134 151794
rect 239514 145308 240134 151558
rect 243234 155834 243854 165000
rect 244414 164389 244474 166950
rect 245334 166950 245500 167010
rect 246438 166950 246588 167010
rect 247542 166950 247676 167010
rect 248278 166950 248356 167010
rect 248646 166950 248764 167010
rect 250064 167010 250124 167106
rect 250744 167010 250804 167106
rect 251288 167010 251348 167106
rect 252376 167010 252436 167106
rect 253464 167010 253524 167106
rect 250064 166950 250178 167010
rect 244411 164388 244477 164389
rect 244411 164324 244412 164388
rect 244476 164324 244477 164388
rect 244411 164323 244477 164324
rect 245334 164253 245394 166950
rect 246438 164253 246498 166950
rect 247542 165613 247602 166950
rect 247539 165612 247605 165613
rect 247539 165548 247540 165612
rect 247604 165548 247605 165612
rect 247539 165547 247605 165548
rect 245331 164252 245397 164253
rect 245331 164188 245332 164252
rect 245396 164188 245397 164252
rect 245331 164187 245397 164188
rect 246435 164252 246501 164253
rect 246435 164188 246436 164252
rect 246500 164188 246501 164252
rect 246435 164187 246501 164188
rect 243234 155598 243266 155834
rect 243502 155598 243586 155834
rect 243822 155598 243854 155834
rect 243234 155514 243854 155598
rect 243234 155278 243266 155514
rect 243502 155278 243586 155514
rect 243822 155278 243854 155514
rect 243234 145308 243854 155278
rect 246954 157674 247574 165000
rect 248278 164933 248338 166950
rect 248275 164932 248341 164933
rect 248275 164868 248276 164932
rect 248340 164868 248341 164932
rect 248275 164867 248341 164868
rect 248646 164253 248706 166950
rect 250118 164253 250178 166950
rect 250670 166950 250804 167010
rect 251222 166950 251348 167010
rect 252326 166950 252436 167010
rect 253430 166950 253524 167010
rect 253600 167010 253660 167106
rect 254552 167010 254612 167106
rect 255912 167010 255972 167106
rect 253600 166950 253674 167010
rect 250670 164933 250730 166950
rect 250667 164932 250733 164933
rect 250667 164868 250668 164932
rect 250732 164868 250733 164932
rect 250667 164867 250733 164868
rect 251222 164253 251282 166950
rect 252326 164389 252386 166950
rect 252323 164388 252389 164389
rect 252323 164324 252324 164388
rect 252388 164324 252389 164388
rect 252323 164323 252389 164324
rect 253430 164253 253490 166950
rect 253614 166565 253674 166950
rect 254534 166950 254612 167010
rect 255822 166950 255972 167010
rect 256048 167010 256108 167106
rect 257000 167010 257060 167106
rect 258088 167010 258148 167106
rect 258496 167010 258556 167106
rect 256048 166950 256250 167010
rect 253611 166564 253677 166565
rect 253611 166500 253612 166564
rect 253676 166500 253677 166564
rect 253611 166499 253677 166500
rect 248643 164252 248709 164253
rect 248643 164188 248644 164252
rect 248708 164188 248709 164252
rect 248643 164187 248709 164188
rect 250115 164252 250181 164253
rect 250115 164188 250116 164252
rect 250180 164188 250181 164252
rect 250115 164187 250181 164188
rect 251219 164252 251285 164253
rect 251219 164188 251220 164252
rect 251284 164188 251285 164252
rect 251219 164187 251285 164188
rect 253427 164252 253493 164253
rect 253427 164188 253428 164252
rect 253492 164188 253493 164252
rect 253427 164187 253493 164188
rect 246954 157438 246986 157674
rect 247222 157438 247306 157674
rect 247542 157438 247574 157674
rect 246954 157354 247574 157438
rect 246954 157118 246986 157354
rect 247222 157118 247306 157354
rect 247542 157118 247574 157354
rect 246954 145308 247574 157118
rect 253794 147454 254414 165000
rect 254534 164253 254594 166950
rect 255822 164253 255882 166950
rect 256190 164933 256250 166950
rect 256926 166950 257060 167010
rect 258030 166950 258148 167010
rect 258398 166950 258556 167010
rect 259448 167010 259508 167106
rect 260672 167010 260732 167106
rect 261080 167010 261140 167106
rect 261760 167010 261820 167106
rect 262848 167010 262908 167106
rect 259448 166950 259562 167010
rect 256187 164932 256253 164933
rect 256187 164868 256188 164932
rect 256252 164868 256253 164932
rect 256187 164867 256253 164868
rect 256926 164389 256986 166950
rect 258030 165613 258090 166950
rect 258027 165612 258093 165613
rect 258027 165548 258028 165612
rect 258092 165548 258093 165612
rect 258027 165547 258093 165548
rect 256923 164388 256989 164389
rect 256923 164324 256924 164388
rect 256988 164324 256989 164388
rect 256923 164323 256989 164324
rect 254531 164252 254597 164253
rect 254531 164188 254532 164252
rect 254596 164188 254597 164252
rect 254531 164187 254597 164188
rect 255819 164252 255885 164253
rect 255819 164188 255820 164252
rect 255884 164188 255885 164252
rect 255819 164187 255885 164188
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 145308 254414 146898
rect 257514 151174 258134 165000
rect 258398 164933 258458 166950
rect 258395 164932 258461 164933
rect 258395 164868 258396 164932
rect 258460 164868 258461 164932
rect 258395 164867 258461 164868
rect 259502 164253 259562 166950
rect 260606 166950 260732 167010
rect 260974 166950 261140 167010
rect 261710 166950 261820 167010
rect 262814 166950 262908 167010
rect 263528 167010 263588 167106
rect 263936 167010 263996 167106
rect 263528 166950 263794 167010
rect 260606 164389 260666 166950
rect 260974 165205 261034 166950
rect 261710 165613 261770 166950
rect 261707 165612 261773 165613
rect 261707 165548 261708 165612
rect 261772 165548 261773 165612
rect 261707 165547 261773 165548
rect 260971 165204 261037 165205
rect 260971 165140 260972 165204
rect 261036 165140 261037 165204
rect 260971 165139 261037 165140
rect 260603 164388 260669 164389
rect 260603 164324 260604 164388
rect 260668 164324 260669 164388
rect 260603 164323 260669 164324
rect 259499 164252 259565 164253
rect 259499 164188 259500 164252
rect 259564 164188 259565 164252
rect 259499 164187 259565 164188
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 145308 258134 150618
rect 261234 154894 261854 165000
rect 262814 164253 262874 166950
rect 263734 165205 263794 166950
rect 263918 166950 263996 167010
rect 265296 167010 265356 167106
rect 265976 167010 266036 167106
rect 266384 167010 266444 167106
rect 267608 167010 267668 167106
rect 265296 166950 265450 167010
rect 263731 165204 263797 165205
rect 263731 165140 263732 165204
rect 263796 165140 263797 165204
rect 263731 165139 263797 165140
rect 263918 164253 263978 166950
rect 265390 165205 265450 166950
rect 265942 166950 266036 167010
rect 266310 166950 266444 167010
rect 267598 166950 267668 167010
rect 268288 167010 268348 167106
rect 268696 167010 268756 167106
rect 269784 167010 269844 167106
rect 271008 167010 271068 167106
rect 268288 166950 268394 167010
rect 268696 166950 268762 167010
rect 269784 166950 269866 167010
rect 265942 166565 266002 166950
rect 265939 166564 266005 166565
rect 265939 166500 265940 166564
rect 266004 166500 266005 166564
rect 265939 166499 266005 166500
rect 265387 165204 265453 165205
rect 265387 165140 265388 165204
rect 265452 165140 265453 165204
rect 265387 165139 265453 165140
rect 262811 164252 262877 164253
rect 262811 164188 262812 164252
rect 262876 164188 262877 164252
rect 262811 164187 262877 164188
rect 263915 164252 263981 164253
rect 263915 164188 263916 164252
rect 263980 164188 263981 164252
rect 263915 164187 263981 164188
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 145308 261854 154338
rect 264954 158614 265574 165000
rect 266310 164253 266370 166950
rect 267598 164389 267658 166950
rect 268334 165069 268394 166950
rect 268331 165068 268397 165069
rect 268331 165004 268332 165068
rect 268396 165004 268397 165068
rect 268331 165003 268397 165004
rect 267595 164388 267661 164389
rect 267595 164324 267596 164388
rect 267660 164324 267661 164388
rect 267595 164323 267661 164324
rect 268702 164253 268762 166950
rect 269806 164253 269866 166950
rect 270910 166950 271068 167010
rect 271144 167010 271204 167106
rect 272232 167010 272292 167106
rect 271144 166950 271338 167010
rect 270910 166565 270970 166950
rect 270907 166564 270973 166565
rect 270907 166500 270908 166564
rect 270972 166500 270973 166564
rect 270907 166499 270973 166500
rect 271278 164253 271338 166950
rect 272198 166950 272292 167010
rect 272198 165205 272258 166950
rect 273320 166290 273380 167106
rect 273592 166290 273652 167106
rect 274408 166290 274468 167106
rect 275768 166290 275828 167106
rect 273302 166230 273380 166290
rect 273486 166230 273652 166290
rect 274406 166230 274468 166290
rect 275694 166230 275828 166290
rect 276040 166290 276100 167106
rect 276992 166290 277052 167106
rect 276040 166230 276122 166290
rect 272195 165204 272261 165205
rect 272195 165140 272196 165204
rect 272260 165140 272261 165204
rect 272195 165139 272261 165140
rect 266307 164252 266373 164253
rect 266307 164188 266308 164252
rect 266372 164188 266373 164252
rect 266307 164187 266373 164188
rect 268699 164252 268765 164253
rect 268699 164188 268700 164252
rect 268764 164188 268765 164252
rect 268699 164187 268765 164188
rect 269803 164252 269869 164253
rect 269803 164188 269804 164252
rect 269868 164188 269869 164252
rect 269803 164187 269869 164188
rect 271275 164252 271341 164253
rect 271275 164188 271276 164252
rect 271340 164188 271341 164252
rect 271275 164187 271341 164188
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 145308 265574 158058
rect 271794 148394 272414 165000
rect 273302 164253 273362 166230
rect 273486 165613 273546 166230
rect 273483 165612 273549 165613
rect 273483 165548 273484 165612
rect 273548 165548 273549 165612
rect 273483 165547 273549 165548
rect 274406 164389 274466 166230
rect 275694 165205 275754 166230
rect 276062 165613 276122 166230
rect 276982 166230 277052 166290
rect 278080 166290 278140 167106
rect 278488 166290 278548 167106
rect 278080 166230 278146 166290
rect 276059 165612 276125 165613
rect 276059 165548 276060 165612
rect 276124 165548 276125 165612
rect 276059 165547 276125 165548
rect 275691 165204 275757 165205
rect 275691 165140 275692 165204
rect 275756 165140 275757 165204
rect 275691 165139 275757 165140
rect 274403 164388 274469 164389
rect 274403 164324 274404 164388
rect 274468 164324 274469 164388
rect 274403 164323 274469 164324
rect 273299 164252 273365 164253
rect 273299 164188 273300 164252
rect 273364 164188 273365 164252
rect 273299 164187 273365 164188
rect 271794 148158 271826 148394
rect 272062 148158 272146 148394
rect 272382 148158 272414 148394
rect 271794 148074 272414 148158
rect 271794 147838 271826 148074
rect 272062 147838 272146 148074
rect 272382 147838 272414 148074
rect 271794 145308 272414 147838
rect 275514 152114 276134 165000
rect 276982 164253 277042 166230
rect 278086 164253 278146 166230
rect 278454 166230 278548 166290
rect 279168 166290 279228 167106
rect 280936 166290 280996 167106
rect 283520 166290 283580 167106
rect 279168 166230 279250 166290
rect 278454 165613 278514 166230
rect 278451 165612 278517 165613
rect 278451 165548 278452 165612
rect 278516 165548 278517 165612
rect 278451 165547 278517 165548
rect 279190 165205 279250 166230
rect 280846 166230 280996 166290
rect 283422 166230 283580 166290
rect 285968 166290 286028 167106
rect 288280 166701 288340 167106
rect 288277 166700 288343 166701
rect 288277 166636 288278 166700
rect 288342 166636 288343 166700
rect 288277 166635 288343 166636
rect 291000 166565 291060 167106
rect 290997 166564 291063 166565
rect 290997 166500 290998 166564
rect 291062 166500 291063 166564
rect 290997 166499 291063 166500
rect 293448 166290 293508 167106
rect 295896 166701 295956 167106
rect 298480 166837 298540 167106
rect 298477 166836 298543 166837
rect 298477 166772 298478 166836
rect 298542 166772 298543 166836
rect 298477 166771 298543 166772
rect 295893 166700 295959 166701
rect 295893 166636 295894 166700
rect 295958 166636 295959 166700
rect 295893 166635 295959 166636
rect 300928 166290 300988 167106
rect 303512 166837 303572 167106
rect 303509 166836 303575 166837
rect 303509 166772 303510 166836
rect 303574 166772 303575 166836
rect 303509 166771 303575 166772
rect 305960 166701 306020 167106
rect 308544 166701 308604 167106
rect 310992 166834 311052 167106
rect 313440 166837 313500 167106
rect 313437 166836 313503 166837
rect 310992 166774 311082 166834
rect 305957 166700 306023 166701
rect 305957 166636 305958 166700
rect 306022 166636 306023 166700
rect 305957 166635 306023 166636
rect 308541 166700 308607 166701
rect 308541 166636 308542 166700
rect 308606 166636 308607 166700
rect 308541 166635 308607 166636
rect 285968 166230 286058 166290
rect 280846 165613 280906 166230
rect 280843 165612 280909 165613
rect 280843 165548 280844 165612
rect 280908 165548 280909 165612
rect 280843 165547 280909 165548
rect 283422 165341 283482 166230
rect 285998 165613 286058 166230
rect 293358 166230 293508 166290
rect 300902 166230 300988 166290
rect 293358 165613 293418 166230
rect 300902 165613 300962 166230
rect 311022 165613 311082 166774
rect 313437 166772 313438 166836
rect 313502 166772 313503 166836
rect 313437 166771 313503 166772
rect 315888 166701 315948 167106
rect 315885 166700 315951 166701
rect 315885 166636 315886 166700
rect 315950 166636 315951 166700
rect 318472 166698 318532 167106
rect 315885 166635 315951 166636
rect 318382 166638 318532 166698
rect 320920 166698 320980 167106
rect 323368 166698 323428 167106
rect 320920 166638 321018 166698
rect 285995 165612 286061 165613
rect 285995 165548 285996 165612
rect 286060 165548 286061 165612
rect 285995 165547 286061 165548
rect 293355 165612 293421 165613
rect 293355 165548 293356 165612
rect 293420 165548 293421 165612
rect 293355 165547 293421 165548
rect 300899 165612 300965 165613
rect 300899 165548 300900 165612
rect 300964 165548 300965 165612
rect 300899 165547 300965 165548
rect 311019 165612 311085 165613
rect 311019 165548 311020 165612
rect 311084 165548 311085 165612
rect 311019 165547 311085 165548
rect 318382 165477 318442 166638
rect 318379 165476 318445 165477
rect 318379 165412 318380 165476
rect 318444 165412 318445 165476
rect 318379 165411 318445 165412
rect 283419 165340 283485 165341
rect 283419 165276 283420 165340
rect 283484 165276 283485 165340
rect 283419 165275 283485 165276
rect 279187 165204 279253 165205
rect 279187 165140 279188 165204
rect 279252 165140 279253 165204
rect 279187 165139 279253 165140
rect 276979 164252 277045 164253
rect 276979 164188 276980 164252
rect 277044 164188 277045 164252
rect 276979 164187 277045 164188
rect 278083 164252 278149 164253
rect 278083 164188 278084 164252
rect 278148 164188 278149 164252
rect 278083 164187 278149 164188
rect 275514 151878 275546 152114
rect 275782 151878 275866 152114
rect 276102 151878 276134 152114
rect 275514 151794 276134 151878
rect 275514 151558 275546 151794
rect 275782 151558 275866 151794
rect 276102 151558 276134 151794
rect 275514 145308 276134 151558
rect 279234 155834 279854 165000
rect 279234 155598 279266 155834
rect 279502 155598 279586 155834
rect 279822 155598 279854 155834
rect 279234 155514 279854 155598
rect 279234 155278 279266 155514
rect 279502 155278 279586 155514
rect 279822 155278 279854 155514
rect 279234 145308 279854 155278
rect 282954 157674 283574 165000
rect 282954 157438 282986 157674
rect 283222 157438 283306 157674
rect 283542 157438 283574 157674
rect 282954 157354 283574 157438
rect 282954 157118 282986 157354
rect 283222 157118 283306 157354
rect 283542 157118 283574 157354
rect 282954 145308 283574 157118
rect 289794 147454 290414 165000
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 145308 290414 146898
rect 293514 151174 294134 165000
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 145308 294134 150618
rect 297234 154894 297854 165000
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 145308 297854 154338
rect 300954 158614 301574 165000
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 145308 301574 158058
rect 307794 148394 308414 165000
rect 307794 148158 307826 148394
rect 308062 148158 308146 148394
rect 308382 148158 308414 148394
rect 307794 148074 308414 148158
rect 307794 147838 307826 148074
rect 308062 147838 308146 148074
rect 308382 147838 308414 148074
rect 307794 145308 308414 147838
rect 311514 152114 312134 165000
rect 311514 151878 311546 152114
rect 311782 151878 311866 152114
rect 312102 151878 312134 152114
rect 311514 151794 312134 151878
rect 311514 151558 311546 151794
rect 311782 151558 311866 151794
rect 312102 151558 312134 151794
rect 311514 145308 312134 151558
rect 315234 155834 315854 165000
rect 315234 155598 315266 155834
rect 315502 155598 315586 155834
rect 315822 155598 315854 155834
rect 315234 155514 315854 155598
rect 315234 155278 315266 155514
rect 315502 155278 315586 155514
rect 315822 155278 315854 155514
rect 315234 145308 315854 155278
rect 318954 157674 319574 165000
rect 320958 163981 321018 166638
rect 323350 166638 323428 166698
rect 323350 164797 323410 166638
rect 325952 166290 326012 167106
rect 343224 166290 343284 167106
rect 325926 166230 326012 166290
rect 343222 166230 343284 166290
rect 343360 166290 343420 167106
rect 343360 166230 343466 166290
rect 325926 165613 325986 166230
rect 343222 165613 343282 166230
rect 325923 165612 325989 165613
rect 325923 165548 325924 165612
rect 325988 165548 325989 165612
rect 325923 165547 325989 165548
rect 343219 165612 343285 165613
rect 343219 165548 343220 165612
rect 343284 165548 343285 165612
rect 343219 165547 343285 165548
rect 323347 164796 323413 164797
rect 323347 164732 323348 164796
rect 323412 164732 323413 164796
rect 323347 164731 323413 164732
rect 320955 163980 321021 163981
rect 320955 163916 320956 163980
rect 321020 163916 321021 163980
rect 320955 163915 321021 163916
rect 318954 157438 318986 157674
rect 319222 157438 319306 157674
rect 319542 157438 319574 157674
rect 318954 157354 319574 157438
rect 318954 157118 318986 157354
rect 319222 157118 319306 157354
rect 319542 157118 319574 157354
rect 318954 145308 319574 157118
rect 325794 147454 326414 165000
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 145308 326414 146898
rect 329514 151174 330134 165000
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 145308 330134 150618
rect 333234 154894 333854 165000
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 145308 333854 154338
rect 336954 158614 337574 165000
rect 343406 164933 343466 166230
rect 343403 164932 343469 164933
rect 343403 164868 343404 164932
rect 343468 164868 343469 164932
rect 343403 164867 343469 164868
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 145308 337574 158058
rect 343794 148394 344414 165000
rect 343794 148158 343826 148394
rect 344062 148158 344146 148394
rect 344382 148158 344414 148394
rect 343794 148074 344414 148158
rect 343794 147838 343826 148074
rect 344062 147838 344146 148074
rect 344382 147838 344414 148074
rect 343794 145308 344414 147838
rect 347514 152114 348134 165000
rect 347514 151878 347546 152114
rect 347782 151878 347866 152114
rect 348102 151878 348134 152114
rect 347514 151794 348134 151878
rect 347514 151558 347546 151794
rect 347782 151558 347866 151794
rect 348102 151558 348134 151794
rect 347514 145308 348134 151558
rect 351234 155834 351854 165000
rect 351234 155598 351266 155834
rect 351502 155598 351586 155834
rect 351822 155598 351854 155834
rect 351234 155514 351854 155598
rect 351234 155278 351266 155514
rect 351502 155278 351586 155514
rect 351822 155278 351854 155514
rect 351234 145308 351854 155278
rect 354954 157674 355574 165000
rect 354954 157438 354986 157674
rect 355222 157438 355306 157674
rect 355542 157438 355574 157674
rect 354954 157354 355574 157438
rect 354954 157118 354986 157354
rect 355222 157118 355306 157354
rect 355542 157118 355574 157354
rect 354954 145308 355574 157118
rect 338435 144940 338501 144941
rect 338435 144876 338436 144940
rect 338500 144876 338501 144940
rect 338435 144875 338501 144876
rect 339723 144940 339789 144941
rect 339723 144876 339724 144940
rect 339788 144876 339789 144940
rect 339723 144875 339789 144876
rect 350947 144940 351013 144941
rect 350947 144876 350948 144940
rect 351012 144876 351013 144940
rect 350947 144875 351013 144876
rect 338438 143850 338498 144875
rect 339726 143850 339786 144875
rect 350950 143850 351010 144875
rect 338438 143790 338524 143850
rect 338464 143202 338524 143790
rect 339688 143790 339786 143850
rect 350840 143790 351010 143850
rect 339688 143202 339748 143790
rect 350840 143202 350900 143790
rect 220272 129454 220620 129486
rect 220272 129218 220328 129454
rect 220564 129218 220620 129454
rect 220272 129134 220620 129218
rect 220272 128898 220328 129134
rect 220564 128898 220620 129134
rect 220272 128866 220620 128898
rect 356000 129454 356348 129486
rect 356000 129218 356056 129454
rect 356292 129218 356348 129454
rect 356000 129134 356348 129218
rect 356000 128898 356056 129134
rect 356292 128898 356348 129134
rect 356000 128866 356348 128898
rect 220952 111454 221300 111486
rect 220952 111218 221008 111454
rect 221244 111218 221300 111454
rect 220952 111134 221300 111218
rect 220952 110898 221008 111134
rect 221244 110898 221300 111134
rect 220952 110866 221300 110898
rect 355320 111454 355668 111486
rect 355320 111218 355376 111454
rect 355612 111218 355668 111454
rect 355320 111134 355668 111218
rect 355320 110898 355376 111134
rect 355612 110898 355668 111134
rect 355320 110866 355668 110898
rect 220272 93454 220620 93486
rect 220272 93218 220328 93454
rect 220564 93218 220620 93454
rect 220272 93134 220620 93218
rect 220272 92898 220328 93134
rect 220564 92898 220620 93134
rect 220272 92866 220620 92898
rect 356000 93454 356348 93486
rect 356000 93218 356056 93454
rect 356292 93218 356348 93454
rect 356000 93134 356348 93218
rect 356000 92898 356056 93134
rect 356292 92898 356348 93134
rect 356000 92866 356348 92898
rect 220952 75454 221300 75486
rect 220952 75218 221008 75454
rect 221244 75218 221300 75454
rect 220952 75134 221300 75218
rect 220952 74898 221008 75134
rect 221244 74898 221300 75134
rect 220952 74866 221300 74898
rect 355320 75454 355668 75486
rect 355320 75218 355376 75454
rect 355612 75218 355668 75454
rect 355320 75134 355668 75218
rect 355320 74898 355376 75134
rect 355612 74898 355668 75134
rect 355320 74866 355668 74898
rect 236056 59530 236116 60106
rect 237144 59530 237204 60106
rect 238232 59530 238292 60106
rect 239592 59530 239652 60106
rect 236056 59470 236194 59530
rect 219203 58580 219269 58581
rect 219203 58516 219204 58580
rect 219268 58516 219269 58580
rect 219203 58515 219269 58516
rect 217547 58444 217613 58445
rect 217547 58380 217548 58444
rect 217612 58380 217613 58444
rect 217547 58379 217613 58380
rect 236134 58173 236194 59470
rect 237054 59470 237204 59530
rect 238158 59470 238292 59530
rect 239262 59470 239652 59530
rect 240544 59530 240604 60106
rect 241768 59530 241828 60106
rect 243128 59530 243188 60106
rect 240544 59470 240610 59530
rect 236131 58172 236197 58173
rect 236131 58108 236132 58172
rect 236196 58108 236197 58172
rect 236131 58107 236197 58108
rect 217363 55044 217429 55045
rect 217363 54980 217364 55044
rect 217428 54980 217429 55044
rect 217363 54979 217429 54980
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 210371 3772 210437 3773
rect 210371 3708 210372 3772
rect 210436 3708 210437 3772
rect 210371 3707 210437 3708
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 39454 218414 58000
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 43174 222134 58000
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 46894 225854 58000
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 50614 229574 58000
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 57454 236414 58000
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 237054 56949 237114 59470
rect 238158 57901 238218 59470
rect 239262 57901 239322 59470
rect 238155 57900 238221 57901
rect 238155 57836 238156 57900
rect 238220 57836 238221 57900
rect 238155 57835 238221 57836
rect 239259 57900 239325 57901
rect 239259 57836 239260 57900
rect 239324 57836 239325 57900
rect 239259 57835 239325 57836
rect 235794 21454 236414 56898
rect 237051 56948 237117 56949
rect 237051 56884 237052 56948
rect 237116 56884 237117 56948
rect 237051 56883 237117 56884
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 25174 240134 58000
rect 240550 57901 240610 59470
rect 241654 59470 241828 59530
rect 242942 59470 243188 59530
rect 244216 59530 244276 60106
rect 245440 59530 245500 60106
rect 246528 59530 246588 60106
rect 244216 59470 244290 59530
rect 241654 57901 241714 59470
rect 242942 57901 243002 59470
rect 240547 57900 240613 57901
rect 240547 57836 240548 57900
rect 240612 57836 240613 57900
rect 240547 57835 240613 57836
rect 241651 57900 241717 57901
rect 241651 57836 241652 57900
rect 241716 57836 241717 57900
rect 241651 57835 241717 57836
rect 242939 57900 243005 57901
rect 242939 57836 242940 57900
rect 243004 57836 243005 57900
rect 242939 57835 243005 57836
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 28894 243854 58000
rect 244230 57901 244290 59470
rect 245334 59470 245500 59530
rect 246438 59470 246588 59530
rect 247616 59530 247676 60106
rect 248296 59530 248356 60106
rect 248704 59530 248764 60106
rect 247616 59470 247786 59530
rect 245334 57901 245394 59470
rect 246438 57901 246498 59470
rect 244227 57900 244293 57901
rect 244227 57836 244228 57900
rect 244292 57836 244293 57900
rect 244227 57835 244293 57836
rect 245331 57900 245397 57901
rect 245331 57836 245332 57900
rect 245396 57836 245397 57900
rect 245331 57835 245397 57836
rect 246435 57900 246501 57901
rect 246435 57836 246436 57900
rect 246500 57836 246501 57900
rect 246435 57835 246501 57836
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 32614 247574 58000
rect 247726 57901 247786 59470
rect 248278 59470 248356 59530
rect 248646 59470 248764 59530
rect 250064 59530 250124 60106
rect 250744 59530 250804 60106
rect 251288 59530 251348 60106
rect 252376 59530 252436 60106
rect 253464 59530 253524 60106
rect 250064 59470 250178 59530
rect 248278 57901 248338 59470
rect 248646 57901 248706 59470
rect 250118 57901 250178 59470
rect 250670 59470 250804 59530
rect 251222 59470 251348 59530
rect 252326 59470 252436 59530
rect 253430 59470 253524 59530
rect 253600 59530 253660 60106
rect 254552 59530 254612 60106
rect 255912 59805 255972 60106
rect 255909 59804 255975 59805
rect 255909 59740 255910 59804
rect 255974 59740 255975 59804
rect 255909 59739 255975 59740
rect 256048 59530 256108 60106
rect 257000 59669 257060 60106
rect 256997 59668 257063 59669
rect 256997 59604 256998 59668
rect 257062 59604 257063 59668
rect 256997 59603 257063 59604
rect 258088 59530 258148 60106
rect 258496 59669 258556 60106
rect 258493 59668 258559 59669
rect 258493 59604 258494 59668
rect 258558 59604 258559 59668
rect 258493 59603 258559 59604
rect 253600 59470 253674 59530
rect 250670 58717 250730 59470
rect 250667 58716 250733 58717
rect 250667 58652 250668 58716
rect 250732 58652 250733 58716
rect 250667 58651 250733 58652
rect 251222 57901 251282 59470
rect 252326 57901 252386 59470
rect 253430 57901 253490 59470
rect 247723 57900 247789 57901
rect 247723 57836 247724 57900
rect 247788 57836 247789 57900
rect 247723 57835 247789 57836
rect 248275 57900 248341 57901
rect 248275 57836 248276 57900
rect 248340 57836 248341 57900
rect 248275 57835 248341 57836
rect 248643 57900 248709 57901
rect 248643 57836 248644 57900
rect 248708 57836 248709 57900
rect 248643 57835 248709 57836
rect 250115 57900 250181 57901
rect 250115 57836 250116 57900
rect 250180 57836 250181 57900
rect 250115 57835 250181 57836
rect 251219 57900 251285 57901
rect 251219 57836 251220 57900
rect 251284 57836 251285 57900
rect 251219 57835 251285 57836
rect 252323 57900 252389 57901
rect 252323 57836 252324 57900
rect 252388 57836 252389 57900
rect 252323 57835 252389 57836
rect 253427 57900 253493 57901
rect 253427 57836 253428 57900
rect 253492 57836 253493 57900
rect 253427 57835 253493 57836
rect 253614 57085 253674 59470
rect 254534 59470 254612 59530
rect 256006 59470 256108 59530
rect 257846 59470 258148 59530
rect 259448 59530 259508 60106
rect 260672 59805 260732 60106
rect 260669 59804 260735 59805
rect 260669 59740 260670 59804
rect 260734 59740 260735 59804
rect 260669 59739 260735 59740
rect 261080 59530 261140 60106
rect 261760 59805 261820 60106
rect 262848 59805 262908 60106
rect 261757 59804 261823 59805
rect 261757 59740 261758 59804
rect 261822 59740 261823 59804
rect 261757 59739 261823 59740
rect 262845 59804 262911 59805
rect 262845 59740 262846 59804
rect 262910 59740 262911 59804
rect 262845 59739 262911 59740
rect 259448 59470 259562 59530
rect 253611 57084 253677 57085
rect 253611 57020 253612 57084
rect 253676 57020 253677 57084
rect 253611 57019 253677 57020
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 39454 254414 58000
rect 254534 57901 254594 59470
rect 254531 57900 254597 57901
rect 254531 57836 254532 57900
rect 254596 57836 254597 57900
rect 254531 57835 254597 57836
rect 256006 57221 256066 59470
rect 257846 58445 257906 59470
rect 259502 59397 259562 59470
rect 260974 59470 261140 59530
rect 263528 59530 263588 60106
rect 263936 59805 263996 60106
rect 263933 59804 263999 59805
rect 263933 59740 263934 59804
rect 263998 59740 263999 59804
rect 263933 59739 263999 59740
rect 265296 59530 265356 60106
rect 265976 59530 266036 60106
rect 266384 59530 266444 60106
rect 267608 59530 267668 60106
rect 263528 59470 263610 59530
rect 259499 59396 259565 59397
rect 259499 59332 259500 59396
rect 259564 59332 259565 59396
rect 259499 59331 259565 59332
rect 257843 58444 257909 58445
rect 257843 58380 257844 58444
rect 257908 58380 257909 58444
rect 257843 58379 257909 58380
rect 256003 57220 256069 57221
rect 256003 57156 256004 57220
rect 256068 57156 256069 57220
rect 256003 57155 256069 57156
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 43174 258134 58000
rect 260974 57357 261034 59470
rect 260971 57356 261037 57357
rect 260971 57292 260972 57356
rect 261036 57292 261037 57356
rect 260971 57291 261037 57292
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 46894 261854 58000
rect 263550 57765 263610 59470
rect 265206 59470 265356 59530
rect 265942 59470 266036 59530
rect 266310 59470 266444 59530
rect 267598 59470 267668 59530
rect 268288 59530 268348 60106
rect 268696 59530 268756 60106
rect 269784 59530 269844 60106
rect 271008 59530 271068 60106
rect 268288 59470 268394 59530
rect 268696 59470 268762 59530
rect 269784 59470 269866 59530
rect 265206 58581 265266 59470
rect 265203 58580 265269 58581
rect 265203 58516 265204 58580
rect 265268 58516 265269 58580
rect 265203 58515 265269 58516
rect 263547 57764 263613 57765
rect 263547 57700 263548 57764
rect 263612 57700 263613 57764
rect 263547 57699 263613 57700
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 50614 265574 58000
rect 265942 57765 266002 59470
rect 265939 57764 266005 57765
rect 265939 57700 265940 57764
rect 266004 57700 266005 57764
rect 265939 57699 266005 57700
rect 266310 57357 266370 59470
rect 267598 57765 267658 59470
rect 268334 57765 268394 59470
rect 268702 57765 268762 59470
rect 269806 57765 269866 59470
rect 270910 59470 271068 59530
rect 271144 59530 271204 60106
rect 272232 59530 272292 60106
rect 273320 59530 273380 60106
rect 273592 59530 273652 60106
rect 274408 59530 274468 60106
rect 275768 59530 275828 60106
rect 271144 59470 271338 59530
rect 270910 57901 270970 59470
rect 271278 57901 271338 59470
rect 272198 59470 272292 59530
rect 273302 59470 273380 59530
rect 273486 59470 273652 59530
rect 274406 59470 274468 59530
rect 275694 59470 275828 59530
rect 276040 59530 276100 60106
rect 276992 59530 277052 60106
rect 276040 59470 276122 59530
rect 272198 58173 272258 59470
rect 272195 58172 272261 58173
rect 272195 58108 272196 58172
rect 272260 58108 272261 58172
rect 272195 58107 272261 58108
rect 270907 57900 270973 57901
rect 270907 57836 270908 57900
rect 270972 57836 270973 57900
rect 270907 57835 270973 57836
rect 271275 57900 271341 57901
rect 271275 57836 271276 57900
rect 271340 57836 271341 57900
rect 271275 57835 271341 57836
rect 267595 57764 267661 57765
rect 267595 57700 267596 57764
rect 267660 57700 267661 57764
rect 267595 57699 267661 57700
rect 268331 57764 268397 57765
rect 268331 57700 268332 57764
rect 268396 57700 268397 57764
rect 268331 57699 268397 57700
rect 268699 57764 268765 57765
rect 268699 57700 268700 57764
rect 268764 57700 268765 57764
rect 268699 57699 268765 57700
rect 269803 57764 269869 57765
rect 269803 57700 269804 57764
rect 269868 57700 269869 57764
rect 269803 57699 269869 57700
rect 271794 57454 272414 58000
rect 273302 57901 273362 59470
rect 273299 57900 273365 57901
rect 273299 57836 273300 57900
rect 273364 57836 273365 57900
rect 273299 57835 273365 57836
rect 273486 57493 273546 59470
rect 274406 57765 274466 59470
rect 275694 58173 275754 59470
rect 276062 58853 276122 59470
rect 276982 59470 277052 59530
rect 278080 59530 278140 60106
rect 278488 59530 278548 60106
rect 279168 59530 279228 60106
rect 280936 59530 280996 60106
rect 283520 59530 283580 60106
rect 278080 59470 278146 59530
rect 276059 58852 276125 58853
rect 276059 58788 276060 58852
rect 276124 58788 276125 58852
rect 276059 58787 276125 58788
rect 275691 58172 275757 58173
rect 275691 58108 275692 58172
rect 275756 58108 275757 58172
rect 275691 58107 275757 58108
rect 274403 57764 274469 57765
rect 274403 57700 274404 57764
rect 274468 57700 274469 57764
rect 274403 57699 274469 57700
rect 266307 57356 266373 57357
rect 266307 57292 266308 57356
rect 266372 57292 266373 57356
rect 266307 57291 266373 57292
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 273483 57492 273549 57493
rect 273483 57428 273484 57492
rect 273548 57428 273549 57492
rect 273483 57427 273549 57428
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 25174 276134 58000
rect 276982 57765 277042 59470
rect 278086 57901 278146 59470
rect 278454 59470 278548 59530
rect 279006 59470 279228 59530
rect 280846 59470 280996 59530
rect 283422 59470 283580 59530
rect 285968 59530 286028 60106
rect 288280 59530 288340 60106
rect 291000 59530 291060 60106
rect 293448 59530 293508 60106
rect 285968 59470 286058 59530
rect 278454 58989 278514 59470
rect 278451 58988 278517 58989
rect 278451 58924 278452 58988
rect 278516 58924 278517 58988
rect 278451 58923 278517 58924
rect 279006 57901 279066 59470
rect 278083 57900 278149 57901
rect 278083 57836 278084 57900
rect 278148 57836 278149 57900
rect 278083 57835 278149 57836
rect 279003 57900 279069 57901
rect 279003 57836 279004 57900
rect 279068 57836 279069 57900
rect 279003 57835 279069 57836
rect 276979 57764 277045 57765
rect 276979 57700 276980 57764
rect 277044 57700 277045 57764
rect 276979 57699 277045 57700
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 28894 279854 58000
rect 280846 57629 280906 59470
rect 283422 59125 283482 59470
rect 283419 59124 283485 59125
rect 283419 59060 283420 59124
rect 283484 59060 283485 59124
rect 283419 59059 283485 59060
rect 280843 57628 280909 57629
rect 280843 57564 280844 57628
rect 280908 57564 280909 57628
rect 280843 57563 280909 57564
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 32614 283574 58000
rect 285998 56677 286058 59470
rect 288206 59470 288340 59530
rect 290966 59470 291060 59530
rect 293358 59470 293508 59530
rect 295896 59530 295956 60106
rect 298480 59530 298540 60106
rect 300928 59530 300988 60106
rect 303512 59530 303572 60106
rect 305960 59530 306020 60106
rect 308544 59669 308604 60106
rect 308541 59668 308607 59669
rect 308541 59604 308542 59668
rect 308606 59604 308607 59668
rect 308541 59603 308607 59604
rect 295896 59470 295994 59530
rect 298480 59470 298570 59530
rect 288206 57901 288266 59470
rect 290966 59261 291026 59470
rect 290963 59260 291029 59261
rect 290963 59196 290964 59260
rect 291028 59196 291029 59260
rect 290963 59195 291029 59196
rect 288203 57900 288269 57901
rect 288203 57836 288204 57900
rect 288268 57836 288269 57900
rect 288203 57835 288269 57836
rect 285995 56676 286061 56677
rect 285995 56612 285996 56676
rect 286060 56612 286061 56676
rect 285995 56611 286061 56612
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 39454 290414 58000
rect 293358 57901 293418 59470
rect 295934 59261 295994 59470
rect 298510 59261 298570 59470
rect 300902 59470 300988 59530
rect 303478 59470 303572 59530
rect 305870 59470 306020 59530
rect 310992 59530 311052 60106
rect 313440 59530 313500 60106
rect 315888 59530 315948 60106
rect 318472 59530 318532 60106
rect 310992 59470 311082 59530
rect 295931 59260 295997 59261
rect 295931 59196 295932 59260
rect 295996 59196 295997 59260
rect 295931 59195 295997 59196
rect 298507 59260 298573 59261
rect 298507 59196 298508 59260
rect 298572 59196 298573 59260
rect 298507 59195 298573 59196
rect 300902 58173 300962 59470
rect 303478 59261 303538 59470
rect 303475 59260 303541 59261
rect 303475 59196 303476 59260
rect 303540 59196 303541 59260
rect 303475 59195 303541 59196
rect 300899 58172 300965 58173
rect 300899 58108 300900 58172
rect 300964 58108 300965 58172
rect 300899 58107 300965 58108
rect 293355 57900 293421 57901
rect 293355 57836 293356 57900
rect 293420 57836 293421 57900
rect 293355 57835 293421 57836
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 43174 294134 58000
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 46894 297854 58000
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 50614 301574 58000
rect 305870 57901 305930 59470
rect 305867 57900 305933 57901
rect 305867 57836 305868 57900
rect 305932 57836 305933 57900
rect 305867 57835 305933 57836
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 57454 308414 58000
rect 311022 57901 311082 59470
rect 313414 59470 313500 59530
rect 315806 59470 315948 59530
rect 318382 59470 318532 59530
rect 320920 59530 320980 60106
rect 323368 59530 323428 60106
rect 325952 59530 326012 60106
rect 343224 59530 343284 60106
rect 320920 59470 321018 59530
rect 311019 57900 311085 57901
rect 311019 57836 311020 57900
rect 311084 57836 311085 57900
rect 311019 57835 311085 57836
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 25174 312134 58000
rect 313414 57901 313474 59470
rect 315806 58173 315866 59470
rect 315803 58172 315869 58173
rect 315803 58108 315804 58172
rect 315868 58108 315869 58172
rect 315803 58107 315869 58108
rect 313411 57900 313477 57901
rect 313411 57836 313412 57900
rect 313476 57836 313477 57900
rect 313411 57835 313477 57836
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 28894 315854 58000
rect 318382 57901 318442 59470
rect 318379 57900 318445 57901
rect 318379 57836 318380 57900
rect 318444 57836 318445 57900
rect 318379 57835 318445 57836
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 32614 319574 58000
rect 320958 56677 321018 59470
rect 323350 59470 323428 59530
rect 325926 59470 326012 59530
rect 343222 59470 343284 59530
rect 343360 59530 343420 60106
rect 343360 59470 343466 59530
rect 323350 56677 323410 59470
rect 325926 58173 325986 59470
rect 325923 58172 325989 58173
rect 325923 58108 325924 58172
rect 325988 58108 325989 58172
rect 325923 58107 325989 58108
rect 320955 56676 321021 56677
rect 320955 56612 320956 56676
rect 321020 56612 321021 56676
rect 320955 56611 321021 56612
rect 323347 56676 323413 56677
rect 323347 56612 323348 56676
rect 323412 56612 323413 56676
rect 323347 56611 323413 56612
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 39454 326414 58000
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 43174 330134 58000
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 46894 333854 58000
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 50614 337574 58000
rect 343222 57901 343282 59470
rect 343406 57901 343466 59470
rect 357942 59261 358002 491131
rect 358123 487796 358189 487797
rect 358123 487732 358124 487796
rect 358188 487732 358189 487796
rect 358123 487731 358189 487732
rect 357939 59260 358005 59261
rect 357939 59196 357940 59260
rect 358004 59196 358005 59260
rect 357939 59195 358005 59196
rect 343219 57900 343285 57901
rect 343219 57836 343220 57900
rect 343284 57836 343285 57900
rect 343219 57835 343285 57836
rect 343403 57900 343469 57901
rect 343403 57836 343404 57900
rect 343468 57836 343469 57900
rect 343403 57835 343469 57836
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 57454 344414 58000
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 25174 348134 58000
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 28894 351854 58000
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 32614 355574 58000
rect 358126 56677 358186 487731
rect 360699 483716 360765 483717
rect 360699 483652 360700 483716
rect 360764 483652 360765 483716
rect 360699 483651 360765 483652
rect 359411 478140 359477 478141
rect 359411 478076 359412 478140
rect 359476 478076 359477 478140
rect 359411 478075 359477 478076
rect 359414 272917 359474 478075
rect 360147 476780 360213 476781
rect 360147 476716 360148 476780
rect 360212 476716 360213 476780
rect 360147 476715 360213 476716
rect 359595 471476 359661 471477
rect 359595 471412 359596 471476
rect 359660 471412 359661 471476
rect 359595 471411 359661 471412
rect 359598 380221 359658 471411
rect 359779 468484 359845 468485
rect 359779 468420 359780 468484
rect 359844 468420 359845 468484
rect 359779 468419 359845 468420
rect 359595 380220 359661 380221
rect 359595 380156 359596 380220
rect 359660 380156 359661 380220
rect 359595 380155 359661 380156
rect 359782 378045 359842 468419
rect 359963 410548 360029 410549
rect 359963 410484 359964 410548
rect 360028 410484 360029 410548
rect 359963 410483 360029 410484
rect 359779 378044 359845 378045
rect 359779 377980 359780 378044
rect 359844 377980 359845 378044
rect 359779 377979 359845 377980
rect 359966 376005 360026 410483
rect 360150 379541 360210 476715
rect 360147 379540 360213 379541
rect 360147 379476 360148 379540
rect 360212 379476 360213 379540
rect 360147 379475 360213 379476
rect 359963 376004 360029 376005
rect 359963 375940 359964 376004
rect 360028 375940 360029 376004
rect 359963 375939 360029 375940
rect 359411 272916 359477 272917
rect 359411 272852 359412 272916
rect 359476 272852 359477 272916
rect 359411 272851 359477 272852
rect 360702 57493 360762 483651
rect 361794 471454 362414 506898
rect 365514 511174 366134 532000
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 363459 496092 363525 496093
rect 363459 496028 363460 496092
rect 363524 496028 363525 496092
rect 363459 496027 363525 496028
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 360699 57492 360765 57493
rect 360699 57428 360700 57492
rect 360764 57428 360765 57492
rect 360699 57427 360765 57428
rect 358123 56676 358189 56677
rect 358123 56612 358124 56676
rect 358188 56612 358189 56676
rect 358123 56611 358189 56612
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 363462 3501 363522 496027
rect 364931 493372 364997 493373
rect 364931 493308 364932 493372
rect 364996 493308 364997 493372
rect 364931 493307 364997 493308
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 363459 3500 363525 3501
rect 363459 3436 363460 3500
rect 363524 3436 363525 3500
rect 363459 3435 363525 3436
rect 364934 3365 364994 493307
rect 365514 475174 366134 510618
rect 369234 514894 369854 532000
rect 370635 529140 370701 529141
rect 370635 529076 370636 529140
rect 370700 529076 370701 529140
rect 370635 529075 370701 529076
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 367875 490924 367941 490925
rect 367875 490860 367876 490924
rect 367940 490860 367941 490924
rect 367875 490859 367941 490860
rect 367691 490788 367757 490789
rect 367691 490724 367692 490788
rect 367756 490724 367757 490788
rect 367691 490723 367757 490724
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 367694 58581 367754 490723
rect 367878 58853 367938 490859
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 370451 474060 370517 474061
rect 370451 473996 370452 474060
rect 370516 473996 370517 474060
rect 370451 473995 370517 473996
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 367875 58852 367941 58853
rect 367875 58788 367876 58852
rect 367940 58788 367941 58852
rect 367875 58787 367941 58788
rect 367691 58580 367757 58581
rect 367691 58516 367692 58580
rect 367756 58516 367757 58580
rect 367691 58515 367757 58516
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 364931 3364 364997 3365
rect 364931 3300 364932 3364
rect 364996 3300 364997 3364
rect 364931 3299 364997 3300
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 46894 369854 82338
rect 370454 57629 370514 473995
rect 370638 149157 370698 529075
rect 371739 526420 371805 526421
rect 371739 526356 371740 526420
rect 371804 526356 371805 526420
rect 371739 526355 371805 526356
rect 370635 149156 370701 149157
rect 370635 149092 370636 149156
rect 370700 149092 370701 149156
rect 370635 149091 370701 149092
rect 370451 57628 370517 57629
rect 370451 57564 370452 57628
rect 370516 57564 370517 57628
rect 370451 57563 370517 57564
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 371742 3637 371802 526355
rect 372954 518614 373574 532000
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 371923 491060 371989 491061
rect 371923 490996 371924 491060
rect 371988 490996 371989 491060
rect 371923 490995 371989 490996
rect 371926 59125 371986 490995
rect 372954 482614 373574 518058
rect 379794 525454 380414 532000
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 374499 490652 374565 490653
rect 374499 490588 374500 490652
rect 374564 490588 374565 490652
rect 374499 490587 374565 490588
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372659 482356 372725 482357
rect 372659 482292 372660 482356
rect 372724 482292 372725 482356
rect 372659 482291 372725 482292
rect 372954 482294 373574 482378
rect 372107 475420 372173 475421
rect 372107 475356 372108 475420
rect 372172 475356 372173 475420
rect 372107 475355 372173 475356
rect 371923 59124 371989 59125
rect 371923 59060 371924 59124
rect 371988 59060 371989 59124
rect 371923 59059 371989 59060
rect 372110 57765 372170 475355
rect 372662 377909 372722 482291
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372659 377908 372725 377909
rect 372659 377844 372660 377908
rect 372724 377844 372725 377908
rect 372659 377843 372725 377844
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372107 57764 372173 57765
rect 372107 57700 372108 57764
rect 372172 57700 372173 57764
rect 372107 57699 372173 57700
rect 372954 50614 373574 86058
rect 374502 58989 374562 490587
rect 375971 490516 376037 490517
rect 375971 490452 375972 490516
rect 376036 490452 376037 490516
rect 375971 490451 376037 490452
rect 374499 58988 374565 58989
rect 374499 58924 374500 58988
rect 374564 58924 374565 58988
rect 374499 58923 374565 58924
rect 375974 58717 376034 490451
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 378915 489156 378981 489157
rect 378915 489092 378916 489156
rect 378980 489092 378981 489156
rect 378915 489091 378981 489092
rect 379794 489134 380414 489218
rect 378731 486436 378797 486437
rect 378731 486372 378732 486436
rect 378796 486372 378797 486436
rect 378731 486371 378797 486372
rect 376155 485076 376221 485077
rect 376155 485012 376156 485076
rect 376220 485012 376221 485076
rect 376155 485011 376221 485012
rect 375971 58716 376037 58717
rect 375971 58652 375972 58716
rect 376036 58652 376037 58716
rect 375971 58651 376037 58652
rect 376158 57357 376218 485011
rect 376339 480996 376405 480997
rect 376339 480932 376340 480996
rect 376404 480932 376405 480996
rect 376339 480931 376405 480932
rect 376155 57356 376221 57357
rect 376155 57292 376156 57356
rect 376220 57292 376221 57356
rect 376155 57291 376221 57292
rect 376342 57085 376402 480931
rect 378179 479500 378245 479501
rect 378179 479436 378180 479500
rect 378244 479436 378245 479500
rect 378179 479435 378245 479436
rect 377259 475556 377325 475557
rect 377259 475492 377260 475556
rect 377324 475492 377325 475556
rect 377259 475491 377325 475492
rect 376707 375324 376773 375325
rect 376707 375260 376708 375324
rect 376772 375260 376773 375324
rect 376707 375259 376773 375260
rect 376710 369870 376770 375259
rect 376710 369810 376954 369870
rect 376894 273325 376954 369810
rect 376891 273324 376957 273325
rect 376891 273260 376892 273324
rect 376956 273260 376957 273324
rect 376891 273259 376957 273260
rect 377262 271421 377322 475491
rect 377443 471340 377509 471341
rect 377443 471276 377444 471340
rect 377508 471276 377509 471340
rect 377443 471275 377509 471276
rect 377446 378725 377506 471275
rect 377627 471204 377693 471205
rect 377627 471140 377628 471204
rect 377692 471140 377693 471204
rect 377627 471139 377693 471140
rect 377630 378861 377690 471139
rect 377811 465900 377877 465901
rect 377811 465836 377812 465900
rect 377876 465836 377877 465900
rect 377811 465835 377877 465836
rect 377627 378860 377693 378861
rect 377627 378796 377628 378860
rect 377692 378796 377693 378860
rect 377627 378795 377693 378796
rect 377443 378724 377509 378725
rect 377443 378660 377444 378724
rect 377508 378660 377509 378724
rect 377443 378659 377509 378660
rect 377814 375325 377874 465835
rect 377811 375324 377877 375325
rect 377811 375260 377812 375324
rect 377876 375260 377877 375324
rect 377811 375259 377877 375260
rect 377995 273324 378061 273325
rect 377995 273260 377996 273324
rect 378060 273260 378061 273324
rect 377995 273259 378061 273260
rect 377998 272781 378058 273259
rect 377995 272780 378061 272781
rect 377995 272716 377996 272780
rect 378060 272716 378061 272780
rect 377995 272715 378061 272716
rect 377259 271420 377325 271421
rect 377259 271356 377260 271420
rect 377324 271356 377325 271420
rect 377259 271355 377325 271356
rect 377995 251836 378061 251837
rect 377995 251772 377996 251836
rect 378060 251772 378061 251836
rect 377995 251771 378061 251772
rect 377259 163028 377325 163029
rect 377259 162964 377260 163028
rect 377324 162964 377325 163028
rect 377259 162963 377325 162964
rect 376339 57084 376405 57085
rect 376339 57020 376340 57084
rect 376404 57020 376405 57084
rect 376339 57019 376405 57020
rect 377262 56541 377322 162963
rect 377998 162621 378058 251771
rect 377995 162620 378061 162621
rect 377995 162556 377996 162620
rect 378060 162556 378061 162620
rect 377995 162555 378061 162556
rect 377811 144124 377877 144125
rect 377811 144060 377812 144124
rect 377876 144060 377877 144124
rect 377811 144059 377877 144060
rect 377259 56540 377325 56541
rect 377259 56476 377260 56540
rect 377324 56476 377325 56540
rect 377259 56475 377325 56476
rect 377814 55181 377874 144059
rect 377998 58445 378058 162555
rect 378182 60621 378242 479435
rect 378363 472564 378429 472565
rect 378363 472500 378364 472564
rect 378428 472500 378429 472564
rect 378363 472499 378429 472500
rect 378366 273325 378426 472499
rect 378363 273324 378429 273325
rect 378363 273260 378364 273324
rect 378428 273260 378429 273324
rect 378363 273259 378429 273260
rect 378179 60620 378245 60621
rect 378179 60556 378180 60620
rect 378244 60556 378245 60620
rect 378179 60555 378245 60556
rect 377995 58444 378061 58445
rect 377995 58380 377996 58444
rect 378060 58380 378061 58444
rect 377995 58379 378061 58380
rect 378734 57221 378794 486371
rect 378918 165205 378978 489091
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379467 481132 379533 481133
rect 379467 481068 379468 481132
rect 379532 481130 379533 481132
rect 379532 481070 379714 481130
rect 379532 481068 379533 481070
rect 379467 481067 379533 481068
rect 379654 277410 379714 481070
rect 379794 466308 380414 488898
rect 383514 529174 384134 532000
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 466308 384134 492618
rect 387234 496894 387854 532000
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 466308 387854 496338
rect 390954 500614 391574 532000
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 466308 391574 500058
rect 397794 507454 398414 532000
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 466308 398414 470898
rect 401514 511174 402134 532000
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 466308 402134 474618
rect 405234 514894 405854 532000
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 466308 405854 478338
rect 408954 518614 409574 532000
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 466308 409574 482058
rect 415794 525454 416414 532000
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 466308 416414 488898
rect 419514 529174 420134 532000
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 466308 420134 492618
rect 423234 496894 423854 532000
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 466308 423854 496338
rect 426954 500614 427574 532000
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 466308 427574 500058
rect 433794 507454 434414 532000
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 466308 434414 470898
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 466308 438134 474618
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 466308 441854 478338
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 466308 445574 482058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 466308 452414 488898
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 642000 459854 676338
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 642000 463574 644058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 642000 470414 650898
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 642000 474134 654618
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 642000 477854 658338
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 642000 481574 662058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 642000 488414 668898
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 642000 492134 672618
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 642000 495854 676338
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 642000 499574 644058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 642000 506414 650898
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 642000 510134 654618
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 476067 639980 476133 639981
rect 476067 639916 476068 639980
rect 476132 639916 476133 639980
rect 476067 639915 476133 639916
rect 488579 639980 488645 639981
rect 488579 639916 488580 639980
rect 488644 639916 488645 639980
rect 488579 639915 488645 639916
rect 506611 639980 506677 639981
rect 506611 639916 506612 639980
rect 506676 639916 506677 639980
rect 506611 639915 506677 639916
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 464208 615454 464528 615486
rect 464208 615218 464250 615454
rect 464486 615218 464528 615454
rect 464208 615134 464528 615218
rect 464208 614898 464250 615134
rect 464486 614898 464528 615134
rect 464208 614866 464528 614898
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 466308 456134 492618
rect 459234 568894 459854 588000
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 466308 459854 496338
rect 462954 572614 463574 588000
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 466308 463574 500058
rect 469794 579454 470414 588000
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 466308 470414 470898
rect 473514 583174 474134 588000
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 476070 496093 476130 639915
rect 479568 633454 479888 633486
rect 479568 633218 479610 633454
rect 479846 633218 479888 633454
rect 479568 633134 479888 633218
rect 479568 632898 479610 633134
rect 479846 632898 479888 633134
rect 479568 632866 479888 632898
rect 479568 597454 479888 597486
rect 479568 597218 479610 597454
rect 479846 597218 479888 597454
rect 479568 597134 479888 597218
rect 479568 596898 479610 597134
rect 479846 596898 479888 597134
rect 479568 596866 479888 596898
rect 477234 586894 477854 588000
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 476067 496092 476133 496093
rect 476067 496028 476068 496092
rect 476132 496028 476133 496092
rect 476067 496027 476133 496028
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 466308 474134 474618
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 466308 477854 478338
rect 480954 554614 481574 588000
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 466308 481574 482058
rect 487794 561454 488414 588000
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 488582 491877 488642 639915
rect 494928 615454 495248 615486
rect 494928 615218 494970 615454
rect 495206 615218 495248 615454
rect 494928 615134 495248 615218
rect 494928 614898 494970 615134
rect 495206 614898 495248 615134
rect 494928 614866 495248 614898
rect 491514 565174 492134 588000
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 488579 491876 488645 491877
rect 488579 491812 488580 491876
rect 488644 491812 488645 491876
rect 488579 491811 488645 491812
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 466308 488414 488898
rect 491514 466308 492134 492618
rect 495234 568894 495854 588000
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 466308 495854 496338
rect 498954 572614 499574 588000
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498515 466580 498581 466581
rect 498515 466516 498516 466580
rect 498580 466516 498581 466580
rect 498515 466515 498581 466516
rect 498518 464810 498578 466515
rect 498954 466308 499574 500058
rect 505794 579454 506414 588000
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 506614 472701 506674 639915
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 509514 583174 510134 588000
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 506611 472700 506677 472701
rect 506611 472636 506612 472700
rect 506676 472636 506677 472700
rect 506611 472635 506677 472636
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 499803 466580 499869 466581
rect 499803 466516 499804 466580
rect 499868 466516 499869 466580
rect 499803 466515 499869 466516
rect 499806 464810 499866 466515
rect 505794 466308 506414 470898
rect 509514 466308 510134 474618
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 510843 466580 510909 466581
rect 510843 466516 510844 466580
rect 510908 466516 510909 466580
rect 510843 466515 510909 466516
rect 510846 464810 510906 466515
rect 513234 466308 513854 478338
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 466308 517574 482058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 498464 464750 498578 464810
rect 499688 464750 499866 464810
rect 510840 464750 510906 464810
rect 498464 464202 498524 464750
rect 499688 464202 499748 464750
rect 510840 464202 510900 464750
rect 380272 453454 380620 453486
rect 380272 453218 380328 453454
rect 380564 453218 380620 453454
rect 380272 453134 380620 453218
rect 380272 452898 380328 453134
rect 380564 452898 380620 453134
rect 380272 452866 380620 452898
rect 516000 453454 516348 453486
rect 516000 453218 516056 453454
rect 516292 453218 516348 453454
rect 516000 453134 516348 453218
rect 516000 452898 516056 453134
rect 516292 452898 516348 453134
rect 516000 452866 516348 452898
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 380952 435454 381300 435486
rect 380952 435218 381008 435454
rect 381244 435218 381300 435454
rect 380952 435134 381300 435218
rect 380952 434898 381008 435134
rect 381244 434898 381300 435134
rect 380952 434866 381300 434898
rect 515320 435454 515668 435486
rect 515320 435218 515376 435454
rect 515612 435218 515668 435454
rect 515320 435134 515668 435218
rect 515320 434898 515376 435134
rect 515612 434898 515668 435134
rect 515320 434866 515668 434898
rect 380272 417454 380620 417486
rect 380272 417218 380328 417454
rect 380564 417218 380620 417454
rect 380272 417134 380620 417218
rect 380272 416898 380328 417134
rect 380564 416898 380620 417134
rect 380272 416866 380620 416898
rect 516000 417454 516348 417486
rect 516000 417218 516056 417454
rect 516292 417218 516348 417454
rect 516000 417134 516348 417218
rect 516000 416898 516056 417134
rect 516292 416898 516348 417134
rect 516000 416866 516348 416898
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 380952 399454 381300 399486
rect 380952 399218 381008 399454
rect 381244 399218 381300 399454
rect 380952 399134 381300 399218
rect 380952 398898 381008 399134
rect 381244 398898 381300 399134
rect 380952 398866 381300 398898
rect 515320 399454 515668 399486
rect 515320 399218 515376 399454
rect 515612 399218 515668 399454
rect 515320 399134 515668 399218
rect 515320 398898 515376 399134
rect 515612 398898 515668 399134
rect 515320 398866 515668 398898
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 396056 380490 396116 381106
rect 397144 380490 397204 381106
rect 396030 380430 396116 380490
rect 397134 380430 397204 380490
rect 398232 380490 398292 381106
rect 399592 380490 399652 381106
rect 400544 380490 400604 381106
rect 401768 380490 401828 381106
rect 403128 380490 403188 381106
rect 404216 380629 404276 381106
rect 405440 380629 405500 381106
rect 404213 380628 404279 380629
rect 404213 380564 404214 380628
rect 404278 380564 404279 380628
rect 404213 380563 404279 380564
rect 405437 380628 405503 380629
rect 405437 380564 405438 380628
rect 405502 380564 405503 380628
rect 405437 380563 405503 380564
rect 406528 380490 406588 381106
rect 398232 380430 398298 380490
rect 396030 379405 396090 380430
rect 397134 379405 397194 380430
rect 398238 379405 398298 380430
rect 399526 380430 399652 380490
rect 400446 380430 400604 380490
rect 401734 380430 401828 380490
rect 403022 380430 403188 380490
rect 406518 380430 406588 380490
rect 407616 380490 407676 381106
rect 408296 380490 408356 381106
rect 408704 380490 408764 381106
rect 410064 380490 410124 381106
rect 407616 380430 407682 380490
rect 408296 380430 408418 380490
rect 408704 380430 408786 380490
rect 399526 379405 399586 380430
rect 396027 379404 396093 379405
rect 396027 379340 396028 379404
rect 396092 379340 396093 379404
rect 396027 379339 396093 379340
rect 397131 379404 397197 379405
rect 397131 379340 397132 379404
rect 397196 379340 397197 379404
rect 397131 379339 397197 379340
rect 398235 379404 398301 379405
rect 398235 379340 398236 379404
rect 398300 379340 398301 379404
rect 398235 379339 398301 379340
rect 399523 379404 399589 379405
rect 399523 379340 399524 379404
rect 399588 379340 399589 379404
rect 399523 379339 399589 379340
rect 400446 379133 400506 380430
rect 401734 379269 401794 380430
rect 403022 379269 403082 380430
rect 406518 379405 406578 380430
rect 407622 379405 407682 380430
rect 408358 379405 408418 380430
rect 406515 379404 406581 379405
rect 406515 379340 406516 379404
rect 406580 379340 406581 379404
rect 406515 379339 406581 379340
rect 407619 379404 407685 379405
rect 407619 379340 407620 379404
rect 407684 379340 407685 379404
rect 407619 379339 407685 379340
rect 408355 379404 408421 379405
rect 408355 379340 408356 379404
rect 408420 379340 408421 379404
rect 408355 379339 408421 379340
rect 401731 379268 401797 379269
rect 401731 379204 401732 379268
rect 401796 379204 401797 379268
rect 401731 379203 401797 379204
rect 403019 379268 403085 379269
rect 403019 379204 403020 379268
rect 403084 379204 403085 379268
rect 403019 379203 403085 379204
rect 400443 379132 400509 379133
rect 400443 379068 400444 379132
rect 400508 379068 400509 379132
rect 400443 379067 400509 379068
rect 379794 364394 380414 379000
rect 379794 364158 379826 364394
rect 380062 364158 380146 364394
rect 380382 364158 380414 364394
rect 379794 364074 380414 364158
rect 379794 363838 379826 364074
rect 380062 363838 380146 364074
rect 380382 363838 380414 364074
rect 379794 359308 380414 363838
rect 383514 368114 384134 379000
rect 383514 367878 383546 368114
rect 383782 367878 383866 368114
rect 384102 367878 384134 368114
rect 383514 367794 384134 367878
rect 383514 367558 383546 367794
rect 383782 367558 383866 367794
rect 384102 367558 384134 367794
rect 383514 359308 384134 367558
rect 387234 369954 387854 379000
rect 387234 369718 387266 369954
rect 387502 369718 387586 369954
rect 387822 369718 387854 369954
rect 387234 369634 387854 369718
rect 387234 369398 387266 369634
rect 387502 369398 387586 369634
rect 387822 369398 387854 369634
rect 387234 359308 387854 369398
rect 390954 373674 391574 379000
rect 390954 373438 390986 373674
rect 391222 373438 391306 373674
rect 391542 373438 391574 373674
rect 390954 373354 391574 373438
rect 390954 373118 390986 373354
rect 391222 373118 391306 373354
rect 391542 373118 391574 373354
rect 390954 359308 391574 373118
rect 397794 363454 398414 379000
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 359308 398414 362898
rect 401514 367174 402134 379000
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 359308 402134 366618
rect 405234 370894 405854 379000
rect 408726 378589 408786 380430
rect 410014 380430 410124 380490
rect 410744 380490 410804 381106
rect 411288 380490 411348 381106
rect 412376 380490 412436 381106
rect 413464 380629 413524 381106
rect 413600 380901 413660 381106
rect 413597 380900 413663 380901
rect 413597 380836 413598 380900
rect 413662 380836 413663 380900
rect 413597 380835 413663 380836
rect 413461 380628 413527 380629
rect 413461 380564 413462 380628
rect 413526 380564 413527 380628
rect 413461 380563 413527 380564
rect 414552 380490 414612 381106
rect 415912 380490 415972 381106
rect 410744 380430 410810 380490
rect 411288 380430 411362 380490
rect 412376 380430 412466 380490
rect 414552 380430 414674 380490
rect 408723 378588 408789 378589
rect 408723 378524 408724 378588
rect 408788 378524 408789 378588
rect 408723 378523 408789 378524
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 359308 405854 370338
rect 408954 374614 409574 379000
rect 410014 378181 410074 380430
rect 410750 379405 410810 380430
rect 411302 379405 411362 380430
rect 412406 379405 412466 380430
rect 410747 379404 410813 379405
rect 410747 379340 410748 379404
rect 410812 379340 410813 379404
rect 410747 379339 410813 379340
rect 411299 379404 411365 379405
rect 411299 379340 411300 379404
rect 411364 379340 411365 379404
rect 411299 379339 411365 379340
rect 412403 379404 412469 379405
rect 412403 379340 412404 379404
rect 412468 379340 412469 379404
rect 412403 379339 412469 379340
rect 414614 379269 414674 380430
rect 415902 380430 415972 380490
rect 416048 380490 416108 381106
rect 417000 380490 417060 381106
rect 418088 380490 418148 381106
rect 418496 380490 418556 381106
rect 419448 380490 419508 381106
rect 416048 380430 416146 380490
rect 417000 380430 417066 380490
rect 418088 380430 418170 380490
rect 415902 379269 415962 380430
rect 416086 379269 416146 380430
rect 414611 379268 414677 379269
rect 414611 379204 414612 379268
rect 414676 379204 414677 379268
rect 414611 379203 414677 379204
rect 415899 379268 415965 379269
rect 415899 379204 415900 379268
rect 415964 379204 415965 379268
rect 415899 379203 415965 379204
rect 416083 379268 416149 379269
rect 416083 379204 416084 379268
rect 416148 379204 416149 379268
rect 416083 379203 416149 379204
rect 410011 378180 410077 378181
rect 410011 378116 410012 378180
rect 410076 378116 410077 378180
rect 410011 378115 410077 378116
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 359308 409574 374058
rect 415794 364394 416414 379000
rect 417006 378181 417066 380430
rect 418110 378181 418170 380430
rect 418478 380430 418556 380490
rect 419398 380430 419508 380490
rect 420672 380490 420732 381106
rect 421080 380901 421140 381106
rect 421077 380900 421143 380901
rect 421077 380836 421078 380900
rect 421142 380836 421143 380900
rect 421077 380835 421143 380836
rect 421760 380490 421820 381106
rect 422848 380490 422908 381106
rect 423528 380490 423588 381106
rect 420672 380430 420746 380490
rect 421760 380430 421850 380490
rect 422848 380430 422954 380490
rect 418478 378589 418538 380430
rect 419398 379133 419458 380430
rect 420686 379405 420746 380430
rect 420683 379404 420749 379405
rect 420683 379340 420684 379404
rect 420748 379340 420749 379404
rect 420683 379339 420749 379340
rect 419395 379132 419461 379133
rect 419395 379068 419396 379132
rect 419460 379068 419461 379132
rect 419395 379067 419461 379068
rect 418475 378588 418541 378589
rect 418475 378524 418476 378588
rect 418540 378524 418541 378588
rect 418475 378523 418541 378524
rect 417003 378180 417069 378181
rect 417003 378116 417004 378180
rect 417068 378116 417069 378180
rect 417003 378115 417069 378116
rect 418107 378180 418173 378181
rect 418107 378116 418108 378180
rect 418172 378116 418173 378180
rect 418107 378115 418173 378116
rect 415794 364158 415826 364394
rect 416062 364158 416146 364394
rect 416382 364158 416414 364394
rect 415794 364074 416414 364158
rect 415794 363838 415826 364074
rect 416062 363838 416146 364074
rect 416382 363838 416414 364074
rect 415794 359308 416414 363838
rect 419514 368114 420134 379000
rect 421790 378589 421850 380430
rect 421787 378588 421853 378589
rect 421787 378524 421788 378588
rect 421852 378524 421853 378588
rect 421787 378523 421853 378524
rect 422894 378317 422954 380430
rect 423446 380430 423588 380490
rect 423936 380490 423996 381106
rect 425296 380490 425356 381106
rect 425976 380901 426036 381106
rect 425973 380900 426039 380901
rect 425973 380836 425974 380900
rect 426038 380836 426039 380900
rect 425973 380835 426039 380836
rect 423936 380430 424058 380490
rect 423446 379269 423506 380430
rect 423443 379268 423509 379269
rect 423443 379204 423444 379268
rect 423508 379204 423509 379268
rect 423443 379203 423509 379204
rect 422891 378316 422957 378317
rect 422891 378252 422892 378316
rect 422956 378252 422957 378316
rect 422891 378251 422957 378252
rect 419514 367878 419546 368114
rect 419782 367878 419866 368114
rect 420102 367878 420134 368114
rect 419514 367794 420134 367878
rect 419514 367558 419546 367794
rect 419782 367558 419866 367794
rect 420102 367558 420134 367794
rect 419514 359308 420134 367558
rect 423234 369954 423854 379000
rect 423998 378181 424058 380430
rect 425286 380430 425356 380490
rect 426384 380490 426444 381106
rect 427608 380490 427668 381106
rect 428288 380490 428348 381106
rect 428696 380490 428756 381106
rect 429784 380490 429844 381106
rect 431008 380490 431068 381106
rect 426384 380430 426450 380490
rect 425286 378181 425346 380430
rect 426390 378181 426450 380430
rect 427494 380430 427668 380490
rect 428230 380430 428348 380490
rect 428598 380430 428756 380490
rect 429702 380430 429844 380490
rect 430990 380430 431068 380490
rect 431144 380490 431204 381106
rect 432232 380490 432292 381106
rect 433320 380490 433380 381106
rect 433592 380901 433652 381106
rect 433589 380900 433655 380901
rect 433589 380836 433590 380900
rect 433654 380836 433655 380900
rect 433589 380835 433655 380836
rect 434408 380490 434468 381106
rect 431144 380430 431234 380490
rect 432232 380430 432338 380490
rect 433320 380430 433442 380490
rect 427494 380221 427554 380430
rect 427491 380220 427557 380221
rect 427491 380156 427492 380220
rect 427556 380156 427557 380220
rect 427491 380155 427557 380156
rect 428230 379405 428290 380430
rect 428227 379404 428293 379405
rect 428227 379340 428228 379404
rect 428292 379340 428293 379404
rect 428227 379339 428293 379340
rect 423995 378180 424061 378181
rect 423995 378116 423996 378180
rect 424060 378116 424061 378180
rect 423995 378115 424061 378116
rect 425283 378180 425349 378181
rect 425283 378116 425284 378180
rect 425348 378116 425349 378180
rect 425283 378115 425349 378116
rect 426387 378180 426453 378181
rect 426387 378116 426388 378180
rect 426452 378116 426453 378180
rect 426387 378115 426453 378116
rect 423234 369718 423266 369954
rect 423502 369718 423586 369954
rect 423822 369718 423854 369954
rect 423234 369634 423854 369718
rect 423234 369398 423266 369634
rect 423502 369398 423586 369634
rect 423822 369398 423854 369634
rect 423234 359308 423854 369398
rect 426954 373674 427574 379000
rect 428598 378181 428658 380430
rect 429702 378861 429762 380430
rect 429699 378860 429765 378861
rect 429699 378796 429700 378860
rect 429764 378796 429765 378860
rect 429699 378795 429765 378796
rect 430990 378589 431050 380430
rect 431174 379405 431234 380430
rect 431171 379404 431237 379405
rect 431171 379340 431172 379404
rect 431236 379340 431237 379404
rect 431171 379339 431237 379340
rect 430987 378588 431053 378589
rect 430987 378524 430988 378588
rect 431052 378524 431053 378588
rect 430987 378523 431053 378524
rect 432278 378181 432338 380430
rect 433382 378725 433442 380430
rect 434302 380430 434468 380490
rect 435768 380490 435828 381106
rect 436040 380901 436100 381106
rect 436037 380900 436103 380901
rect 436037 380836 436038 380900
rect 436102 380836 436103 380900
rect 436037 380835 436103 380836
rect 436992 380490 437052 381106
rect 438080 380490 438140 381106
rect 438488 380765 438548 381106
rect 438485 380764 438551 380765
rect 438485 380700 438486 380764
rect 438550 380700 438551 380764
rect 438485 380699 438551 380700
rect 439168 380490 439228 381106
rect 440936 380765 440996 381106
rect 443520 380765 443580 381106
rect 440933 380764 440999 380765
rect 440933 380700 440934 380764
rect 440998 380700 440999 380764
rect 440933 380699 440999 380700
rect 443517 380764 443583 380765
rect 443517 380700 443518 380764
rect 443582 380700 443583 380764
rect 443517 380699 443583 380700
rect 445968 380629 446028 381106
rect 448280 380765 448340 381106
rect 448277 380764 448343 380765
rect 448277 380700 448278 380764
rect 448342 380700 448343 380764
rect 448277 380699 448343 380700
rect 445965 380628 446031 380629
rect 445965 380564 445966 380628
rect 446030 380564 446031 380628
rect 445965 380563 446031 380564
rect 435768 380430 435834 380490
rect 434302 379405 434362 380430
rect 434299 379404 434365 379405
rect 434299 379340 434300 379404
rect 434364 379340 434365 379404
rect 434299 379339 434365 379340
rect 433379 378724 433445 378725
rect 433379 378660 433380 378724
rect 433444 378660 433445 378724
rect 433379 378659 433445 378660
rect 428595 378180 428661 378181
rect 428595 378116 428596 378180
rect 428660 378116 428661 378180
rect 428595 378115 428661 378116
rect 432275 378180 432341 378181
rect 432275 378116 432276 378180
rect 432340 378116 432341 378180
rect 432275 378115 432341 378116
rect 426954 373438 426986 373674
rect 427222 373438 427306 373674
rect 427542 373438 427574 373674
rect 426954 373354 427574 373438
rect 426954 373118 426986 373354
rect 427222 373118 427306 373354
rect 427542 373118 427574 373354
rect 426954 359308 427574 373118
rect 433794 363454 434414 379000
rect 435774 378181 435834 380430
rect 436878 380430 437052 380490
rect 437982 380430 438140 380490
rect 439086 380430 439228 380490
rect 451000 380490 451060 381106
rect 453448 380490 453508 381106
rect 455896 380490 455956 381106
rect 458480 380490 458540 381106
rect 451000 380430 451106 380490
rect 436878 378589 436938 380430
rect 437982 379405 438042 380430
rect 437979 379404 438045 379405
rect 437979 379340 437980 379404
rect 438044 379340 438045 379404
rect 437979 379339 438045 379340
rect 436875 378588 436941 378589
rect 436875 378524 436876 378588
rect 436940 378524 436941 378588
rect 436875 378523 436941 378524
rect 435771 378180 435837 378181
rect 435771 378116 435772 378180
rect 435836 378116 435837 378180
rect 435771 378115 435837 378116
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 359308 434414 362898
rect 437514 367174 438134 379000
rect 439086 378181 439146 380430
rect 451046 379405 451106 380430
rect 453438 380430 453508 380490
rect 455830 380430 455956 380490
rect 458406 380430 458540 380490
rect 460928 380490 460988 381106
rect 463512 380490 463572 381106
rect 465960 380490 466020 381106
rect 468544 380490 468604 381106
rect 470992 380490 471052 381106
rect 460928 380430 461042 380490
rect 463512 380430 463618 380490
rect 453438 379405 453498 380430
rect 455830 379405 455890 380430
rect 451043 379404 451109 379405
rect 451043 379340 451044 379404
rect 451108 379340 451109 379404
rect 451043 379339 451109 379340
rect 453435 379404 453501 379405
rect 453435 379340 453436 379404
rect 453500 379340 453501 379404
rect 453435 379339 453501 379340
rect 455827 379404 455893 379405
rect 455827 379340 455828 379404
rect 455892 379340 455893 379404
rect 455827 379339 455893 379340
rect 439083 378180 439149 378181
rect 439083 378116 439084 378180
rect 439148 378116 439149 378180
rect 439083 378115 439149 378116
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 359308 438134 366618
rect 441234 370894 441854 379000
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 359308 441854 370338
rect 444954 374614 445574 379000
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 359308 445574 374058
rect 451794 364394 452414 379000
rect 451794 364158 451826 364394
rect 452062 364158 452146 364394
rect 452382 364158 452414 364394
rect 451794 364074 452414 364158
rect 451794 363838 451826 364074
rect 452062 363838 452146 364074
rect 452382 363838 452414 364074
rect 451794 359308 452414 363838
rect 455514 368114 456134 379000
rect 458406 378181 458466 380430
rect 460982 379405 461042 380430
rect 463558 379405 463618 380430
rect 465950 380430 466020 380490
rect 468526 380430 468604 380490
rect 470918 380430 471052 380490
rect 473440 380490 473500 381106
rect 475888 380490 475948 381106
rect 478472 380490 478532 381106
rect 480920 380490 480980 381106
rect 473440 380430 473554 380490
rect 460979 379404 461045 379405
rect 460979 379340 460980 379404
rect 461044 379340 461045 379404
rect 460979 379339 461045 379340
rect 463555 379404 463621 379405
rect 463555 379340 463556 379404
rect 463620 379340 463621 379404
rect 463555 379339 463621 379340
rect 465950 379133 466010 380430
rect 465947 379132 466013 379133
rect 465947 379068 465948 379132
rect 466012 379068 466013 379132
rect 465947 379067 466013 379068
rect 458403 378180 458469 378181
rect 458403 378116 458404 378180
rect 458468 378116 458469 378180
rect 458403 378115 458469 378116
rect 455514 367878 455546 368114
rect 455782 367878 455866 368114
rect 456102 367878 456134 368114
rect 455514 367794 456134 367878
rect 455514 367558 455546 367794
rect 455782 367558 455866 367794
rect 456102 367558 456134 367794
rect 455514 359308 456134 367558
rect 459234 369954 459854 379000
rect 459234 369718 459266 369954
rect 459502 369718 459586 369954
rect 459822 369718 459854 369954
rect 459234 369634 459854 369718
rect 459234 369398 459266 369634
rect 459502 369398 459586 369634
rect 459822 369398 459854 369634
rect 459234 359308 459854 369398
rect 462954 373674 463574 379000
rect 468526 378861 468586 380430
rect 468523 378860 468589 378861
rect 468523 378796 468524 378860
rect 468588 378796 468589 378860
rect 468523 378795 468589 378796
rect 462954 373438 462986 373674
rect 463222 373438 463306 373674
rect 463542 373438 463574 373674
rect 462954 373354 463574 373438
rect 462954 373118 462986 373354
rect 463222 373118 463306 373354
rect 463542 373118 463574 373354
rect 462954 359308 463574 373118
rect 469794 363454 470414 379000
rect 470918 378997 470978 380430
rect 473494 379405 473554 380430
rect 475886 380430 475948 380490
rect 478462 380430 478532 380490
rect 480854 380430 480980 380490
rect 483368 380490 483428 381106
rect 485952 380490 486012 381106
rect 503224 380490 503284 381106
rect 503360 380629 503420 381106
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 503357 380628 503423 380629
rect 503357 380564 503358 380628
rect 503422 380564 503423 380628
rect 503357 380563 503423 380564
rect 483368 380430 483490 380490
rect 485952 380430 486066 380490
rect 503224 380430 503362 380490
rect 473491 379404 473557 379405
rect 473491 379340 473492 379404
rect 473556 379340 473557 379404
rect 473491 379339 473557 379340
rect 470915 378996 470981 378997
rect 470915 378932 470916 378996
rect 470980 378932 470981 378996
rect 470915 378931 470981 378932
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 359308 470414 362898
rect 473514 367174 474134 379000
rect 475886 378861 475946 380430
rect 475883 378860 475949 378861
rect 475883 378796 475884 378860
rect 475948 378796 475949 378860
rect 475883 378795 475949 378796
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 359308 474134 366618
rect 477234 370894 477854 379000
rect 478462 378861 478522 380430
rect 480854 379405 480914 380430
rect 480851 379404 480917 379405
rect 480851 379340 480852 379404
rect 480916 379340 480917 379404
rect 480851 379339 480917 379340
rect 478459 378860 478525 378861
rect 478459 378796 478460 378860
rect 478524 378796 478525 378860
rect 478459 378795 478525 378796
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 359308 477854 370338
rect 480954 374614 481574 379000
rect 483430 378861 483490 380430
rect 486006 379405 486066 380430
rect 503302 379405 503362 380430
rect 486003 379404 486069 379405
rect 486003 379340 486004 379404
rect 486068 379340 486069 379404
rect 486003 379339 486069 379340
rect 503299 379404 503365 379405
rect 503299 379340 503300 379404
rect 503364 379340 503365 379404
rect 503299 379339 503365 379340
rect 483427 378860 483493 378861
rect 483427 378796 483428 378860
rect 483492 378796 483493 378860
rect 483427 378795 483493 378796
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 359308 481574 374058
rect 487794 364394 488414 379000
rect 487794 364158 487826 364394
rect 488062 364158 488146 364394
rect 488382 364158 488414 364394
rect 487794 364074 488414 364158
rect 487794 363838 487826 364074
rect 488062 363838 488146 364074
rect 488382 363838 488414 364074
rect 487794 359308 488414 363838
rect 491514 368114 492134 379000
rect 491514 367878 491546 368114
rect 491782 367878 491866 368114
rect 492102 367878 492134 368114
rect 491514 367794 492134 367878
rect 491514 367558 491546 367794
rect 491782 367558 491866 367794
rect 492102 367558 492134 367794
rect 491514 359308 492134 367558
rect 495234 369954 495854 379000
rect 495234 369718 495266 369954
rect 495502 369718 495586 369954
rect 495822 369718 495854 369954
rect 495234 369634 495854 369718
rect 495234 369398 495266 369634
rect 495502 369398 495586 369634
rect 495822 369398 495854 369634
rect 495234 359308 495854 369398
rect 498954 373674 499574 379000
rect 498954 373438 498986 373674
rect 499222 373438 499306 373674
rect 499542 373438 499574 373674
rect 498954 373354 499574 373438
rect 498954 373118 498986 373354
rect 499222 373118 499306 373354
rect 499542 373118 499574 373354
rect 498954 359308 499574 373118
rect 505794 363454 506414 379000
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 359308 506414 362898
rect 509514 367174 510134 379000
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 359308 510134 366618
rect 513234 370894 513854 379000
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 359308 513854 370338
rect 516954 374614 517574 379000
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 359308 517574 374058
rect 498515 358868 498581 358869
rect 498515 358804 498516 358868
rect 498580 358804 498581 358868
rect 498515 358803 498581 358804
rect 499803 358868 499869 358869
rect 499803 358804 499804 358868
rect 499868 358804 499869 358868
rect 499803 358803 499869 358804
rect 510843 358868 510909 358869
rect 510843 358804 510844 358868
rect 510908 358804 510909 358868
rect 510843 358803 510909 358804
rect 498518 358050 498578 358803
rect 499806 358050 499866 358803
rect 510846 358050 510906 358803
rect 498464 357990 498578 358050
rect 499688 357990 499866 358050
rect 510840 357990 510906 358050
rect 498464 357202 498524 357990
rect 499688 357202 499748 357990
rect 510840 357202 510900 357990
rect 380272 345454 380620 345486
rect 380272 345218 380328 345454
rect 380564 345218 380620 345454
rect 380272 345134 380620 345218
rect 380272 344898 380328 345134
rect 380564 344898 380620 345134
rect 380272 344866 380620 344898
rect 516000 345454 516348 345486
rect 516000 345218 516056 345454
rect 516292 345218 516348 345454
rect 516000 345134 516348 345218
rect 516000 344898 516056 345134
rect 516292 344898 516348 345134
rect 516000 344866 516348 344898
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 380952 327454 381300 327486
rect 380952 327218 381008 327454
rect 381244 327218 381300 327454
rect 380952 327134 381300 327218
rect 380952 326898 381008 327134
rect 381244 326898 381300 327134
rect 380952 326866 381300 326898
rect 515320 327454 515668 327486
rect 515320 327218 515376 327454
rect 515612 327218 515668 327454
rect 515320 327134 515668 327218
rect 515320 326898 515376 327134
rect 515612 326898 515668 327134
rect 515320 326866 515668 326898
rect 380272 309454 380620 309486
rect 380272 309218 380328 309454
rect 380564 309218 380620 309454
rect 380272 309134 380620 309218
rect 380272 308898 380328 309134
rect 380564 308898 380620 309134
rect 380272 308866 380620 308898
rect 516000 309454 516348 309486
rect 516000 309218 516056 309454
rect 516292 309218 516348 309454
rect 516000 309134 516348 309218
rect 516000 308898 516056 309134
rect 516292 308898 516348 309134
rect 516000 308866 516348 308898
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 380952 291454 381300 291486
rect 380952 291218 381008 291454
rect 381244 291218 381300 291454
rect 380952 291134 381300 291218
rect 380952 290898 381008 291134
rect 381244 290898 381300 291134
rect 380952 290866 381300 290898
rect 515320 291454 515668 291486
rect 515320 291218 515376 291454
rect 515612 291218 515668 291454
rect 515320 291134 515668 291218
rect 515320 290898 515376 291134
rect 515612 290898 515668 291134
rect 515320 290866 515668 290898
rect 379470 277350 379714 277410
rect 379470 271557 379530 277350
rect 396056 273730 396116 274040
rect 397144 273730 397204 274040
rect 398232 273730 398292 274040
rect 399592 273730 399652 274040
rect 400544 273730 400604 274040
rect 401768 273730 401828 274040
rect 403128 273730 403188 274040
rect 404216 273730 404276 274040
rect 405440 273730 405500 274040
rect 406528 273730 406588 274040
rect 396030 273670 396116 273730
rect 397134 273670 397204 273730
rect 397502 273670 398292 273730
rect 399526 273670 399652 273730
rect 400446 273670 400604 273730
rect 401734 273670 401828 273730
rect 403022 273670 403188 273730
rect 404126 273670 404276 273730
rect 405046 273670 405500 273730
rect 406518 273670 406588 273730
rect 407616 273730 407676 274040
rect 408296 273730 408356 274040
rect 407616 273670 407682 273730
rect 379467 271556 379533 271557
rect 379467 271492 379468 271556
rect 379532 271492 379533 271556
rect 379467 271491 379533 271492
rect 379794 256394 380414 272000
rect 379794 256158 379826 256394
rect 380062 256158 380146 256394
rect 380382 256158 380414 256394
rect 379794 256074 380414 256158
rect 379794 255838 379826 256074
rect 380062 255838 380146 256074
rect 380382 255838 380414 256074
rect 379794 252308 380414 255838
rect 383514 260114 384134 272000
rect 383514 259878 383546 260114
rect 383782 259878 383866 260114
rect 384102 259878 384134 260114
rect 383514 259794 384134 259878
rect 383514 259558 383546 259794
rect 383782 259558 383866 259794
rect 384102 259558 384134 259794
rect 383514 252308 384134 259558
rect 387234 261954 387854 272000
rect 387234 261718 387266 261954
rect 387502 261718 387586 261954
rect 387822 261718 387854 261954
rect 387234 261634 387854 261718
rect 387234 261398 387266 261634
rect 387502 261398 387586 261634
rect 387822 261398 387854 261634
rect 387234 252308 387854 261398
rect 390954 265674 391574 272000
rect 396030 270605 396090 273670
rect 397134 271285 397194 273670
rect 397131 271284 397197 271285
rect 397131 271220 397132 271284
rect 397196 271220 397197 271284
rect 397131 271219 397197 271220
rect 397502 270605 397562 273670
rect 396027 270604 396093 270605
rect 396027 270540 396028 270604
rect 396092 270540 396093 270604
rect 396027 270539 396093 270540
rect 397499 270604 397565 270605
rect 397499 270540 397500 270604
rect 397564 270540 397565 270604
rect 397499 270539 397565 270540
rect 390954 265438 390986 265674
rect 391222 265438 391306 265674
rect 391542 265438 391574 265674
rect 390954 265354 391574 265438
rect 390954 265118 390986 265354
rect 391222 265118 391306 265354
rect 391542 265118 391574 265354
rect 390954 252308 391574 265118
rect 397794 255454 398414 272000
rect 399526 270605 399586 273670
rect 400446 270605 400506 273670
rect 401734 272237 401794 273670
rect 401731 272236 401797 272237
rect 401731 272172 401732 272236
rect 401796 272172 401797 272236
rect 401731 272171 401797 272172
rect 399523 270604 399589 270605
rect 399523 270540 399524 270604
rect 399588 270540 399589 270604
rect 399523 270539 399589 270540
rect 400443 270604 400509 270605
rect 400443 270540 400444 270604
rect 400508 270540 400509 270604
rect 400443 270539 400509 270540
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 252308 398414 254898
rect 401514 259174 402134 272000
rect 403022 270605 403082 273670
rect 404126 271829 404186 273670
rect 404123 271828 404189 271829
rect 404123 271764 404124 271828
rect 404188 271764 404189 271828
rect 404123 271763 404189 271764
rect 405046 270605 405106 273670
rect 403019 270604 403085 270605
rect 403019 270540 403020 270604
rect 403084 270540 403085 270604
rect 403019 270539 403085 270540
rect 405043 270604 405109 270605
rect 405043 270540 405044 270604
rect 405108 270540 405109 270604
rect 405043 270539 405109 270540
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 252308 402134 258618
rect 405234 262894 405854 272000
rect 406518 270605 406578 273670
rect 407622 270605 407682 273670
rect 408174 273670 408356 273730
rect 408704 273730 408764 274040
rect 410064 273730 410124 274040
rect 408704 273670 408786 273730
rect 408174 271421 408234 273670
rect 408171 271420 408237 271421
rect 408171 271356 408172 271420
rect 408236 271356 408237 271420
rect 408171 271355 408237 271356
rect 408726 270605 408786 273670
rect 410014 273670 410124 273730
rect 410744 273730 410804 274040
rect 411288 273730 411348 274040
rect 412376 273730 412436 274040
rect 413464 273730 413524 274040
rect 410744 273670 410810 273730
rect 411288 273670 411362 273730
rect 412376 273670 412466 273730
rect 406515 270604 406581 270605
rect 406515 270540 406516 270604
rect 406580 270540 406581 270604
rect 406515 270539 406581 270540
rect 407619 270604 407685 270605
rect 407619 270540 407620 270604
rect 407684 270540 407685 270604
rect 407619 270539 407685 270540
rect 408723 270604 408789 270605
rect 408723 270540 408724 270604
rect 408788 270540 408789 270604
rect 408723 270539 408789 270540
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 252308 405854 262338
rect 408954 266614 409574 272000
rect 410014 270605 410074 273670
rect 410750 271013 410810 273670
rect 410747 271012 410813 271013
rect 410747 270948 410748 271012
rect 410812 270948 410813 271012
rect 410747 270947 410813 270948
rect 411302 270741 411362 273670
rect 411299 270740 411365 270741
rect 411299 270676 411300 270740
rect 411364 270676 411365 270740
rect 411299 270675 411365 270676
rect 412406 270605 412466 273670
rect 413326 273670 413524 273730
rect 413600 273730 413660 274040
rect 414552 273730 414612 274040
rect 415912 273730 415972 274040
rect 413600 273670 413754 273730
rect 413326 270605 413386 273670
rect 413694 271557 413754 273670
rect 414430 273670 414612 273730
rect 415534 273670 415972 273730
rect 413691 271556 413757 271557
rect 413691 271492 413692 271556
rect 413756 271492 413757 271556
rect 413691 271491 413757 271492
rect 414430 270605 414490 273670
rect 415534 270605 415594 273670
rect 416048 273597 416108 274040
rect 417000 273730 417060 274040
rect 418088 273730 418148 274040
rect 418496 273730 418556 274040
rect 419448 273730 419508 274040
rect 417000 273670 417066 273730
rect 418088 273670 418170 273730
rect 416045 273596 416111 273597
rect 416045 273532 416046 273596
rect 416110 273532 416111 273596
rect 416045 273531 416111 273532
rect 410011 270604 410077 270605
rect 410011 270540 410012 270604
rect 410076 270540 410077 270604
rect 410011 270539 410077 270540
rect 412403 270604 412469 270605
rect 412403 270540 412404 270604
rect 412468 270540 412469 270604
rect 412403 270539 412469 270540
rect 413323 270604 413389 270605
rect 413323 270540 413324 270604
rect 413388 270540 413389 270604
rect 413323 270539 413389 270540
rect 414427 270604 414493 270605
rect 414427 270540 414428 270604
rect 414492 270540 414493 270604
rect 414427 270539 414493 270540
rect 415531 270604 415597 270605
rect 415531 270540 415532 270604
rect 415596 270540 415597 270604
rect 415531 270539 415597 270540
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 252308 409574 266058
rect 415794 256394 416414 272000
rect 417006 271285 417066 273670
rect 418110 273270 418170 273670
rect 418478 273670 418556 273730
rect 419214 273670 419508 273730
rect 420672 273730 420732 274040
rect 421080 273730 421140 274040
rect 420672 273670 420746 273730
rect 418110 273210 418354 273270
rect 417003 271284 417069 271285
rect 417003 271220 417004 271284
rect 417068 271220 417069 271284
rect 417003 271219 417069 271220
rect 418294 270605 418354 273210
rect 418478 271421 418538 273670
rect 418475 271420 418541 271421
rect 418475 271356 418476 271420
rect 418540 271356 418541 271420
rect 418475 271355 418541 271356
rect 419214 270605 419274 273670
rect 418291 270604 418357 270605
rect 418291 270540 418292 270604
rect 418356 270540 418357 270604
rect 418291 270539 418357 270540
rect 419211 270604 419277 270605
rect 419211 270540 419212 270604
rect 419276 270540 419277 270604
rect 419211 270539 419277 270540
rect 415794 256158 415826 256394
rect 416062 256158 416146 256394
rect 416382 256158 416414 256394
rect 415794 256074 416414 256158
rect 415794 255838 415826 256074
rect 416062 255838 416146 256074
rect 416382 255838 416414 256074
rect 415794 252308 416414 255838
rect 419514 260114 420134 272000
rect 420686 270605 420746 273670
rect 421054 273670 421140 273730
rect 421760 273730 421820 274040
rect 422848 273730 422908 274040
rect 423528 273730 423588 274040
rect 423936 273730 423996 274040
rect 425296 273730 425356 274040
rect 421760 273670 421850 273730
rect 422848 273670 422954 273730
rect 421054 271149 421114 273670
rect 421051 271148 421117 271149
rect 421051 271084 421052 271148
rect 421116 271084 421117 271148
rect 421051 271083 421117 271084
rect 421790 270605 421850 273670
rect 422894 272781 422954 273670
rect 423446 273670 423588 273730
rect 423814 273670 423996 273730
rect 425286 273670 425356 273730
rect 425976 273730 426036 274040
rect 426384 273730 426444 274040
rect 425976 273670 426082 273730
rect 426384 273670 426450 273730
rect 423446 272917 423506 273670
rect 423814 272917 423874 273670
rect 423443 272916 423509 272917
rect 423443 272852 423444 272916
rect 423508 272852 423509 272916
rect 423443 272851 423509 272852
rect 423811 272916 423877 272917
rect 423811 272852 423812 272916
rect 423876 272852 423877 272916
rect 423811 272851 423877 272852
rect 422891 272780 422957 272781
rect 422891 272716 422892 272780
rect 422956 272716 422957 272780
rect 422891 272715 422957 272716
rect 420683 270604 420749 270605
rect 420683 270540 420684 270604
rect 420748 270540 420749 270604
rect 420683 270539 420749 270540
rect 421787 270604 421853 270605
rect 421787 270540 421788 270604
rect 421852 270540 421853 270604
rect 421787 270539 421853 270540
rect 419514 259878 419546 260114
rect 419782 259878 419866 260114
rect 420102 259878 420134 260114
rect 419514 259794 420134 259878
rect 419514 259558 419546 259794
rect 419782 259558 419866 259794
rect 420102 259558 420134 259794
rect 419514 252308 420134 259558
rect 423234 261954 423854 272000
rect 425286 271829 425346 273670
rect 426022 272781 426082 273670
rect 426390 272917 426450 273670
rect 427608 273597 427668 274040
rect 428288 273730 428348 274040
rect 428696 273730 428756 274040
rect 429784 273730 429844 274040
rect 431008 273730 431068 274040
rect 428230 273670 428348 273730
rect 428598 273670 428756 273730
rect 429702 273670 429844 273730
rect 430990 273670 431068 273730
rect 431144 273730 431204 274040
rect 432232 273730 432292 274040
rect 431144 273670 431234 273730
rect 432232 273670 432338 273730
rect 427605 273596 427671 273597
rect 427605 273532 427606 273596
rect 427670 273532 427671 273596
rect 427605 273531 427671 273532
rect 428230 272917 428290 273670
rect 426387 272916 426453 272917
rect 426387 272852 426388 272916
rect 426452 272852 426453 272916
rect 426387 272851 426453 272852
rect 428227 272916 428293 272917
rect 428227 272852 428228 272916
rect 428292 272852 428293 272916
rect 428227 272851 428293 272852
rect 426019 272780 426085 272781
rect 426019 272716 426020 272780
rect 426084 272716 426085 272780
rect 426019 272715 426085 272716
rect 425283 271828 425349 271829
rect 425283 271764 425284 271828
rect 425348 271764 425349 271828
rect 425283 271763 425349 271764
rect 423234 261718 423266 261954
rect 423502 261718 423586 261954
rect 423822 261718 423854 261954
rect 423234 261634 423854 261718
rect 423234 261398 423266 261634
rect 423502 261398 423586 261634
rect 423822 261398 423854 261634
rect 423234 252308 423854 261398
rect 426954 265674 427574 272000
rect 428598 271829 428658 273670
rect 428595 271828 428661 271829
rect 428595 271764 428596 271828
rect 428660 271764 428661 271828
rect 428595 271763 428661 271764
rect 429702 271013 429762 273670
rect 430990 273325 431050 273670
rect 430987 273324 431053 273325
rect 430987 273260 430988 273324
rect 431052 273260 431053 273324
rect 430987 273259 431053 273260
rect 429699 271012 429765 271013
rect 429699 270948 429700 271012
rect 429764 270948 429765 271012
rect 429699 270947 429765 270948
rect 431174 269789 431234 273670
rect 432278 270741 432338 273670
rect 433320 273597 433380 274040
rect 433592 273730 433652 274040
rect 433566 273670 433652 273730
rect 434408 273730 434468 274040
rect 435768 273730 435828 274040
rect 436040 273730 436100 274040
rect 436992 273730 437052 274040
rect 434408 273670 434730 273730
rect 435768 273670 435834 273730
rect 433317 273596 433383 273597
rect 433317 273532 433318 273596
rect 433382 273532 433383 273596
rect 433317 273531 433383 273532
rect 433566 271285 433626 273670
rect 433563 271284 433629 271285
rect 433563 271220 433564 271284
rect 433628 271220 433629 271284
rect 433563 271219 433629 271220
rect 432275 270740 432341 270741
rect 432275 270676 432276 270740
rect 432340 270676 432341 270740
rect 432275 270675 432341 270676
rect 431171 269788 431237 269789
rect 431171 269724 431172 269788
rect 431236 269724 431237 269788
rect 431171 269723 431237 269724
rect 426954 265438 426986 265674
rect 427222 265438 427306 265674
rect 427542 265438 427574 265674
rect 426954 265354 427574 265438
rect 426954 265118 426986 265354
rect 427222 265118 427306 265354
rect 427542 265118 427574 265354
rect 426954 252308 427574 265118
rect 433794 255454 434414 272000
rect 434670 269925 434730 273670
rect 435774 270469 435834 273670
rect 435958 273670 436100 273730
rect 436878 273670 437052 273730
rect 438080 273730 438140 274040
rect 438488 273730 438548 274040
rect 439168 273730 439228 274040
rect 440936 273733 440996 274040
rect 440933 273732 440999 273733
rect 438080 273670 438410 273730
rect 438488 273670 438594 273730
rect 439168 273670 439330 273730
rect 435958 271421 436018 273670
rect 435955 271420 436021 271421
rect 435955 271356 435956 271420
rect 436020 271356 436021 271420
rect 435955 271355 436021 271356
rect 436878 270605 436938 273670
rect 436875 270604 436941 270605
rect 436875 270540 436876 270604
rect 436940 270540 436941 270604
rect 436875 270539 436941 270540
rect 435771 270468 435837 270469
rect 435771 270404 435772 270468
rect 435836 270404 435837 270468
rect 435771 270403 435837 270404
rect 434667 269924 434733 269925
rect 434667 269860 434668 269924
rect 434732 269860 434733 269924
rect 434667 269859 434733 269860
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 252308 434414 254898
rect 437514 259174 438134 272000
rect 438350 271013 438410 273670
rect 438534 271285 438594 273670
rect 439270 271829 439330 273670
rect 440933 273668 440934 273732
rect 440998 273668 440999 273732
rect 443520 273730 443580 274040
rect 445968 273730 446028 274040
rect 440933 273667 440999 273668
rect 443502 273670 443580 273730
rect 445894 273670 446028 273730
rect 448280 273730 448340 274040
rect 451000 273730 451060 274040
rect 453448 273730 453508 274040
rect 455896 273730 455956 274040
rect 458480 273730 458540 274040
rect 448280 273670 448346 273730
rect 451000 273670 451106 273730
rect 439267 271828 439333 271829
rect 439267 271764 439268 271828
rect 439332 271764 439333 271828
rect 439267 271763 439333 271764
rect 438531 271284 438597 271285
rect 438531 271220 438532 271284
rect 438596 271220 438597 271284
rect 438531 271219 438597 271220
rect 438347 271012 438413 271013
rect 438347 270948 438348 271012
rect 438412 270948 438413 271012
rect 438347 270947 438413 270948
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 252308 438134 258618
rect 441234 262894 441854 272000
rect 443502 271557 443562 273670
rect 443499 271556 443565 271557
rect 443499 271492 443500 271556
rect 443564 271492 443565 271556
rect 443499 271491 443565 271492
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 252308 441854 262338
rect 444954 266614 445574 272000
rect 445894 271421 445954 273670
rect 448286 271829 448346 273670
rect 451046 271829 451106 273670
rect 453438 273670 453508 273730
rect 455830 273670 455956 273730
rect 458406 273670 458540 273730
rect 460928 273730 460988 274040
rect 463512 273730 463572 274040
rect 465960 273730 466020 274040
rect 468544 273730 468604 274040
rect 470992 273730 471052 274040
rect 460928 273670 461042 273730
rect 448283 271828 448349 271829
rect 448283 271764 448284 271828
rect 448348 271764 448349 271828
rect 448283 271763 448349 271764
rect 451043 271828 451109 271829
rect 451043 271764 451044 271828
rect 451108 271764 451109 271828
rect 451043 271763 451109 271764
rect 445891 271420 445957 271421
rect 445891 271356 445892 271420
rect 445956 271356 445957 271420
rect 445891 271355 445957 271356
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 252308 445574 266058
rect 451794 256394 452414 272000
rect 453438 271829 453498 273670
rect 455830 272237 455890 273670
rect 455827 272236 455893 272237
rect 455827 272172 455828 272236
rect 455892 272172 455893 272236
rect 455827 272171 455893 272172
rect 453435 271828 453501 271829
rect 453435 271764 453436 271828
rect 453500 271764 453501 271828
rect 453435 271763 453501 271764
rect 451794 256158 451826 256394
rect 452062 256158 452146 256394
rect 452382 256158 452414 256394
rect 451794 256074 452414 256158
rect 451794 255838 451826 256074
rect 452062 255838 452146 256074
rect 452382 255838 452414 256074
rect 451794 252308 452414 255838
rect 455514 260114 456134 272000
rect 458406 271829 458466 273670
rect 458403 271828 458469 271829
rect 458403 271764 458404 271828
rect 458468 271764 458469 271828
rect 458403 271763 458469 271764
rect 455514 259878 455546 260114
rect 455782 259878 455866 260114
rect 456102 259878 456134 260114
rect 455514 259794 456134 259878
rect 455514 259558 455546 259794
rect 455782 259558 455866 259794
rect 456102 259558 456134 259794
rect 455514 252308 456134 259558
rect 459234 261954 459854 272000
rect 460982 271829 461042 273670
rect 462638 273670 463572 273730
rect 465950 273670 466020 273730
rect 468526 273670 468604 273730
rect 470918 273670 471052 273730
rect 473440 273730 473500 274040
rect 475888 273730 475948 274040
rect 478472 273730 478532 274040
rect 480920 273730 480980 274040
rect 483368 273730 483428 274040
rect 473440 273670 473554 273730
rect 460979 271828 461045 271829
rect 460979 271764 460980 271828
rect 461044 271764 461045 271828
rect 460979 271763 461045 271764
rect 462638 270877 462698 273670
rect 462635 270876 462701 270877
rect 462635 270812 462636 270876
rect 462700 270812 462701 270876
rect 462635 270811 462701 270812
rect 459234 261718 459266 261954
rect 459502 261718 459586 261954
rect 459822 261718 459854 261954
rect 459234 261634 459854 261718
rect 459234 261398 459266 261634
rect 459502 261398 459586 261634
rect 459822 261398 459854 261634
rect 459234 252308 459854 261398
rect 462954 265674 463574 272000
rect 465950 271693 466010 273670
rect 468526 272917 468586 273670
rect 470918 272917 470978 273670
rect 468523 272916 468589 272917
rect 468523 272852 468524 272916
rect 468588 272852 468589 272916
rect 468523 272851 468589 272852
rect 470915 272916 470981 272917
rect 470915 272852 470916 272916
rect 470980 272852 470981 272916
rect 470915 272851 470981 272852
rect 473494 272645 473554 273670
rect 475886 273670 475948 273730
rect 478462 273670 478532 273730
rect 480854 273670 480980 273730
rect 483246 273670 483428 273730
rect 485952 273730 486012 274040
rect 503224 273730 503284 274040
rect 485952 273670 486066 273730
rect 475886 272645 475946 273670
rect 478462 272781 478522 273670
rect 480854 272781 480914 273670
rect 483246 273053 483306 273670
rect 486006 273189 486066 273670
rect 503118 273670 503284 273730
rect 503360 273730 503420 274040
rect 503360 273670 503546 273730
rect 486003 273188 486069 273189
rect 486003 273124 486004 273188
rect 486068 273124 486069 273188
rect 486003 273123 486069 273124
rect 483243 273052 483309 273053
rect 483243 272988 483244 273052
rect 483308 272988 483309 273052
rect 483243 272987 483309 272988
rect 478459 272780 478525 272781
rect 478459 272716 478460 272780
rect 478524 272716 478525 272780
rect 478459 272715 478525 272716
rect 480851 272780 480917 272781
rect 480851 272716 480852 272780
rect 480916 272716 480917 272780
rect 480851 272715 480917 272716
rect 473491 272644 473557 272645
rect 473491 272580 473492 272644
rect 473556 272580 473557 272644
rect 473491 272579 473557 272580
rect 475883 272644 475949 272645
rect 475883 272580 475884 272644
rect 475948 272580 475949 272644
rect 475883 272579 475949 272580
rect 465947 271692 466013 271693
rect 465947 271628 465948 271692
rect 466012 271628 466013 271692
rect 465947 271627 466013 271628
rect 462954 265438 462986 265674
rect 463222 265438 463306 265674
rect 463542 265438 463574 265674
rect 462954 265354 463574 265438
rect 462954 265118 462986 265354
rect 463222 265118 463306 265354
rect 463542 265118 463574 265354
rect 462954 252308 463574 265118
rect 469794 255454 470414 272000
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 252308 470414 254898
rect 473514 259174 474134 272000
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 252308 474134 258618
rect 477234 262894 477854 272000
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 252308 477854 262338
rect 480954 266614 481574 272000
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 252308 481574 266058
rect 487794 256394 488414 272000
rect 487794 256158 487826 256394
rect 488062 256158 488146 256394
rect 488382 256158 488414 256394
rect 487794 256074 488414 256158
rect 487794 255838 487826 256074
rect 488062 255838 488146 256074
rect 488382 255838 488414 256074
rect 487794 252308 488414 255838
rect 491514 260114 492134 272000
rect 491514 259878 491546 260114
rect 491782 259878 491866 260114
rect 492102 259878 492134 260114
rect 491514 259794 492134 259878
rect 491514 259558 491546 259794
rect 491782 259558 491866 259794
rect 492102 259558 492134 259794
rect 491514 252308 492134 259558
rect 495234 261954 495854 272000
rect 495234 261718 495266 261954
rect 495502 261718 495586 261954
rect 495822 261718 495854 261954
rect 495234 261634 495854 261718
rect 495234 261398 495266 261634
rect 495502 261398 495586 261634
rect 495822 261398 495854 261634
rect 495234 252308 495854 261398
rect 498954 265674 499574 272000
rect 503118 271421 503178 273670
rect 503486 271557 503546 273670
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 503483 271556 503549 271557
rect 503483 271492 503484 271556
rect 503548 271492 503549 271556
rect 503483 271491 503549 271492
rect 503115 271420 503181 271421
rect 503115 271356 503116 271420
rect 503180 271356 503181 271420
rect 503115 271355 503181 271356
rect 498954 265438 498986 265674
rect 499222 265438 499306 265674
rect 499542 265438 499574 265674
rect 498954 265354 499574 265438
rect 498954 265118 498986 265354
rect 499222 265118 499306 265354
rect 499542 265118 499574 265354
rect 498515 252788 498581 252789
rect 498515 252724 498516 252788
rect 498580 252724 498581 252788
rect 498515 252723 498581 252724
rect 498518 250610 498578 252723
rect 498954 252308 499574 265118
rect 505794 255454 506414 272000
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 499803 253332 499869 253333
rect 499803 253268 499804 253332
rect 499868 253268 499869 253332
rect 499803 253267 499869 253268
rect 499806 250610 499866 253267
rect 505794 252308 506414 254898
rect 509514 259174 510134 272000
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 252308 510134 258618
rect 513234 262894 513854 272000
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 510843 252652 510909 252653
rect 510843 252588 510844 252652
rect 510908 252588 510909 252652
rect 510843 252587 510909 252588
rect 510846 250610 510906 252587
rect 513234 252308 513854 262338
rect 516954 266614 517574 272000
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 252308 517574 266058
rect 498464 250550 498578 250610
rect 499688 250550 499866 250610
rect 510840 250550 510906 250610
rect 498464 250240 498524 250550
rect 499688 250240 499748 250550
rect 510840 250240 510900 250550
rect 380272 237454 380620 237486
rect 380272 237218 380328 237454
rect 380564 237218 380620 237454
rect 380272 237134 380620 237218
rect 380272 236898 380328 237134
rect 380564 236898 380620 237134
rect 380272 236866 380620 236898
rect 516000 237454 516348 237486
rect 516000 237218 516056 237454
rect 516292 237218 516348 237454
rect 516000 237134 516348 237218
rect 516000 236898 516056 237134
rect 516292 236898 516348 237134
rect 516000 236866 516348 236898
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 380952 219454 381300 219486
rect 380952 219218 381008 219454
rect 381244 219218 381300 219454
rect 380952 219134 381300 219218
rect 380952 218898 381008 219134
rect 381244 218898 381300 219134
rect 380952 218866 381300 218898
rect 515320 219454 515668 219486
rect 515320 219218 515376 219454
rect 515612 219218 515668 219454
rect 515320 219134 515668 219218
rect 515320 218898 515376 219134
rect 515612 218898 515668 219134
rect 515320 218866 515668 218898
rect 380272 201454 380620 201486
rect 380272 201218 380328 201454
rect 380564 201218 380620 201454
rect 380272 201134 380620 201218
rect 380272 200898 380328 201134
rect 380564 200898 380620 201134
rect 380272 200866 380620 200898
rect 516000 201454 516348 201486
rect 516000 201218 516056 201454
rect 516292 201218 516348 201454
rect 516000 201134 516348 201218
rect 516000 200898 516056 201134
rect 516292 200898 516348 201134
rect 516000 200866 516348 200898
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 380952 183454 381300 183486
rect 380952 183218 381008 183454
rect 381244 183218 381300 183454
rect 380952 183134 381300 183218
rect 380952 182898 381008 183134
rect 381244 182898 381300 183134
rect 380952 182866 381300 182898
rect 515320 183454 515668 183486
rect 515320 183218 515376 183454
rect 515612 183218 515668 183454
rect 515320 183134 515668 183218
rect 515320 182898 515376 183134
rect 515612 182898 515668 183134
rect 515320 182866 515668 182898
rect 396056 167010 396116 167106
rect 397144 167010 397204 167106
rect 396030 166950 396116 167010
rect 397134 166950 397204 167010
rect 398232 167010 398292 167106
rect 399592 167010 399652 167106
rect 400544 167010 400604 167106
rect 401768 167010 401828 167106
rect 403128 167010 403188 167106
rect 404216 167010 404276 167106
rect 405440 167010 405500 167106
rect 406528 167010 406588 167106
rect 398232 166950 398298 167010
rect 378915 165204 378981 165205
rect 378915 165140 378916 165204
rect 378980 165140 378981 165204
rect 378915 165139 378981 165140
rect 379794 148394 380414 165000
rect 379794 148158 379826 148394
rect 380062 148158 380146 148394
rect 380382 148158 380414 148394
rect 379794 148074 380414 148158
rect 379794 147838 379826 148074
rect 380062 147838 380146 148074
rect 380382 147838 380414 148074
rect 379467 146300 379533 146301
rect 379467 146236 379468 146300
rect 379532 146236 379533 146300
rect 379467 146235 379533 146236
rect 379470 142170 379530 146235
rect 379794 145308 380414 147838
rect 383514 152114 384134 165000
rect 383514 151878 383546 152114
rect 383782 151878 383866 152114
rect 384102 151878 384134 152114
rect 383514 151794 384134 151878
rect 383514 151558 383546 151794
rect 383782 151558 383866 151794
rect 384102 151558 384134 151794
rect 383514 145308 384134 151558
rect 387234 155834 387854 165000
rect 387234 155598 387266 155834
rect 387502 155598 387586 155834
rect 387822 155598 387854 155834
rect 387234 155514 387854 155598
rect 387234 155278 387266 155514
rect 387502 155278 387586 155514
rect 387822 155278 387854 155514
rect 387234 145308 387854 155278
rect 390954 157674 391574 165000
rect 396030 164253 396090 166950
rect 397134 164389 397194 166950
rect 398238 165613 398298 166950
rect 399526 166950 399652 167010
rect 400446 166950 400604 167010
rect 401734 166950 401828 167010
rect 403022 166950 403188 167010
rect 404126 166950 404276 167010
rect 405414 166950 405500 167010
rect 406518 166950 406588 167010
rect 407616 167010 407676 167106
rect 408296 167010 408356 167106
rect 407616 166950 407682 167010
rect 398235 165612 398301 165613
rect 398235 165548 398236 165612
rect 398300 165548 398301 165612
rect 398235 165547 398301 165548
rect 397131 164388 397197 164389
rect 397131 164324 397132 164388
rect 397196 164324 397197 164388
rect 397131 164323 397197 164324
rect 396027 164252 396093 164253
rect 396027 164188 396028 164252
rect 396092 164188 396093 164252
rect 396027 164187 396093 164188
rect 390954 157438 390986 157674
rect 391222 157438 391306 157674
rect 391542 157438 391574 157674
rect 390954 157354 391574 157438
rect 390954 157118 390986 157354
rect 391222 157118 391306 157354
rect 391542 157118 391574 157354
rect 390954 145308 391574 157118
rect 397794 147454 398414 165000
rect 399526 164253 399586 166950
rect 400446 164253 400506 166950
rect 401734 165613 401794 166950
rect 401731 165612 401797 165613
rect 401731 165548 401732 165612
rect 401796 165548 401797 165612
rect 401731 165547 401797 165548
rect 399523 164252 399589 164253
rect 399523 164188 399524 164252
rect 399588 164188 399589 164252
rect 399523 164187 399589 164188
rect 400443 164252 400509 164253
rect 400443 164188 400444 164252
rect 400508 164188 400509 164252
rect 400443 164187 400509 164188
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 145308 398414 146898
rect 401514 151174 402134 165000
rect 403022 164253 403082 166950
rect 404126 164389 404186 166950
rect 405414 165613 405474 166950
rect 405411 165612 405477 165613
rect 405411 165548 405412 165612
rect 405476 165548 405477 165612
rect 405411 165547 405477 165548
rect 404123 164388 404189 164389
rect 404123 164324 404124 164388
rect 404188 164324 404189 164388
rect 404123 164323 404189 164324
rect 403019 164252 403085 164253
rect 403019 164188 403020 164252
rect 403084 164188 403085 164252
rect 403019 164187 403085 164188
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 145308 402134 150618
rect 405234 154894 405854 165000
rect 406518 164253 406578 166950
rect 407622 164253 407682 166950
rect 408174 166950 408356 167010
rect 408174 166293 408234 166950
rect 408171 166292 408237 166293
rect 408171 166228 408172 166292
rect 408236 166228 408237 166292
rect 408704 166290 408764 167106
rect 410064 166290 410124 167106
rect 408704 166230 408786 166290
rect 408171 166227 408237 166228
rect 408726 164253 408786 166230
rect 410014 166230 410124 166290
rect 410744 166290 410804 167106
rect 411288 166290 411348 167106
rect 412376 166290 412436 167106
rect 413464 166290 413524 167106
rect 413600 166565 413660 167106
rect 413597 166564 413663 166565
rect 413597 166500 413598 166564
rect 413662 166500 413663 166564
rect 413597 166499 413663 166500
rect 414552 166290 414612 167106
rect 415912 166290 415972 167106
rect 416048 166837 416108 167106
rect 416045 166836 416111 166837
rect 416045 166772 416046 166836
rect 416110 166772 416111 166836
rect 416045 166771 416111 166772
rect 410744 166230 410810 166290
rect 411288 166230 411362 166290
rect 412376 166230 412466 166290
rect 413464 166230 413570 166290
rect 414552 166230 414674 166290
rect 406515 164252 406581 164253
rect 406515 164188 406516 164252
rect 406580 164188 406581 164252
rect 406515 164187 406581 164188
rect 407619 164252 407685 164253
rect 407619 164188 407620 164252
rect 407684 164188 407685 164252
rect 407619 164187 407685 164188
rect 408723 164252 408789 164253
rect 408723 164188 408724 164252
rect 408788 164188 408789 164252
rect 408723 164187 408789 164188
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 145308 405854 154338
rect 408954 158614 409574 165000
rect 410014 164253 410074 166230
rect 410750 165613 410810 166230
rect 410747 165612 410813 165613
rect 410747 165548 410748 165612
rect 410812 165548 410813 165612
rect 410747 165547 410813 165548
rect 411302 164253 411362 166230
rect 412406 164389 412466 166230
rect 412403 164388 412469 164389
rect 412403 164324 412404 164388
rect 412468 164324 412469 164388
rect 412403 164323 412469 164324
rect 413510 164253 413570 166230
rect 414614 164253 414674 166230
rect 415902 166230 415972 166290
rect 417000 166290 417060 167106
rect 418088 167010 418148 167106
rect 418496 167010 418556 167106
rect 419448 167010 419508 167106
rect 418088 166950 418354 167010
rect 418088 166910 418170 166950
rect 417000 166230 417066 166290
rect 415902 165613 415962 166230
rect 417006 165613 417066 166230
rect 415899 165612 415965 165613
rect 415899 165548 415900 165612
rect 415964 165548 415965 165612
rect 415899 165547 415965 165548
rect 417003 165612 417069 165613
rect 417003 165548 417004 165612
rect 417068 165548 417069 165612
rect 417003 165547 417069 165548
rect 410011 164252 410077 164253
rect 410011 164188 410012 164252
rect 410076 164188 410077 164252
rect 410011 164187 410077 164188
rect 411299 164252 411365 164253
rect 411299 164188 411300 164252
rect 411364 164188 411365 164252
rect 411299 164187 411365 164188
rect 413507 164252 413573 164253
rect 413507 164188 413508 164252
rect 413572 164188 413573 164252
rect 413507 164187 413573 164188
rect 414611 164252 414677 164253
rect 414611 164188 414612 164252
rect 414676 164188 414677 164252
rect 414611 164187 414677 164188
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 145308 409574 158058
rect 415794 148394 416414 165000
rect 418294 164253 418354 166950
rect 418478 166950 418556 167010
rect 419398 166950 419508 167010
rect 420672 167010 420732 167106
rect 421080 167010 421140 167106
rect 420672 166950 420746 167010
rect 418478 166837 418538 166950
rect 418475 166836 418541 166837
rect 418475 166772 418476 166836
rect 418540 166772 418541 166836
rect 418475 166771 418541 166772
rect 419398 165613 419458 166950
rect 419395 165612 419461 165613
rect 419395 165548 419396 165612
rect 419460 165548 419461 165612
rect 419395 165547 419461 165548
rect 418291 164252 418357 164253
rect 418291 164188 418292 164252
rect 418356 164188 418357 164252
rect 418291 164187 418357 164188
rect 415794 148158 415826 148394
rect 416062 148158 416146 148394
rect 416382 148158 416414 148394
rect 415794 148074 416414 148158
rect 415794 147838 415826 148074
rect 416062 147838 416146 148074
rect 416382 147838 416414 148074
rect 415794 145308 416414 147838
rect 419514 152114 420134 165000
rect 420686 164253 420746 166950
rect 421054 166950 421140 167010
rect 421760 167010 421820 167106
rect 422848 167010 422908 167106
rect 423528 167010 423588 167106
rect 423936 167010 423996 167106
rect 425296 167010 425356 167106
rect 421760 166950 421850 167010
rect 422848 166950 422954 167010
rect 421054 164933 421114 166950
rect 421051 164932 421117 164933
rect 421051 164868 421052 164932
rect 421116 164868 421117 164932
rect 421051 164867 421117 164868
rect 421790 164253 421850 166950
rect 422894 164253 422954 166950
rect 423446 166950 423588 167010
rect 423814 166950 423996 167010
rect 425286 166950 425356 167010
rect 425976 167010 426036 167106
rect 426384 167010 426444 167106
rect 427608 167010 427668 167106
rect 428288 167010 428348 167106
rect 425976 166950 426082 167010
rect 426384 166950 426450 167010
rect 423446 166837 423506 166950
rect 423443 166836 423509 166837
rect 423443 166772 423444 166836
rect 423508 166772 423509 166836
rect 423443 166771 423509 166772
rect 423814 165613 423874 166950
rect 423811 165612 423877 165613
rect 423811 165548 423812 165612
rect 423876 165548 423877 165612
rect 423811 165547 423877 165548
rect 420683 164252 420749 164253
rect 420683 164188 420684 164252
rect 420748 164188 420749 164252
rect 420683 164187 420749 164188
rect 421787 164252 421853 164253
rect 421787 164188 421788 164252
rect 421852 164188 421853 164252
rect 421787 164187 421853 164188
rect 422891 164252 422957 164253
rect 422891 164188 422892 164252
rect 422956 164188 422957 164252
rect 422891 164187 422957 164188
rect 419514 151878 419546 152114
rect 419782 151878 419866 152114
rect 420102 151878 420134 152114
rect 419514 151794 420134 151878
rect 419514 151558 419546 151794
rect 419782 151558 419866 151794
rect 420102 151558 420134 151794
rect 419514 145308 420134 151558
rect 423234 155834 423854 165000
rect 425286 164253 425346 166950
rect 426022 166837 426082 166950
rect 426019 166836 426085 166837
rect 426019 166772 426020 166836
rect 426084 166772 426085 166836
rect 426019 166771 426085 166772
rect 426390 164253 426450 166950
rect 427494 166950 427668 167010
rect 428230 166950 428348 167010
rect 428696 167010 428756 167106
rect 429784 167010 429844 167106
rect 431008 167010 431068 167106
rect 428696 166950 428842 167010
rect 427494 165613 427554 166950
rect 428230 166293 428290 166950
rect 428227 166292 428293 166293
rect 428227 166228 428228 166292
rect 428292 166228 428293 166292
rect 428227 166227 428293 166228
rect 427491 165612 427557 165613
rect 427491 165548 427492 165612
rect 427556 165548 427557 165612
rect 427491 165547 427557 165548
rect 425283 164252 425349 164253
rect 425283 164188 425284 164252
rect 425348 164188 425349 164252
rect 425283 164187 425349 164188
rect 426387 164252 426453 164253
rect 426387 164188 426388 164252
rect 426452 164188 426453 164252
rect 426387 164187 426453 164188
rect 423234 155598 423266 155834
rect 423502 155598 423586 155834
rect 423822 155598 423854 155834
rect 423234 155514 423854 155598
rect 423234 155278 423266 155514
rect 423502 155278 423586 155514
rect 423822 155278 423854 155514
rect 423234 145308 423854 155278
rect 426954 157674 427574 165000
rect 428782 164253 428842 166950
rect 429702 166950 429844 167010
rect 430990 166950 431068 167010
rect 431144 167010 431204 167106
rect 432232 167010 432292 167106
rect 433320 167010 433380 167106
rect 433592 167010 433652 167106
rect 431144 166950 431234 167010
rect 432232 166950 432338 167010
rect 433320 166950 433442 167010
rect 429702 164389 429762 166950
rect 429699 164388 429765 164389
rect 429699 164324 429700 164388
rect 429764 164324 429765 164388
rect 429699 164323 429765 164324
rect 430990 164253 431050 166950
rect 431174 164389 431234 166950
rect 431171 164388 431237 164389
rect 431171 164324 431172 164388
rect 431236 164324 431237 164388
rect 431171 164323 431237 164324
rect 432278 164253 432338 166950
rect 433382 165613 433442 166950
rect 433566 166950 433652 167010
rect 434408 167010 434468 167106
rect 435768 167010 435828 167106
rect 436040 167010 436100 167106
rect 436992 167010 437052 167106
rect 438080 167010 438140 167106
rect 434408 166950 434730 167010
rect 435768 166950 435834 167010
rect 433379 165612 433445 165613
rect 433379 165548 433380 165612
rect 433444 165548 433445 165612
rect 433379 165547 433445 165548
rect 433566 164933 433626 166950
rect 433563 164932 433629 164933
rect 433563 164868 433564 164932
rect 433628 164868 433629 164932
rect 433563 164867 433629 164868
rect 428779 164252 428845 164253
rect 428779 164188 428780 164252
rect 428844 164188 428845 164252
rect 428779 164187 428845 164188
rect 430987 164252 431053 164253
rect 430987 164188 430988 164252
rect 431052 164188 431053 164252
rect 430987 164187 431053 164188
rect 432275 164252 432341 164253
rect 432275 164188 432276 164252
rect 432340 164188 432341 164252
rect 432275 164187 432341 164188
rect 426954 157438 426986 157674
rect 427222 157438 427306 157674
rect 427542 157438 427574 157674
rect 426954 157354 427574 157438
rect 426954 157118 426986 157354
rect 427222 157118 427306 157354
rect 427542 157118 427574 157354
rect 426954 145308 427574 157118
rect 433794 147454 434414 165000
rect 434670 164661 434730 166950
rect 434667 164660 434733 164661
rect 434667 164596 434668 164660
rect 434732 164596 434733 164660
rect 434667 164595 434733 164596
rect 435774 164253 435834 166950
rect 435958 166950 436100 167010
rect 436878 166950 437052 167010
rect 437982 166950 438140 167010
rect 438488 167010 438548 167106
rect 439168 167010 439228 167106
rect 440936 167010 440996 167106
rect 443520 167010 443580 167106
rect 445968 167010 446028 167106
rect 438488 166950 438594 167010
rect 439168 166950 439330 167010
rect 435958 165613 436018 166950
rect 435955 165612 436021 165613
rect 435955 165548 435956 165612
rect 436020 165548 436021 165612
rect 435955 165547 436021 165548
rect 436878 164253 436938 166950
rect 437982 165613 438042 166950
rect 437979 165612 438045 165613
rect 437979 165548 437980 165612
rect 438044 165548 438045 165612
rect 437979 165547 438045 165548
rect 438534 165069 438594 166950
rect 438531 165068 438597 165069
rect 438531 165004 438532 165068
rect 438596 165004 438597 165068
rect 438531 165003 438597 165004
rect 435771 164252 435837 164253
rect 435771 164188 435772 164252
rect 435836 164188 435837 164252
rect 435771 164187 435837 164188
rect 436875 164252 436941 164253
rect 436875 164188 436876 164252
rect 436940 164188 436941 164252
rect 436875 164187 436941 164188
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 145308 434414 146898
rect 437514 151174 438134 165000
rect 439270 164253 439330 166950
rect 440926 166950 440996 167010
rect 443502 166950 443580 167010
rect 445894 166950 446028 167010
rect 448280 167010 448340 167106
rect 451000 167010 451060 167106
rect 453448 167010 453508 167106
rect 455896 167010 455956 167106
rect 448280 166950 448346 167010
rect 451000 166950 451106 167010
rect 440926 165613 440986 166950
rect 443502 165613 443562 166950
rect 440923 165612 440989 165613
rect 440923 165548 440924 165612
rect 440988 165548 440989 165612
rect 440923 165547 440989 165548
rect 443499 165612 443565 165613
rect 443499 165548 443500 165612
rect 443564 165548 443565 165612
rect 443499 165547 443565 165548
rect 445894 165069 445954 166950
rect 448286 165613 448346 166950
rect 451046 165613 451106 166950
rect 453438 166950 453508 167010
rect 455830 166950 455956 167010
rect 453438 165613 453498 166950
rect 455830 165613 455890 166950
rect 458480 166290 458540 167106
rect 458406 166230 458540 166290
rect 460928 166290 460988 167106
rect 463512 166290 463572 167106
rect 465960 166290 466020 167106
rect 468544 166290 468604 167106
rect 470992 166837 471052 167106
rect 473440 166837 473500 167106
rect 475888 166837 475948 167106
rect 478472 166837 478532 167106
rect 480920 166837 480980 167106
rect 470989 166836 471055 166837
rect 470989 166772 470990 166836
rect 471054 166772 471055 166836
rect 470989 166771 471055 166772
rect 473437 166836 473503 166837
rect 473437 166772 473438 166836
rect 473502 166772 473503 166836
rect 473437 166771 473503 166772
rect 475885 166836 475951 166837
rect 475885 166772 475886 166836
rect 475950 166772 475951 166836
rect 475885 166771 475951 166772
rect 478469 166836 478535 166837
rect 478469 166772 478470 166836
rect 478534 166772 478535 166836
rect 478469 166771 478535 166772
rect 480917 166836 480983 166837
rect 480917 166772 480918 166836
rect 480982 166772 480983 166836
rect 480917 166771 480983 166772
rect 483368 166701 483428 167106
rect 485952 166701 486012 167106
rect 483365 166700 483431 166701
rect 483365 166636 483366 166700
rect 483430 166636 483431 166700
rect 483365 166635 483431 166636
rect 485949 166700 486015 166701
rect 485949 166636 485950 166700
rect 486014 166636 486015 166700
rect 485949 166635 486015 166636
rect 503224 166565 503284 167106
rect 503221 166564 503287 166565
rect 503221 166500 503222 166564
rect 503286 166500 503287 166564
rect 503221 166499 503287 166500
rect 503360 166290 503420 167106
rect 460928 166230 461042 166290
rect 463512 166230 463618 166290
rect 458406 165613 458466 166230
rect 448283 165612 448349 165613
rect 448283 165548 448284 165612
rect 448348 165548 448349 165612
rect 448283 165547 448349 165548
rect 451043 165612 451109 165613
rect 451043 165548 451044 165612
rect 451108 165548 451109 165612
rect 451043 165547 451109 165548
rect 453435 165612 453501 165613
rect 453435 165548 453436 165612
rect 453500 165548 453501 165612
rect 453435 165547 453501 165548
rect 455827 165612 455893 165613
rect 455827 165548 455828 165612
rect 455892 165548 455893 165612
rect 455827 165547 455893 165548
rect 458403 165612 458469 165613
rect 458403 165548 458404 165612
rect 458468 165548 458469 165612
rect 458403 165547 458469 165548
rect 445891 165068 445957 165069
rect 445891 165004 445892 165068
rect 445956 165004 445957 165068
rect 445891 165003 445957 165004
rect 439267 164252 439333 164253
rect 439267 164188 439268 164252
rect 439332 164188 439333 164252
rect 439267 164187 439333 164188
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 145308 438134 150618
rect 441234 154894 441854 165000
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 145308 441854 154338
rect 444954 158614 445574 165000
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 145308 445574 158058
rect 451794 148394 452414 165000
rect 451794 148158 451826 148394
rect 452062 148158 452146 148394
rect 452382 148158 452414 148394
rect 451794 148074 452414 148158
rect 451794 147838 451826 148074
rect 452062 147838 452146 148074
rect 452382 147838 452414 148074
rect 451794 145308 452414 147838
rect 455514 152114 456134 165000
rect 455514 151878 455546 152114
rect 455782 151878 455866 152114
rect 456102 151878 456134 152114
rect 455514 151794 456134 151878
rect 455514 151558 455546 151794
rect 455782 151558 455866 151794
rect 456102 151558 456134 151794
rect 455514 145308 456134 151558
rect 459234 155834 459854 165000
rect 460982 164797 461042 166230
rect 463558 165205 463618 166230
rect 465950 166230 466020 166290
rect 468526 166230 468604 166290
rect 503302 166230 503420 166290
rect 465950 165341 466010 166230
rect 468526 165477 468586 166230
rect 468523 165476 468589 165477
rect 468523 165412 468524 165476
rect 468588 165412 468589 165476
rect 468523 165411 468589 165412
rect 465947 165340 466013 165341
rect 465947 165276 465948 165340
rect 466012 165276 466013 165340
rect 465947 165275 466013 165276
rect 463555 165204 463621 165205
rect 463555 165140 463556 165204
rect 463620 165140 463621 165204
rect 463555 165139 463621 165140
rect 460979 164796 461045 164797
rect 460979 164732 460980 164796
rect 461044 164732 461045 164796
rect 460979 164731 461045 164732
rect 459234 155598 459266 155834
rect 459502 155598 459586 155834
rect 459822 155598 459854 155834
rect 459234 155514 459854 155598
rect 459234 155278 459266 155514
rect 459502 155278 459586 155514
rect 459822 155278 459854 155514
rect 459234 145308 459854 155278
rect 462954 157674 463574 165000
rect 462954 157438 462986 157674
rect 463222 157438 463306 157674
rect 463542 157438 463574 157674
rect 462954 157354 463574 157438
rect 462954 157118 462986 157354
rect 463222 157118 463306 157354
rect 463542 157118 463574 157354
rect 462954 145308 463574 157118
rect 469794 147454 470414 165000
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 145308 470414 146898
rect 473514 151174 474134 165000
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 145308 474134 150618
rect 477234 154894 477854 165000
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 145308 477854 154338
rect 480954 158614 481574 165000
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 145308 481574 158058
rect 487794 148394 488414 165000
rect 487794 148158 487826 148394
rect 488062 148158 488146 148394
rect 488382 148158 488414 148394
rect 487794 148074 488414 148158
rect 487794 147838 487826 148074
rect 488062 147838 488146 148074
rect 488382 147838 488414 148074
rect 487794 145308 488414 147838
rect 491514 152114 492134 165000
rect 491514 151878 491546 152114
rect 491782 151878 491866 152114
rect 492102 151878 492134 152114
rect 491514 151794 492134 151878
rect 491514 151558 491546 151794
rect 491782 151558 491866 151794
rect 492102 151558 492134 151794
rect 491514 145308 492134 151558
rect 495234 155834 495854 165000
rect 495234 155598 495266 155834
rect 495502 155598 495586 155834
rect 495822 155598 495854 155834
rect 495234 155514 495854 155598
rect 495234 155278 495266 155514
rect 495502 155278 495586 155514
rect 495822 155278 495854 155514
rect 495234 145308 495854 155278
rect 498954 157674 499574 165000
rect 503302 164661 503362 166230
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 503299 164660 503365 164661
rect 503299 164596 503300 164660
rect 503364 164596 503365 164660
rect 503299 164595 503365 164596
rect 498954 157438 498986 157674
rect 499222 157438 499306 157674
rect 499542 157438 499574 157674
rect 498954 157354 499574 157438
rect 498954 157118 498986 157354
rect 499222 157118 499306 157354
rect 499542 157118 499574 157354
rect 498954 145308 499574 157118
rect 505794 147454 506414 165000
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 145308 506414 146898
rect 509514 151174 510134 165000
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 145308 510134 150618
rect 513234 154894 513854 165000
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 510843 146164 510909 146165
rect 510843 146100 510844 146164
rect 510908 146100 510909 146164
rect 510843 146099 510909 146100
rect 498515 144940 498581 144941
rect 498515 144876 498516 144940
rect 498580 144876 498581 144940
rect 498515 144875 498581 144876
rect 499803 144940 499869 144941
rect 499803 144876 499804 144940
rect 499868 144876 499869 144940
rect 499803 144875 499869 144876
rect 498518 143850 498578 144875
rect 499806 143850 499866 144875
rect 510846 143850 510906 146099
rect 513234 145308 513854 154338
rect 516954 158614 517574 165000
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 145308 517574 158058
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 498464 143790 498578 143850
rect 499688 143790 499866 143850
rect 510840 143790 510906 143850
rect 498464 143202 498524 143790
rect 499688 143202 499748 143790
rect 510840 143202 510900 143790
rect 379470 142110 379714 142170
rect 378731 57220 378797 57221
rect 378731 57156 378732 57220
rect 378796 57156 378797 57220
rect 378731 57155 378797 57156
rect 379654 55230 379714 142110
rect 380272 129454 380620 129486
rect 380272 129218 380328 129454
rect 380564 129218 380620 129454
rect 380272 129134 380620 129218
rect 380272 128898 380328 129134
rect 380564 128898 380620 129134
rect 380272 128866 380620 128898
rect 516000 129454 516348 129486
rect 516000 129218 516056 129454
rect 516292 129218 516348 129454
rect 516000 129134 516348 129218
rect 516000 128898 516056 129134
rect 516292 128898 516348 129134
rect 516000 128866 516348 128898
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 380952 111454 381300 111486
rect 380952 111218 381008 111454
rect 381244 111218 381300 111454
rect 380952 111134 381300 111218
rect 380952 110898 381008 111134
rect 381244 110898 381300 111134
rect 380952 110866 381300 110898
rect 515320 111454 515668 111486
rect 515320 111218 515376 111454
rect 515612 111218 515668 111454
rect 515320 111134 515668 111218
rect 515320 110898 515376 111134
rect 515612 110898 515668 111134
rect 515320 110866 515668 110898
rect 380272 93454 380620 93486
rect 380272 93218 380328 93454
rect 380564 93218 380620 93454
rect 380272 93134 380620 93218
rect 380272 92898 380328 93134
rect 380564 92898 380620 93134
rect 380272 92866 380620 92898
rect 516000 93454 516348 93486
rect 516000 93218 516056 93454
rect 516292 93218 516348 93454
rect 516000 93134 516348 93218
rect 516000 92898 516056 93134
rect 516292 92898 516348 93134
rect 516000 92866 516348 92898
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 380952 75454 381300 75486
rect 380952 75218 381008 75454
rect 381244 75218 381300 75454
rect 380952 75134 381300 75218
rect 380952 74898 381008 75134
rect 381244 74898 381300 75134
rect 380952 74866 381300 74898
rect 515320 75454 515668 75486
rect 515320 75218 515376 75454
rect 515612 75218 515668 75454
rect 515320 75134 515668 75218
rect 515320 74898 515376 75134
rect 515612 74898 515668 75134
rect 515320 74866 515668 74898
rect 396056 59805 396116 60106
rect 397144 59805 397204 60106
rect 396053 59804 396119 59805
rect 396053 59740 396054 59804
rect 396118 59740 396119 59804
rect 396053 59739 396119 59740
rect 397141 59804 397207 59805
rect 397141 59740 397142 59804
rect 397206 59740 397207 59804
rect 398232 59802 398292 60106
rect 399592 59802 399652 60106
rect 400544 59802 400604 60106
rect 398232 59742 398298 59802
rect 397141 59739 397207 59740
rect 398238 59397 398298 59742
rect 399526 59742 399652 59802
rect 400446 59742 400604 59802
rect 398235 59396 398301 59397
rect 398235 59332 398236 59396
rect 398300 59332 398301 59396
rect 398235 59331 398301 59332
rect 377811 55180 377877 55181
rect 377811 55116 377812 55180
rect 377876 55116 377877 55180
rect 377811 55115 377877 55116
rect 379470 55170 379714 55230
rect 379794 57454 380414 58000
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379470 55045 379530 55170
rect 379467 55044 379533 55045
rect 379467 54980 379468 55044
rect 379532 54980 379533 55044
rect 379467 54979 379533 54980
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 371739 3636 371805 3637
rect 371739 3572 371740 3636
rect 371804 3572 371805 3636
rect 371739 3571 371805 3572
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 25174 384134 58000
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 28894 387854 58000
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 32614 391574 58000
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 39454 398414 58000
rect 399526 57901 399586 59742
rect 400446 57901 400506 59742
rect 401768 59530 401828 60106
rect 403128 59805 403188 60106
rect 403125 59804 403191 59805
rect 403125 59740 403126 59804
rect 403190 59740 403191 59804
rect 403125 59739 403191 59740
rect 404216 59530 404276 60106
rect 405440 59530 405500 60106
rect 406528 59530 406588 60106
rect 401734 59470 401828 59530
rect 404126 59470 404276 59530
rect 405046 59470 405500 59530
rect 406518 59470 406588 59530
rect 407616 59530 407676 60106
rect 408296 59530 408356 60106
rect 408704 59530 408764 60106
rect 410064 59530 410124 60106
rect 407616 59470 407682 59530
rect 408296 59470 408418 59530
rect 408704 59470 408786 59530
rect 401734 58173 401794 59470
rect 401731 58172 401797 58173
rect 401731 58108 401732 58172
rect 401796 58108 401797 58172
rect 401731 58107 401797 58108
rect 399523 57900 399589 57901
rect 399523 57836 399524 57900
rect 399588 57836 399589 57900
rect 399523 57835 399589 57836
rect 400443 57900 400509 57901
rect 400443 57836 400444 57900
rect 400508 57836 400509 57900
rect 400443 57835 400509 57836
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 43174 402134 58000
rect 404126 57901 404186 59470
rect 405046 57901 405106 59470
rect 404123 57900 404189 57901
rect 404123 57836 404124 57900
rect 404188 57836 404189 57900
rect 404123 57835 404189 57836
rect 405043 57900 405109 57901
rect 405043 57836 405044 57900
rect 405108 57836 405109 57900
rect 405043 57835 405109 57836
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 46894 405854 58000
rect 406518 57901 406578 59470
rect 407622 57901 407682 59470
rect 408358 57901 408418 59470
rect 408726 57901 408786 59470
rect 410014 59470 410124 59530
rect 410744 59530 410804 60106
rect 411288 59530 411348 60106
rect 412376 59530 412436 60106
rect 413464 59530 413524 60106
rect 413600 59805 413660 60106
rect 413597 59804 413663 59805
rect 413597 59740 413598 59804
rect 413662 59740 413663 59804
rect 413597 59739 413663 59740
rect 414552 59530 414612 60106
rect 415912 59805 415972 60106
rect 415909 59804 415975 59805
rect 415909 59740 415910 59804
rect 415974 59740 415975 59804
rect 415909 59739 415975 59740
rect 416048 59530 416108 60106
rect 410744 59470 410810 59530
rect 411288 59470 411362 59530
rect 412376 59470 412466 59530
rect 413464 59470 413570 59530
rect 414552 59470 414674 59530
rect 406515 57900 406581 57901
rect 406515 57836 406516 57900
rect 406580 57836 406581 57900
rect 406515 57835 406581 57836
rect 407619 57900 407685 57901
rect 407619 57836 407620 57900
rect 407684 57836 407685 57900
rect 407619 57835 407685 57836
rect 408355 57900 408421 57901
rect 408355 57836 408356 57900
rect 408420 57836 408421 57900
rect 408355 57835 408421 57836
rect 408723 57900 408789 57901
rect 408723 57836 408724 57900
rect 408788 57836 408789 57900
rect 408723 57835 408789 57836
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 50614 409574 58000
rect 410014 57901 410074 59470
rect 410750 59397 410810 59470
rect 410747 59396 410813 59397
rect 410747 59332 410748 59396
rect 410812 59332 410813 59396
rect 410747 59331 410813 59332
rect 410011 57900 410077 57901
rect 410011 57836 410012 57900
rect 410076 57836 410077 57900
rect 410011 57835 410077 57836
rect 411302 56949 411362 59470
rect 412406 57901 412466 59470
rect 413510 57901 413570 59470
rect 414614 57901 414674 59470
rect 415534 59470 416108 59530
rect 417000 59530 417060 60106
rect 418088 59530 418148 60106
rect 418496 59530 418556 60106
rect 419448 59805 419508 60106
rect 419445 59804 419511 59805
rect 419445 59740 419446 59804
rect 419510 59740 419511 59804
rect 419445 59739 419511 59740
rect 417000 59470 417066 59530
rect 418088 59470 418170 59530
rect 412403 57900 412469 57901
rect 412403 57836 412404 57900
rect 412468 57836 412469 57900
rect 412403 57835 412469 57836
rect 413507 57900 413573 57901
rect 413507 57836 413508 57900
rect 413572 57836 413573 57900
rect 413507 57835 413573 57836
rect 414611 57900 414677 57901
rect 414611 57836 414612 57900
rect 414676 57836 414677 57900
rect 414611 57835 414677 57836
rect 415534 57085 415594 59470
rect 417006 59397 417066 59470
rect 418110 59397 418170 59470
rect 418478 59470 418556 59530
rect 420672 59530 420732 60106
rect 421080 59530 421140 60106
rect 420672 59470 420746 59530
rect 417003 59396 417069 59397
rect 417003 59332 417004 59396
rect 417068 59332 417069 59396
rect 417003 59331 417069 59332
rect 418107 59396 418173 59397
rect 418107 59332 418108 59396
rect 418172 59332 418173 59396
rect 418107 59331 418173 59332
rect 415794 57454 416414 58000
rect 418478 57901 418538 59470
rect 420686 58445 420746 59470
rect 421054 59470 421140 59530
rect 421760 59530 421820 60106
rect 422848 59530 422908 60106
rect 423528 59669 423588 60106
rect 423525 59668 423591 59669
rect 423525 59604 423526 59668
rect 423590 59604 423591 59668
rect 423525 59603 423591 59604
rect 423936 59530 423996 60106
rect 425296 59530 425356 60106
rect 421760 59470 421850 59530
rect 422848 59470 422954 59530
rect 423936 59470 424058 59530
rect 421054 59397 421114 59470
rect 421790 59397 421850 59470
rect 421051 59396 421117 59397
rect 421051 59332 421052 59396
rect 421116 59332 421117 59396
rect 421051 59331 421117 59332
rect 421787 59396 421853 59397
rect 421787 59332 421788 59396
rect 421852 59332 421853 59396
rect 421787 59331 421853 59332
rect 420683 58444 420749 58445
rect 420683 58380 420684 58444
rect 420748 58380 420749 58444
rect 420683 58379 420749 58380
rect 418475 57900 418541 57901
rect 418475 57836 418476 57900
rect 418540 57836 418541 57900
rect 418475 57835 418541 57836
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415531 57084 415597 57085
rect 415531 57020 415532 57084
rect 415596 57020 415597 57084
rect 415531 57019 415597 57020
rect 411299 56948 411365 56949
rect 411299 56884 411300 56948
rect 411364 56884 411365 56948
rect 411299 56883 411365 56884
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 25174 420134 58000
rect 422894 57901 422954 59470
rect 422891 57900 422957 57901
rect 422891 57836 422892 57900
rect 422956 57836 422957 57900
rect 422891 57835 422957 57836
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 28894 423854 58000
rect 423998 57901 424058 59470
rect 425286 59470 425356 59530
rect 425976 59530 426036 60106
rect 426384 59530 426444 60106
rect 427608 59530 427668 60106
rect 428288 59530 428348 60106
rect 428696 59530 428756 60106
rect 429784 59530 429844 60106
rect 431008 59530 431068 60106
rect 425976 59470 426082 59530
rect 426384 59470 426450 59530
rect 427608 59470 427738 59530
rect 425286 59397 425346 59470
rect 426022 59397 426082 59470
rect 425283 59396 425349 59397
rect 425283 59332 425284 59396
rect 425348 59332 425349 59396
rect 425283 59331 425349 59332
rect 426019 59396 426085 59397
rect 426019 59332 426020 59396
rect 426084 59332 426085 59396
rect 426019 59331 426085 59332
rect 426390 57901 426450 59470
rect 423995 57900 424061 57901
rect 423995 57836 423996 57900
rect 424060 57836 424061 57900
rect 423995 57835 424061 57836
rect 426387 57900 426453 57901
rect 426387 57836 426388 57900
rect 426452 57836 426453 57900
rect 426387 57835 426453 57836
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 32614 427574 58000
rect 427678 57901 427738 59470
rect 428230 59470 428348 59530
rect 428598 59470 428756 59530
rect 429702 59470 429844 59530
rect 430990 59470 431068 59530
rect 431144 59530 431204 60106
rect 432232 59530 432292 60106
rect 433320 59530 433380 60106
rect 433592 59530 433652 60106
rect 431144 59470 431234 59530
rect 432232 59470 432338 59530
rect 433320 59470 433442 59530
rect 428230 59397 428290 59470
rect 428227 59396 428293 59397
rect 428227 59332 428228 59396
rect 428292 59332 428293 59396
rect 428227 59331 428293 59332
rect 428598 57901 428658 59470
rect 429702 57901 429762 59470
rect 430990 57901 431050 59470
rect 427675 57900 427741 57901
rect 427675 57836 427676 57900
rect 427740 57836 427741 57900
rect 427675 57835 427741 57836
rect 428595 57900 428661 57901
rect 428595 57836 428596 57900
rect 428660 57836 428661 57900
rect 428595 57835 428661 57836
rect 429699 57900 429765 57901
rect 429699 57836 429700 57900
rect 429764 57836 429765 57900
rect 429699 57835 429765 57836
rect 430987 57900 431053 57901
rect 430987 57836 430988 57900
rect 431052 57836 431053 57900
rect 430987 57835 431053 57836
rect 431174 57085 431234 59470
rect 432278 57901 432338 59470
rect 433382 57901 433442 59470
rect 433566 59470 433652 59530
rect 434408 59530 434468 60106
rect 435768 59530 435828 60106
rect 436040 59530 436100 60106
rect 436992 59530 437052 60106
rect 434408 59470 434730 59530
rect 435768 59470 435834 59530
rect 433566 57901 433626 59470
rect 432275 57900 432341 57901
rect 432275 57836 432276 57900
rect 432340 57836 432341 57900
rect 432275 57835 432341 57836
rect 433379 57900 433445 57901
rect 433379 57836 433380 57900
rect 433444 57836 433445 57900
rect 433379 57835 433445 57836
rect 433563 57900 433629 57901
rect 433563 57836 433564 57900
rect 433628 57836 433629 57900
rect 433563 57835 433629 57836
rect 431171 57084 431237 57085
rect 431171 57020 431172 57084
rect 431236 57020 431237 57084
rect 431171 57019 431237 57020
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 39454 434414 58000
rect 434670 57493 434730 59470
rect 435774 57901 435834 59470
rect 435958 59470 436100 59530
rect 436878 59470 437052 59530
rect 438080 59530 438140 60106
rect 438488 59530 438548 60106
rect 439168 59530 439228 60106
rect 440936 59530 440996 60106
rect 443520 59530 443580 60106
rect 445968 59530 446028 60106
rect 438080 59470 438410 59530
rect 438488 59470 438594 59530
rect 435958 57901 436018 59470
rect 435771 57900 435837 57901
rect 435771 57836 435772 57900
rect 435836 57836 435837 57900
rect 435771 57835 435837 57836
rect 435955 57900 436021 57901
rect 435955 57836 435956 57900
rect 436020 57836 436021 57900
rect 435955 57835 436021 57836
rect 436878 57493 436938 59470
rect 434667 57492 434733 57493
rect 434667 57428 434668 57492
rect 434732 57428 434733 57492
rect 434667 57427 434733 57428
rect 436875 57492 436941 57493
rect 436875 57428 436876 57492
rect 436940 57428 436941 57492
rect 436875 57427 436941 57428
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 43174 438134 58000
rect 438350 56677 438410 59470
rect 438534 57901 438594 59470
rect 439086 59470 439228 59530
rect 440926 59470 440996 59530
rect 443502 59470 443580 59530
rect 445894 59470 446028 59530
rect 448280 59530 448340 60106
rect 451000 59530 451060 60106
rect 453448 59530 453508 60106
rect 455896 59530 455956 60106
rect 458480 59530 458540 60106
rect 448280 59470 448346 59530
rect 451000 59470 451106 59530
rect 438531 57900 438597 57901
rect 438531 57836 438532 57900
rect 438596 57836 438597 57900
rect 438531 57835 438597 57836
rect 439086 57493 439146 59470
rect 439083 57492 439149 57493
rect 439083 57428 439084 57492
rect 439148 57428 439149 57492
rect 439083 57427 439149 57428
rect 440926 57085 440986 59470
rect 440923 57084 440989 57085
rect 440923 57020 440924 57084
rect 440988 57020 440989 57084
rect 440923 57019 440989 57020
rect 438347 56676 438413 56677
rect 438347 56612 438348 56676
rect 438412 56612 438413 56676
rect 438347 56611 438413 56612
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 46894 441854 58000
rect 443502 56813 443562 59470
rect 443499 56812 443565 56813
rect 443499 56748 443500 56812
rect 443564 56748 443565 56812
rect 443499 56747 443565 56748
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 50614 445574 58000
rect 445894 57221 445954 59470
rect 448286 57357 448346 59470
rect 451046 57629 451106 59470
rect 453438 59470 453508 59530
rect 455830 59470 455956 59530
rect 458406 59470 458540 59530
rect 460928 59530 460988 60106
rect 463512 59530 463572 60106
rect 465960 59530 466020 60106
rect 468544 59530 468604 60106
rect 470992 59530 471052 60106
rect 460928 59470 461042 59530
rect 463512 59470 463618 59530
rect 453438 58581 453498 59470
rect 453435 58580 453501 58581
rect 453435 58516 453436 58580
rect 453500 58516 453501 58580
rect 453435 58515 453501 58516
rect 455830 58173 455890 59470
rect 458406 58853 458466 59470
rect 458403 58852 458469 58853
rect 458403 58788 458404 58852
rect 458468 58788 458469 58852
rect 458403 58787 458469 58788
rect 455827 58172 455893 58173
rect 455827 58108 455828 58172
rect 455892 58108 455893 58172
rect 455827 58107 455893 58108
rect 451043 57628 451109 57629
rect 451043 57564 451044 57628
rect 451108 57564 451109 57628
rect 451043 57563 451109 57564
rect 451794 57454 452414 58000
rect 448283 57356 448349 57357
rect 448283 57292 448284 57356
rect 448348 57292 448349 57356
rect 448283 57291 448349 57292
rect 445891 57220 445957 57221
rect 445891 57156 445892 57220
rect 445956 57156 445957 57220
rect 445891 57155 445957 57156
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 25174 456134 58000
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 28894 459854 58000
rect 460982 57901 461042 59470
rect 463558 58717 463618 59470
rect 465950 59470 466020 59530
rect 468526 59470 468604 59530
rect 470918 59470 471052 59530
rect 473440 59530 473500 60106
rect 475888 59530 475948 60106
rect 478472 59530 478532 60106
rect 480920 59530 480980 60106
rect 473440 59470 473554 59530
rect 463555 58716 463621 58717
rect 463555 58652 463556 58716
rect 463620 58652 463621 58716
rect 463555 58651 463621 58652
rect 460979 57900 461045 57901
rect 460979 57836 460980 57900
rect 461044 57836 461045 57900
rect 460979 57835 461045 57836
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 32614 463574 58000
rect 465950 57901 466010 59470
rect 468526 59397 468586 59470
rect 468523 59396 468589 59397
rect 468523 59332 468524 59396
rect 468588 59332 468589 59396
rect 468523 59331 468589 59332
rect 465947 57900 466013 57901
rect 465947 57836 465948 57900
rect 466012 57836 466013 57900
rect 465947 57835 466013 57836
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 39454 470414 58000
rect 470918 57901 470978 59470
rect 473494 58989 473554 59470
rect 475886 59470 475948 59530
rect 478462 59470 478532 59530
rect 480670 59470 480980 59530
rect 483368 59530 483428 60106
rect 485952 59530 486012 60106
rect 503224 59669 503284 60106
rect 503221 59668 503287 59669
rect 503221 59604 503222 59668
rect 503286 59604 503287 59668
rect 503221 59603 503287 59604
rect 503360 59530 503420 60106
rect 483368 59470 483490 59530
rect 485952 59470 486066 59530
rect 473491 58988 473557 58989
rect 473491 58924 473492 58988
rect 473556 58924 473557 58988
rect 473491 58923 473557 58924
rect 470915 57900 470981 57901
rect 470915 57836 470916 57900
rect 470980 57836 470981 57900
rect 470915 57835 470981 57836
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 43174 474134 58000
rect 475886 57901 475946 59470
rect 478462 59261 478522 59470
rect 478459 59260 478525 59261
rect 478459 59196 478460 59260
rect 478524 59196 478525 59260
rect 478459 59195 478525 59196
rect 475883 57900 475949 57901
rect 475883 57836 475884 57900
rect 475948 57836 475949 57900
rect 475883 57835 475949 57836
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 46894 477854 58000
rect 480670 57901 480730 59470
rect 480667 57900 480733 57901
rect 480667 57836 480668 57900
rect 480732 57836 480733 57900
rect 480667 57835 480733 57836
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 50614 481574 58000
rect 483430 57901 483490 59470
rect 486006 59125 486066 59470
rect 503302 59470 503420 59530
rect 486003 59124 486069 59125
rect 486003 59060 486004 59124
rect 486068 59060 486069 59124
rect 486003 59059 486069 59060
rect 483427 57900 483493 57901
rect 483427 57836 483428 57900
rect 483492 57836 483493 57900
rect 483427 57835 483493 57836
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 57454 488414 58000
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 25174 492134 58000
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 28894 495854 58000
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 32614 499574 58000
rect 503302 57901 503362 59470
rect 503299 57900 503365 57901
rect 503299 57836 503300 57900
rect 503364 57836 503365 57900
rect 503299 57835 503365 57836
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 39454 506414 58000
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 43174 510134 58000
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 46894 513854 58000
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 50614 517574 58000
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 79610 633218 79846 633454
rect 79610 632898 79846 633134
rect 110330 633218 110566 633454
rect 110330 632898 110566 633134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 64250 615218 64486 615454
rect 64250 614898 64486 615134
rect 94970 615218 95206 615454
rect 94970 614898 95206 615134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 79610 597218 79846 597454
rect 79610 596898 79846 597134
rect 110330 597218 110566 597454
rect 110330 596898 110566 597134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 73826 562158 74062 562394
rect 74146 562158 74382 562394
rect 73826 561838 74062 562074
rect 74146 561838 74382 562074
rect 77546 565878 77782 566114
rect 77866 565878 78102 566114
rect 77546 565558 77782 565794
rect 77866 565558 78102 565794
rect 81266 567718 81502 567954
rect 81586 567718 81822 567954
rect 81266 567398 81502 567634
rect 81586 567398 81822 567634
rect 84986 571438 85222 571674
rect 85306 571438 85542 571674
rect 84986 571118 85222 571354
rect 85306 571118 85542 571354
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 109826 562158 110062 562394
rect 110146 562158 110382 562394
rect 109826 561838 110062 562074
rect 110146 561838 110382 562074
rect 113546 565878 113782 566114
rect 113866 565878 114102 566114
rect 113546 565558 113782 565794
rect 113866 565558 114102 565794
rect 117266 567718 117502 567954
rect 117586 567718 117822 567954
rect 117266 567398 117502 567634
rect 117586 567398 117822 567634
rect 120986 571438 121222 571674
rect 121306 571438 121542 571674
rect 120986 571118 121222 571354
rect 121306 571118 121542 571354
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 169610 633218 169846 633454
rect 169610 632898 169846 633134
rect 200330 633218 200566 633454
rect 200330 632898 200566 633134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 154250 615218 154486 615454
rect 154250 614898 154486 615134
rect 184970 615218 185206 615454
rect 184970 614898 185206 615134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 169610 597218 169846 597454
rect 169610 596898 169846 597134
rect 200330 597218 200566 597454
rect 200330 596898 200566 597134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 145826 562158 146062 562394
rect 146146 562158 146382 562394
rect 145826 561838 146062 562074
rect 146146 561838 146382 562074
rect 149546 565878 149782 566114
rect 149866 565878 150102 566114
rect 149546 565558 149782 565794
rect 149866 565558 150102 565794
rect 153266 567718 153502 567954
rect 153586 567718 153822 567954
rect 153266 567398 153502 567634
rect 153586 567398 153822 567634
rect 156986 571438 157222 571674
rect 157306 571438 157542 571674
rect 156986 571118 157222 571354
rect 157306 571118 157542 571354
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 181826 562158 182062 562394
rect 182146 562158 182382 562394
rect 181826 561838 182062 562074
rect 182146 561838 182382 562074
rect 185546 565878 185782 566114
rect 185866 565878 186102 566114
rect 185546 565558 185782 565794
rect 185866 565558 186102 565794
rect 189266 567718 189502 567954
rect 189586 567718 189822 567954
rect 189266 567398 189502 567634
rect 189586 567398 189822 567634
rect 192986 571438 193222 571674
rect 193306 571438 193542 571674
rect 192986 571118 193222 571354
rect 193306 571118 193542 571354
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 217826 562158 218062 562394
rect 218146 562158 218382 562394
rect 217826 561838 218062 562074
rect 218146 561838 218382 562074
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 565878 221782 566114
rect 221866 565878 222102 566114
rect 221546 565558 221782 565794
rect 221866 565558 222102 565794
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 567718 225502 567954
rect 225586 567718 225822 567954
rect 225266 567398 225502 567634
rect 225586 567398 225822 567634
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 571438 229222 571674
rect 229306 571438 229542 571674
rect 228986 571118 229222 571354
rect 229306 571118 229542 571354
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 259610 633218 259846 633454
rect 259610 632898 259846 633134
rect 290330 633218 290566 633454
rect 290330 632898 290566 633134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 244250 615218 244486 615454
rect 244250 614898 244486 615134
rect 274970 615218 275206 615454
rect 274970 614898 275206 615134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 259610 597218 259846 597454
rect 259610 596898 259846 597134
rect 290330 597218 290566 597454
rect 290330 596898 290566 597134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 253826 562158 254062 562394
rect 254146 562158 254382 562394
rect 253826 561838 254062 562074
rect 254146 561838 254382 562074
rect 257546 565878 257782 566114
rect 257866 565878 258102 566114
rect 257546 565558 257782 565794
rect 257866 565558 258102 565794
rect 261266 567718 261502 567954
rect 261586 567718 261822 567954
rect 261266 567398 261502 567634
rect 261586 567398 261822 567634
rect 264986 571438 265222 571674
rect 265306 571438 265542 571674
rect 264986 571118 265222 571354
rect 265306 571118 265542 571354
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 289826 562158 290062 562394
rect 290146 562158 290382 562394
rect 289826 561838 290062 562074
rect 290146 561838 290382 562074
rect 293546 565878 293782 566114
rect 293866 565878 294102 566114
rect 293546 565558 293782 565794
rect 293866 565558 294102 565794
rect 297266 567718 297502 567954
rect 297586 567718 297822 567954
rect 297266 567398 297502 567634
rect 297586 567398 297822 567634
rect 300986 571438 301222 571674
rect 301306 571438 301542 571674
rect 300986 571118 301222 571354
rect 301306 571118 301542 571354
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 64250 543218 64486 543454
rect 64250 542898 64486 543134
rect 94970 543218 95206 543454
rect 94970 542898 95206 543134
rect 125690 543218 125926 543454
rect 125690 542898 125926 543134
rect 156410 543218 156646 543454
rect 156410 542898 156646 543134
rect 187130 543218 187366 543454
rect 187130 542898 187366 543134
rect 217850 543218 218086 543454
rect 217850 542898 218086 543134
rect 248570 543218 248806 543454
rect 248570 542898 248806 543134
rect 279290 543218 279526 543454
rect 279290 542898 279526 543134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 79610 525218 79846 525454
rect 79610 524898 79846 525134
rect 110330 525218 110566 525454
rect 110330 524898 110566 525134
rect 141050 525218 141286 525454
rect 141050 524898 141286 525134
rect 171770 525218 172006 525454
rect 171770 524898 172006 525134
rect 202490 525218 202726 525454
rect 202490 524898 202726 525134
rect 233210 525218 233446 525454
rect 233210 524898 233446 525134
rect 263930 525218 264166 525454
rect 263930 524898 264166 525134
rect 294650 525218 294886 525454
rect 294650 524898 294886 525134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 64250 507218 64486 507454
rect 64250 506898 64486 507134
rect 94970 507218 95206 507454
rect 94970 506898 95206 507134
rect 125690 507218 125926 507454
rect 125690 506898 125926 507134
rect 156410 507218 156646 507454
rect 156410 506898 156646 507134
rect 187130 507218 187366 507454
rect 187130 506898 187366 507134
rect 217850 507218 218086 507454
rect 217850 506898 218086 507134
rect 248570 507218 248806 507454
rect 248570 506898 248806 507134
rect 279290 507218 279526 507454
rect 279290 506898 279526 507134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 59546 475878 59782 476114
rect 59866 475878 60102 476114
rect 59546 475558 59782 475794
rect 59866 475558 60102 475794
rect 63266 479598 63502 479834
rect 63586 479598 63822 479834
rect 63266 479278 63502 479514
rect 63586 479278 63822 479514
rect 66986 481438 67222 481674
rect 67306 481438 67542 481674
rect 66986 481118 67222 481354
rect 67306 481118 67542 481354
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 95546 475878 95782 476114
rect 95866 475878 96102 476114
rect 95546 475558 95782 475794
rect 95866 475558 96102 475794
rect 99266 479598 99502 479834
rect 99586 479598 99822 479834
rect 99266 479278 99502 479514
rect 99586 479278 99822 479514
rect 102986 481438 103222 481674
rect 103306 481438 103542 481674
rect 102986 481118 103222 481354
rect 103306 481118 103542 481354
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 131546 475878 131782 476114
rect 131866 475878 132102 476114
rect 131546 475558 131782 475794
rect 131866 475558 132102 475794
rect 135266 479598 135502 479834
rect 135586 479598 135822 479834
rect 135266 479278 135502 479514
rect 135586 479278 135822 479514
rect 138986 481438 139222 481674
rect 139306 481438 139542 481674
rect 138986 481118 139222 481354
rect 139306 481118 139542 481354
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 167546 475878 167782 476114
rect 167866 475878 168102 476114
rect 167546 475558 167782 475794
rect 167866 475558 168102 475794
rect 171266 479598 171502 479834
rect 171586 479598 171822 479834
rect 171266 479278 171502 479514
rect 171586 479278 171822 479514
rect 174986 481438 175222 481674
rect 175306 481438 175542 481674
rect 174986 481118 175222 481354
rect 175306 481118 175542 481354
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 60328 453218 60564 453454
rect 60328 452898 60564 453134
rect 196056 453218 196292 453454
rect 196056 452898 196292 453134
rect 61008 435218 61244 435454
rect 61008 434898 61244 435134
rect 195376 435218 195612 435454
rect 195376 434898 195612 435134
rect 60328 417218 60564 417454
rect 60328 416898 60564 417134
rect 196056 417218 196292 417454
rect 196056 416898 196292 417134
rect 61008 399218 61244 399454
rect 61008 398898 61244 399134
rect 195376 399218 195612 399454
rect 195376 398898 195612 399134
rect 59546 367878 59782 368114
rect 59866 367878 60102 368114
rect 59546 367558 59782 367794
rect 59866 367558 60102 367794
rect 63266 369718 63502 369954
rect 63586 369718 63822 369954
rect 63266 369398 63502 369634
rect 63586 369398 63822 369634
rect 66986 373438 67222 373674
rect 67306 373438 67542 373674
rect 66986 373118 67222 373354
rect 67306 373118 67542 373354
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 91826 364158 92062 364394
rect 92146 364158 92382 364394
rect 91826 363838 92062 364074
rect 92146 363838 92382 364074
rect 95546 367878 95782 368114
rect 95866 367878 96102 368114
rect 95546 367558 95782 367794
rect 95866 367558 96102 367794
rect 99266 369718 99502 369954
rect 99586 369718 99822 369954
rect 99266 369398 99502 369634
rect 99586 369398 99822 369634
rect 102986 373438 103222 373674
rect 103306 373438 103542 373674
rect 102986 373118 103222 373354
rect 103306 373118 103542 373354
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 127826 364158 128062 364394
rect 128146 364158 128382 364394
rect 127826 363838 128062 364074
rect 128146 363838 128382 364074
rect 131546 367878 131782 368114
rect 131866 367878 132102 368114
rect 131546 367558 131782 367794
rect 131866 367558 132102 367794
rect 135266 369718 135502 369954
rect 135586 369718 135822 369954
rect 135266 369398 135502 369634
rect 135586 369398 135822 369634
rect 138986 373438 139222 373674
rect 139306 373438 139542 373674
rect 138986 373118 139222 373354
rect 139306 373118 139542 373354
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 163826 364158 164062 364394
rect 164146 364158 164382 364394
rect 163826 363838 164062 364074
rect 164146 363838 164382 364074
rect 167546 367878 167782 368114
rect 167866 367878 168102 368114
rect 167546 367558 167782 367794
rect 167866 367558 168102 367794
rect 171266 369718 171502 369954
rect 171586 369718 171822 369954
rect 171266 369398 171502 369634
rect 171586 369398 171822 369634
rect 174986 373438 175222 373674
rect 175306 373438 175542 373674
rect 174986 373118 175222 373354
rect 175306 373118 175542 373354
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 60328 345218 60564 345454
rect 60328 344898 60564 345134
rect 196056 345218 196292 345454
rect 196056 344898 196292 345134
rect 61008 327218 61244 327454
rect 61008 326898 61244 327134
rect 195376 327218 195612 327454
rect 195376 326898 195612 327134
rect 60328 309218 60564 309454
rect 60328 308898 60564 309134
rect 196056 309218 196292 309454
rect 196056 308898 196292 309134
rect 61008 291218 61244 291454
rect 61008 290898 61244 291134
rect 195376 291218 195612 291454
rect 195376 290898 195612 291134
rect 59546 259878 59782 260114
rect 59866 259878 60102 260114
rect 59546 259558 59782 259794
rect 59866 259558 60102 259794
rect 63266 261718 63502 261954
rect 63586 261718 63822 261954
rect 63266 261398 63502 261634
rect 63586 261398 63822 261634
rect 66986 265438 67222 265674
rect 67306 265438 67542 265674
rect 66986 265118 67222 265354
rect 67306 265118 67542 265354
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 91826 256158 92062 256394
rect 92146 256158 92382 256394
rect 91826 255838 92062 256074
rect 92146 255838 92382 256074
rect 95546 259878 95782 260114
rect 95866 259878 96102 260114
rect 95546 259558 95782 259794
rect 95866 259558 96102 259794
rect 99266 261718 99502 261954
rect 99586 261718 99822 261954
rect 99266 261398 99502 261634
rect 99586 261398 99822 261634
rect 102986 265438 103222 265674
rect 103306 265438 103542 265674
rect 102986 265118 103222 265354
rect 103306 265118 103542 265354
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 127826 256158 128062 256394
rect 128146 256158 128382 256394
rect 127826 255838 128062 256074
rect 128146 255838 128382 256074
rect 131546 259878 131782 260114
rect 131866 259878 132102 260114
rect 131546 259558 131782 259794
rect 131866 259558 132102 259794
rect 135266 261718 135502 261954
rect 135586 261718 135822 261954
rect 135266 261398 135502 261634
rect 135586 261398 135822 261634
rect 138986 265438 139222 265674
rect 139306 265438 139542 265674
rect 138986 265118 139222 265354
rect 139306 265118 139542 265354
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 163826 256158 164062 256394
rect 164146 256158 164382 256394
rect 163826 255838 164062 256074
rect 164146 255838 164382 256074
rect 167546 259878 167782 260114
rect 167866 259878 168102 260114
rect 167546 259558 167782 259794
rect 167866 259558 168102 259794
rect 171266 261718 171502 261954
rect 171586 261718 171822 261954
rect 171266 261398 171502 261634
rect 171586 261398 171822 261634
rect 174986 265438 175222 265674
rect 175306 265438 175542 265674
rect 174986 265118 175222 265354
rect 175306 265118 175542 265354
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 60328 237218 60564 237454
rect 60328 236898 60564 237134
rect 196056 237218 196292 237454
rect 196056 236898 196292 237134
rect 61008 219218 61244 219454
rect 61008 218898 61244 219134
rect 195376 219218 195612 219454
rect 195376 218898 195612 219134
rect 60328 201218 60564 201454
rect 60328 200898 60564 201134
rect 196056 201218 196292 201454
rect 196056 200898 196292 201134
rect 61008 183218 61244 183454
rect 61008 182898 61244 183134
rect 195376 183218 195612 183454
rect 195376 182898 195612 183134
rect 59546 151878 59782 152114
rect 59866 151878 60102 152114
rect 59546 151558 59782 151794
rect 59866 151558 60102 151794
rect 63266 155598 63502 155834
rect 63586 155598 63822 155834
rect 63266 155278 63502 155514
rect 63586 155278 63822 155514
rect 66986 157438 67222 157674
rect 67306 157438 67542 157674
rect 66986 157118 67222 157354
rect 67306 157118 67542 157354
rect 73826 147218 74062 147454
rect 74146 147218 74382 147454
rect 73826 146898 74062 147134
rect 74146 146898 74382 147134
rect 77546 150938 77782 151174
rect 77866 150938 78102 151174
rect 77546 150618 77782 150854
rect 77866 150618 78102 150854
rect 81266 154658 81502 154894
rect 81586 154658 81822 154894
rect 81266 154338 81502 154574
rect 81586 154338 81822 154574
rect 84986 158378 85222 158614
rect 85306 158378 85542 158614
rect 84986 158058 85222 158294
rect 85306 158058 85542 158294
rect 91826 148158 92062 148394
rect 92146 148158 92382 148394
rect 91826 147838 92062 148074
rect 92146 147838 92382 148074
rect 95546 151878 95782 152114
rect 95866 151878 96102 152114
rect 95546 151558 95782 151794
rect 95866 151558 96102 151794
rect 99266 155598 99502 155834
rect 99586 155598 99822 155834
rect 99266 155278 99502 155514
rect 99586 155278 99822 155514
rect 102986 157438 103222 157674
rect 103306 157438 103542 157674
rect 102986 157118 103222 157354
rect 103306 157118 103542 157354
rect 109826 147218 110062 147454
rect 110146 147218 110382 147454
rect 109826 146898 110062 147134
rect 110146 146898 110382 147134
rect 113546 150938 113782 151174
rect 113866 150938 114102 151174
rect 113546 150618 113782 150854
rect 113866 150618 114102 150854
rect 117266 154658 117502 154894
rect 117586 154658 117822 154894
rect 117266 154338 117502 154574
rect 117586 154338 117822 154574
rect 120986 158378 121222 158614
rect 121306 158378 121542 158614
rect 120986 158058 121222 158294
rect 121306 158058 121542 158294
rect 127826 148158 128062 148394
rect 128146 148158 128382 148394
rect 127826 147838 128062 148074
rect 128146 147838 128382 148074
rect 131546 151878 131782 152114
rect 131866 151878 132102 152114
rect 131546 151558 131782 151794
rect 131866 151558 132102 151794
rect 135266 155598 135502 155834
rect 135586 155598 135822 155834
rect 135266 155278 135502 155514
rect 135586 155278 135822 155514
rect 138986 157438 139222 157674
rect 139306 157438 139542 157674
rect 138986 157118 139222 157354
rect 139306 157118 139542 157354
rect 145826 147218 146062 147454
rect 146146 147218 146382 147454
rect 145826 146898 146062 147134
rect 146146 146898 146382 147134
rect 149546 150938 149782 151174
rect 149866 150938 150102 151174
rect 149546 150618 149782 150854
rect 149866 150618 150102 150854
rect 153266 154658 153502 154894
rect 153586 154658 153822 154894
rect 153266 154338 153502 154574
rect 153586 154338 153822 154574
rect 156986 158378 157222 158614
rect 157306 158378 157542 158614
rect 156986 158058 157222 158294
rect 157306 158058 157542 158294
rect 163826 148158 164062 148394
rect 164146 148158 164382 148394
rect 163826 147838 164062 148074
rect 164146 147838 164382 148074
rect 167546 151878 167782 152114
rect 167866 151878 168102 152114
rect 167546 151558 167782 151794
rect 167866 151558 168102 151794
rect 171266 155598 171502 155834
rect 171586 155598 171822 155834
rect 171266 155278 171502 155514
rect 171586 155278 171822 155514
rect 174986 157438 175222 157674
rect 175306 157438 175542 157674
rect 174986 157118 175222 157354
rect 175306 157118 175542 157354
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 60328 129218 60564 129454
rect 60328 128898 60564 129134
rect 196056 129218 196292 129454
rect 196056 128898 196292 129134
rect 61008 111218 61244 111454
rect 61008 110898 61244 111134
rect 195376 111218 195612 111454
rect 195376 110898 195612 111134
rect 60328 93218 60564 93454
rect 60328 92898 60564 93134
rect 196056 93218 196292 93454
rect 196056 92898 196292 93134
rect 61008 75218 61244 75454
rect 61008 74898 61244 75134
rect 195376 75218 195612 75454
rect 195376 74898 195612 75134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 364158 200062 364394
rect 200146 364158 200382 364394
rect 199826 363838 200062 364074
rect 200146 363838 200382 364074
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 256158 200062 256394
rect 200146 256158 200382 256394
rect 199826 255838 200062 256074
rect 200146 255838 200382 256074
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 148158 200062 148394
rect 200146 148158 200382 148394
rect 199826 147838 200062 148074
rect 200146 147838 200382 148074
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 203546 475878 203782 476114
rect 203866 475878 204102 476114
rect 203546 475558 203782 475794
rect 203866 475558 204102 475794
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 367878 203782 368114
rect 203866 367878 204102 368114
rect 203546 367558 203782 367794
rect 203866 367558 204102 367794
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 203546 276938 203782 277174
rect 203866 276938 204102 277174
rect 203546 276618 203782 276854
rect 203866 276618 204102 276854
rect 203546 259878 203782 260114
rect 203866 259878 204102 260114
rect 203546 259558 203782 259794
rect 203866 259558 204102 259794
rect 203546 240938 203782 241174
rect 203866 240938 204102 241174
rect 203546 240618 203782 240854
rect 203866 240618 204102 240854
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 151878 203782 152114
rect 203866 151878 204102 152114
rect 203546 151558 203782 151794
rect 203866 151558 204102 151794
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 207266 479598 207502 479834
rect 207586 479598 207822 479834
rect 207266 479278 207502 479514
rect 207586 479278 207822 479514
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 369718 207502 369954
rect 207586 369718 207822 369954
rect 207266 369398 207502 369634
rect 207586 369398 207822 369634
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 207266 280658 207502 280894
rect 207586 280658 207822 280894
rect 207266 280338 207502 280574
rect 207586 280338 207822 280574
rect 207266 261718 207502 261954
rect 207586 261718 207822 261954
rect 207266 261398 207502 261634
rect 207586 261398 207822 261634
rect 207266 244658 207502 244894
rect 207586 244658 207822 244894
rect 207266 244338 207502 244574
rect 207586 244338 207822 244574
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 155598 207502 155834
rect 207586 155598 207822 155834
rect 207266 155278 207502 155514
rect 207586 155278 207822 155514
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 210986 481438 211222 481674
rect 211306 481438 211542 481674
rect 210986 481118 211222 481354
rect 211306 481118 211542 481354
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 373438 211222 373674
rect 211306 373438 211542 373674
rect 210986 373118 211222 373354
rect 211306 373118 211542 373354
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 210986 284378 211222 284614
rect 211306 284378 211542 284614
rect 210986 284058 211222 284294
rect 211306 284058 211542 284294
rect 210986 265438 211222 265674
rect 211306 265438 211542 265674
rect 210986 265118 211222 265354
rect 211306 265118 211542 265354
rect 210986 248378 211222 248614
rect 211306 248378 211542 248614
rect 210986 248058 211222 248294
rect 211306 248058 211542 248294
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 210986 157438 211222 157674
rect 211306 157438 211542 157674
rect 210986 157118 211222 157354
rect 211306 157118 211542 157354
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 217826 147218 218062 147454
rect 218146 147218 218382 147454
rect 217826 146898 218062 147134
rect 218146 146898 218382 147134
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 239546 475878 239782 476114
rect 239866 475878 240102 476114
rect 239546 475558 239782 475794
rect 239866 475558 240102 475794
rect 243266 479598 243502 479834
rect 243586 479598 243822 479834
rect 243266 479278 243502 479514
rect 243586 479278 243822 479514
rect 246986 481438 247222 481674
rect 247306 481438 247542 481674
rect 246986 481118 247222 481354
rect 247306 481118 247542 481354
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 275546 475878 275782 476114
rect 275866 475878 276102 476114
rect 275546 475558 275782 475794
rect 275866 475558 276102 475794
rect 279266 479598 279502 479834
rect 279586 479598 279822 479834
rect 279266 479278 279502 479514
rect 279586 479278 279822 479514
rect 282986 481438 283222 481674
rect 283306 481438 283542 481674
rect 282986 481118 283222 481354
rect 283306 481118 283542 481354
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 344610 633218 344846 633454
rect 344610 632898 344846 633134
rect 375330 633218 375566 633454
rect 375330 632898 375566 633134
rect 406050 633218 406286 633454
rect 406050 632898 406286 633134
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 329250 615218 329486 615454
rect 329250 614898 329486 615134
rect 359970 615218 360206 615454
rect 359970 614898 360206 615134
rect 390690 615218 390926 615454
rect 390690 614898 390926 615134
rect 421410 615218 421646 615454
rect 421410 614898 421646 615134
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 344610 597218 344846 597454
rect 344610 596898 344846 597134
rect 375330 597218 375566 597454
rect 375330 596898 375566 597134
rect 406050 597218 406286 597454
rect 406050 596898 406286 597134
rect 329250 579218 329486 579454
rect 329250 578898 329486 579134
rect 359970 579218 360206 579454
rect 359970 578898 360206 579134
rect 390690 579218 390926 579454
rect 390690 578898 390926 579134
rect 421410 579218 421646 579454
rect 421410 578898 421646 579134
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 344610 561218 344846 561454
rect 344610 560898 344846 561134
rect 375330 561218 375566 561454
rect 375330 560898 375566 561134
rect 406050 561218 406286 561454
rect 406050 560898 406286 561134
rect 329250 543218 329486 543454
rect 329250 542898 329486 543134
rect 359970 543218 360206 543454
rect 359970 542898 360206 543134
rect 390690 543218 390926 543454
rect 390690 542898 390926 543134
rect 421410 543218 421646 543454
rect 421410 542898 421646 543134
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 220328 453218 220564 453454
rect 220328 452898 220564 453134
rect 356056 453218 356292 453454
rect 356056 452898 356292 453134
rect 221008 435218 221244 435454
rect 221008 434898 221244 435134
rect 355376 435218 355612 435454
rect 355376 434898 355612 435134
rect 220328 417218 220564 417454
rect 220328 416898 220564 417134
rect 356056 417218 356292 417454
rect 356056 416898 356292 417134
rect 221008 399218 221244 399454
rect 221008 398898 221244 399134
rect 355376 399218 355612 399454
rect 355376 398898 355612 399134
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 235826 364158 236062 364394
rect 236146 364158 236382 364394
rect 235826 363838 236062 364074
rect 236146 363838 236382 364074
rect 239546 367878 239782 368114
rect 239866 367878 240102 368114
rect 239546 367558 239782 367794
rect 239866 367558 240102 367794
rect 243266 369718 243502 369954
rect 243586 369718 243822 369954
rect 243266 369398 243502 369634
rect 243586 369398 243822 369634
rect 246986 373438 247222 373674
rect 247306 373438 247542 373674
rect 246986 373118 247222 373354
rect 247306 373118 247542 373354
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 271826 364158 272062 364394
rect 272146 364158 272382 364394
rect 271826 363838 272062 364074
rect 272146 363838 272382 364074
rect 275546 367878 275782 368114
rect 275866 367878 276102 368114
rect 275546 367558 275782 367794
rect 275866 367558 276102 367794
rect 279266 369718 279502 369954
rect 279586 369718 279822 369954
rect 279266 369398 279502 369634
rect 279586 369398 279822 369634
rect 282986 373438 283222 373674
rect 283306 373438 283542 373674
rect 282986 373118 283222 373354
rect 283306 373118 283542 373354
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 307826 364158 308062 364394
rect 308146 364158 308382 364394
rect 307826 363838 308062 364074
rect 308146 363838 308382 364074
rect 311546 367878 311782 368114
rect 311866 367878 312102 368114
rect 311546 367558 311782 367794
rect 311866 367558 312102 367794
rect 315266 369718 315502 369954
rect 315586 369718 315822 369954
rect 315266 369398 315502 369634
rect 315586 369398 315822 369634
rect 318986 373438 319222 373674
rect 319306 373438 319542 373674
rect 318986 373118 319222 373354
rect 319306 373118 319542 373354
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 343826 364158 344062 364394
rect 344146 364158 344382 364394
rect 343826 363838 344062 364074
rect 344146 363838 344382 364074
rect 347546 367878 347782 368114
rect 347866 367878 348102 368114
rect 347546 367558 347782 367794
rect 347866 367558 348102 367794
rect 351266 369718 351502 369954
rect 351586 369718 351822 369954
rect 351266 369398 351502 369634
rect 351586 369398 351822 369634
rect 354986 373438 355222 373674
rect 355306 373438 355542 373674
rect 354986 373118 355222 373354
rect 355306 373118 355542 373354
rect 220328 345218 220564 345454
rect 220328 344898 220564 345134
rect 356056 345218 356292 345454
rect 356056 344898 356292 345134
rect 221008 327218 221244 327454
rect 221008 326898 221244 327134
rect 355376 327218 355612 327454
rect 355376 326898 355612 327134
rect 220328 309218 220564 309454
rect 220328 308898 220564 309134
rect 356056 309218 356292 309454
rect 356056 308898 356292 309134
rect 221008 291218 221244 291454
rect 221008 290898 221244 291134
rect 355376 291218 355612 291454
rect 355376 290898 355612 291134
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 235826 256158 236062 256394
rect 236146 256158 236382 256394
rect 235826 255838 236062 256074
rect 236146 255838 236382 256074
rect 239546 259878 239782 260114
rect 239866 259878 240102 260114
rect 239546 259558 239782 259794
rect 239866 259558 240102 259794
rect 243266 261718 243502 261954
rect 243586 261718 243822 261954
rect 243266 261398 243502 261634
rect 243586 261398 243822 261634
rect 246986 265438 247222 265674
rect 247306 265438 247542 265674
rect 246986 265118 247222 265354
rect 247306 265118 247542 265354
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 271826 256158 272062 256394
rect 272146 256158 272382 256394
rect 271826 255838 272062 256074
rect 272146 255838 272382 256074
rect 275546 259878 275782 260114
rect 275866 259878 276102 260114
rect 275546 259558 275782 259794
rect 275866 259558 276102 259794
rect 279266 261718 279502 261954
rect 279586 261718 279822 261954
rect 279266 261398 279502 261634
rect 279586 261398 279822 261634
rect 282986 265438 283222 265674
rect 283306 265438 283542 265674
rect 282986 265118 283222 265354
rect 283306 265118 283542 265354
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 307826 256158 308062 256394
rect 308146 256158 308382 256394
rect 307826 255838 308062 256074
rect 308146 255838 308382 256074
rect 311546 259878 311782 260114
rect 311866 259878 312102 260114
rect 311546 259558 311782 259794
rect 311866 259558 312102 259794
rect 315266 261718 315502 261954
rect 315586 261718 315822 261954
rect 315266 261398 315502 261634
rect 315586 261398 315822 261634
rect 318986 265438 319222 265674
rect 319306 265438 319542 265674
rect 318986 265118 319222 265354
rect 319306 265118 319542 265354
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 343826 256158 344062 256394
rect 344146 256158 344382 256394
rect 343826 255838 344062 256074
rect 344146 255838 344382 256074
rect 347546 259878 347782 260114
rect 347866 259878 348102 260114
rect 347546 259558 347782 259794
rect 347866 259558 348102 259794
rect 351266 261718 351502 261954
rect 351586 261718 351822 261954
rect 351266 261398 351502 261634
rect 351586 261398 351822 261634
rect 354986 265438 355222 265674
rect 355306 265438 355542 265674
rect 354986 265118 355222 265354
rect 355306 265118 355542 265354
rect 220328 237218 220564 237454
rect 220328 236898 220564 237134
rect 356056 237218 356292 237454
rect 356056 236898 356292 237134
rect 221008 219218 221244 219454
rect 221008 218898 221244 219134
rect 355376 219218 355612 219454
rect 355376 218898 355612 219134
rect 220328 201218 220564 201454
rect 220328 200898 220564 201134
rect 356056 201218 356292 201454
rect 356056 200898 356292 201134
rect 221008 183218 221244 183454
rect 221008 182898 221244 183134
rect 355376 183218 355612 183454
rect 355376 182898 355612 183134
rect 221546 150938 221782 151174
rect 221866 150938 222102 151174
rect 221546 150618 221782 150854
rect 221866 150618 222102 150854
rect 225266 154658 225502 154894
rect 225586 154658 225822 154894
rect 225266 154338 225502 154574
rect 225586 154338 225822 154574
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 235826 148158 236062 148394
rect 236146 148158 236382 148394
rect 235826 147838 236062 148074
rect 236146 147838 236382 148074
rect 239546 151878 239782 152114
rect 239866 151878 240102 152114
rect 239546 151558 239782 151794
rect 239866 151558 240102 151794
rect 243266 155598 243502 155834
rect 243586 155598 243822 155834
rect 243266 155278 243502 155514
rect 243586 155278 243822 155514
rect 246986 157438 247222 157674
rect 247306 157438 247542 157674
rect 246986 157118 247222 157354
rect 247306 157118 247542 157354
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 271826 148158 272062 148394
rect 272146 148158 272382 148394
rect 271826 147838 272062 148074
rect 272146 147838 272382 148074
rect 275546 151878 275782 152114
rect 275866 151878 276102 152114
rect 275546 151558 275782 151794
rect 275866 151558 276102 151794
rect 279266 155598 279502 155834
rect 279586 155598 279822 155834
rect 279266 155278 279502 155514
rect 279586 155278 279822 155514
rect 282986 157438 283222 157674
rect 283306 157438 283542 157674
rect 282986 157118 283222 157354
rect 283306 157118 283542 157354
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 307826 148158 308062 148394
rect 308146 148158 308382 148394
rect 307826 147838 308062 148074
rect 308146 147838 308382 148074
rect 311546 151878 311782 152114
rect 311866 151878 312102 152114
rect 311546 151558 311782 151794
rect 311866 151558 312102 151794
rect 315266 155598 315502 155834
rect 315586 155598 315822 155834
rect 315266 155278 315502 155514
rect 315586 155278 315822 155514
rect 318986 157438 319222 157674
rect 319306 157438 319542 157674
rect 318986 157118 319222 157354
rect 319306 157118 319542 157354
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 343826 148158 344062 148394
rect 344146 148158 344382 148394
rect 343826 147838 344062 148074
rect 344146 147838 344382 148074
rect 347546 151878 347782 152114
rect 347866 151878 348102 152114
rect 347546 151558 347782 151794
rect 347866 151558 348102 151794
rect 351266 155598 351502 155834
rect 351586 155598 351822 155834
rect 351266 155278 351502 155514
rect 351586 155278 351822 155514
rect 354986 157438 355222 157674
rect 355306 157438 355542 157674
rect 354986 157118 355222 157354
rect 355306 157118 355542 157354
rect 220328 129218 220564 129454
rect 220328 128898 220564 129134
rect 356056 129218 356292 129454
rect 356056 128898 356292 129134
rect 221008 111218 221244 111454
rect 221008 110898 221244 111134
rect 355376 111218 355612 111454
rect 355376 110898 355612 111134
rect 220328 93218 220564 93454
rect 220328 92898 220564 93134
rect 356056 93218 356292 93454
rect 356056 92898 356292 93134
rect 221008 75218 221244 75454
rect 221008 74898 221244 75134
rect 355376 75218 355612 75454
rect 355376 74898 355612 75134
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 464250 615218 464486 615454
rect 464250 614898 464486 615134
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 479610 633218 479846 633454
rect 479610 632898 479846 633134
rect 479610 597218 479846 597454
rect 479610 596898 479846 597134
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 494970 615218 495206 615454
rect 494970 614898 495206 615134
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 380328 453218 380564 453454
rect 380328 452898 380564 453134
rect 516056 453218 516292 453454
rect 516056 452898 516292 453134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 381008 435218 381244 435454
rect 381008 434898 381244 435134
rect 515376 435218 515612 435454
rect 515376 434898 515612 435134
rect 380328 417218 380564 417454
rect 380328 416898 380564 417134
rect 516056 417218 516292 417454
rect 516056 416898 516292 417134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 381008 399218 381244 399454
rect 381008 398898 381244 399134
rect 515376 399218 515612 399454
rect 515376 398898 515612 399134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 379826 364158 380062 364394
rect 380146 364158 380382 364394
rect 379826 363838 380062 364074
rect 380146 363838 380382 364074
rect 383546 367878 383782 368114
rect 383866 367878 384102 368114
rect 383546 367558 383782 367794
rect 383866 367558 384102 367794
rect 387266 369718 387502 369954
rect 387586 369718 387822 369954
rect 387266 369398 387502 369634
rect 387586 369398 387822 369634
rect 390986 373438 391222 373674
rect 391306 373438 391542 373674
rect 390986 373118 391222 373354
rect 391306 373118 391542 373354
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 415826 364158 416062 364394
rect 416146 364158 416382 364394
rect 415826 363838 416062 364074
rect 416146 363838 416382 364074
rect 419546 367878 419782 368114
rect 419866 367878 420102 368114
rect 419546 367558 419782 367794
rect 419866 367558 420102 367794
rect 423266 369718 423502 369954
rect 423586 369718 423822 369954
rect 423266 369398 423502 369634
rect 423586 369398 423822 369634
rect 426986 373438 427222 373674
rect 427306 373438 427542 373674
rect 426986 373118 427222 373354
rect 427306 373118 427542 373354
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 451826 364158 452062 364394
rect 452146 364158 452382 364394
rect 451826 363838 452062 364074
rect 452146 363838 452382 364074
rect 455546 367878 455782 368114
rect 455866 367878 456102 368114
rect 455546 367558 455782 367794
rect 455866 367558 456102 367794
rect 459266 369718 459502 369954
rect 459586 369718 459822 369954
rect 459266 369398 459502 369634
rect 459586 369398 459822 369634
rect 462986 373438 463222 373674
rect 463306 373438 463542 373674
rect 462986 373118 463222 373354
rect 463306 373118 463542 373354
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 487826 364158 488062 364394
rect 488146 364158 488382 364394
rect 487826 363838 488062 364074
rect 488146 363838 488382 364074
rect 491546 367878 491782 368114
rect 491866 367878 492102 368114
rect 491546 367558 491782 367794
rect 491866 367558 492102 367794
rect 495266 369718 495502 369954
rect 495586 369718 495822 369954
rect 495266 369398 495502 369634
rect 495586 369398 495822 369634
rect 498986 373438 499222 373674
rect 499306 373438 499542 373674
rect 498986 373118 499222 373354
rect 499306 373118 499542 373354
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 380328 345218 380564 345454
rect 380328 344898 380564 345134
rect 516056 345218 516292 345454
rect 516056 344898 516292 345134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 381008 327218 381244 327454
rect 381008 326898 381244 327134
rect 515376 327218 515612 327454
rect 515376 326898 515612 327134
rect 380328 309218 380564 309454
rect 380328 308898 380564 309134
rect 516056 309218 516292 309454
rect 516056 308898 516292 309134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 381008 291218 381244 291454
rect 381008 290898 381244 291134
rect 515376 291218 515612 291454
rect 515376 290898 515612 291134
rect 379826 256158 380062 256394
rect 380146 256158 380382 256394
rect 379826 255838 380062 256074
rect 380146 255838 380382 256074
rect 383546 259878 383782 260114
rect 383866 259878 384102 260114
rect 383546 259558 383782 259794
rect 383866 259558 384102 259794
rect 387266 261718 387502 261954
rect 387586 261718 387822 261954
rect 387266 261398 387502 261634
rect 387586 261398 387822 261634
rect 390986 265438 391222 265674
rect 391306 265438 391542 265674
rect 390986 265118 391222 265354
rect 391306 265118 391542 265354
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 415826 256158 416062 256394
rect 416146 256158 416382 256394
rect 415826 255838 416062 256074
rect 416146 255838 416382 256074
rect 419546 259878 419782 260114
rect 419866 259878 420102 260114
rect 419546 259558 419782 259794
rect 419866 259558 420102 259794
rect 423266 261718 423502 261954
rect 423586 261718 423822 261954
rect 423266 261398 423502 261634
rect 423586 261398 423822 261634
rect 426986 265438 427222 265674
rect 427306 265438 427542 265674
rect 426986 265118 427222 265354
rect 427306 265118 427542 265354
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 451826 256158 452062 256394
rect 452146 256158 452382 256394
rect 451826 255838 452062 256074
rect 452146 255838 452382 256074
rect 455546 259878 455782 260114
rect 455866 259878 456102 260114
rect 455546 259558 455782 259794
rect 455866 259558 456102 259794
rect 459266 261718 459502 261954
rect 459586 261718 459822 261954
rect 459266 261398 459502 261634
rect 459586 261398 459822 261634
rect 462986 265438 463222 265674
rect 463306 265438 463542 265674
rect 462986 265118 463222 265354
rect 463306 265118 463542 265354
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 487826 256158 488062 256394
rect 488146 256158 488382 256394
rect 487826 255838 488062 256074
rect 488146 255838 488382 256074
rect 491546 259878 491782 260114
rect 491866 259878 492102 260114
rect 491546 259558 491782 259794
rect 491866 259558 492102 259794
rect 495266 261718 495502 261954
rect 495586 261718 495822 261954
rect 495266 261398 495502 261634
rect 495586 261398 495822 261634
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 498986 265438 499222 265674
rect 499306 265438 499542 265674
rect 498986 265118 499222 265354
rect 499306 265118 499542 265354
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 380328 237218 380564 237454
rect 380328 236898 380564 237134
rect 516056 237218 516292 237454
rect 516056 236898 516292 237134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 381008 219218 381244 219454
rect 381008 218898 381244 219134
rect 515376 219218 515612 219454
rect 515376 218898 515612 219134
rect 380328 201218 380564 201454
rect 380328 200898 380564 201134
rect 516056 201218 516292 201454
rect 516056 200898 516292 201134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 381008 183218 381244 183454
rect 381008 182898 381244 183134
rect 515376 183218 515612 183454
rect 515376 182898 515612 183134
rect 379826 148158 380062 148394
rect 380146 148158 380382 148394
rect 379826 147838 380062 148074
rect 380146 147838 380382 148074
rect 383546 151878 383782 152114
rect 383866 151878 384102 152114
rect 383546 151558 383782 151794
rect 383866 151558 384102 151794
rect 387266 155598 387502 155834
rect 387586 155598 387822 155834
rect 387266 155278 387502 155514
rect 387586 155278 387822 155514
rect 390986 157438 391222 157674
rect 391306 157438 391542 157674
rect 390986 157118 391222 157354
rect 391306 157118 391542 157354
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 415826 148158 416062 148394
rect 416146 148158 416382 148394
rect 415826 147838 416062 148074
rect 416146 147838 416382 148074
rect 419546 151878 419782 152114
rect 419866 151878 420102 152114
rect 419546 151558 419782 151794
rect 419866 151558 420102 151794
rect 423266 155598 423502 155834
rect 423586 155598 423822 155834
rect 423266 155278 423502 155514
rect 423586 155278 423822 155514
rect 426986 157438 427222 157674
rect 427306 157438 427542 157674
rect 426986 157118 427222 157354
rect 427306 157118 427542 157354
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 451826 148158 452062 148394
rect 452146 148158 452382 148394
rect 451826 147838 452062 148074
rect 452146 147838 452382 148074
rect 455546 151878 455782 152114
rect 455866 151878 456102 152114
rect 455546 151558 455782 151794
rect 455866 151558 456102 151794
rect 459266 155598 459502 155834
rect 459586 155598 459822 155834
rect 459266 155278 459502 155514
rect 459586 155278 459822 155514
rect 462986 157438 463222 157674
rect 463306 157438 463542 157674
rect 462986 157118 463222 157354
rect 463306 157118 463542 157354
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 487826 148158 488062 148394
rect 488146 148158 488382 148394
rect 487826 147838 488062 148074
rect 488146 147838 488382 148074
rect 491546 151878 491782 152114
rect 491866 151878 492102 152114
rect 491546 151558 491782 151794
rect 491866 151558 492102 151794
rect 495266 155598 495502 155834
rect 495586 155598 495822 155834
rect 495266 155278 495502 155514
rect 495586 155278 495822 155514
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 498986 157438 499222 157674
rect 499306 157438 499542 157674
rect 498986 157118 499222 157354
rect 499306 157118 499542 157354
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 380328 129218 380564 129454
rect 380328 128898 380564 129134
rect 516056 129218 516292 129454
rect 516056 128898 516292 129134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 381008 111218 381244 111454
rect 381008 110898 381244 111134
rect 515376 111218 515612 111454
rect 515376 110898 515612 111134
rect 380328 93218 380564 93454
rect 380328 92898 380564 93134
rect 516056 93218 516292 93454
rect 516056 92898 516292 93134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 381008 75218 381244 75454
rect 381008 74898 381244 75134
rect 515376 75218 515612 75454
rect 515376 74898 515612 75134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 79610 633454
rect 79846 633218 110330 633454
rect 110566 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 169610 633454
rect 169846 633218 200330 633454
rect 200566 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 259610 633454
rect 259846 633218 290330 633454
rect 290566 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 344610 633454
rect 344846 633218 375330 633454
rect 375566 633218 406050 633454
rect 406286 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 479610 633454
rect 479846 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 79610 633134
rect 79846 632898 110330 633134
rect 110566 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 169610 633134
rect 169846 632898 200330 633134
rect 200566 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 259610 633134
rect 259846 632898 290330 633134
rect 290566 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 344610 633134
rect 344846 632898 375330 633134
rect 375566 632898 406050 633134
rect 406286 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 479610 633134
rect 479846 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 64250 615454
rect 64486 615218 94970 615454
rect 95206 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 154250 615454
rect 154486 615218 184970 615454
rect 185206 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 244250 615454
rect 244486 615218 274970 615454
rect 275206 615218 329250 615454
rect 329486 615218 359970 615454
rect 360206 615218 390690 615454
rect 390926 615218 421410 615454
rect 421646 615218 464250 615454
rect 464486 615218 494970 615454
rect 495206 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 64250 615134
rect 64486 614898 94970 615134
rect 95206 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 154250 615134
rect 154486 614898 184970 615134
rect 185206 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 244250 615134
rect 244486 614898 274970 615134
rect 275206 614898 329250 615134
rect 329486 614898 359970 615134
rect 360206 614898 390690 615134
rect 390926 614898 421410 615134
rect 421646 614898 464250 615134
rect 464486 614898 494970 615134
rect 495206 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 79610 597454
rect 79846 597218 110330 597454
rect 110566 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 169610 597454
rect 169846 597218 200330 597454
rect 200566 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 259610 597454
rect 259846 597218 290330 597454
rect 290566 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 344610 597454
rect 344846 597218 375330 597454
rect 375566 597218 406050 597454
rect 406286 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 479610 597454
rect 479846 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 79610 597134
rect 79846 596898 110330 597134
rect 110566 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 169610 597134
rect 169846 596898 200330 597134
rect 200566 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 259610 597134
rect 259846 596898 290330 597134
rect 290566 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 344610 597134
rect 344846 596898 375330 597134
rect 375566 596898 406050 597134
rect 406286 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 479610 597134
rect 479846 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 329250 579454
rect 329486 579218 359970 579454
rect 360206 579218 390690 579454
rect 390926 579218 421410 579454
rect 421646 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 329250 579134
rect 329486 578898 359970 579134
rect 360206 578898 390690 579134
rect 390926 578898 421410 579134
rect 421646 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect 84954 571674 301574 571706
rect 84954 571438 84986 571674
rect 85222 571438 85306 571674
rect 85542 571438 120986 571674
rect 121222 571438 121306 571674
rect 121542 571438 156986 571674
rect 157222 571438 157306 571674
rect 157542 571438 192986 571674
rect 193222 571438 193306 571674
rect 193542 571438 228986 571674
rect 229222 571438 229306 571674
rect 229542 571438 264986 571674
rect 265222 571438 265306 571674
rect 265542 571438 300986 571674
rect 301222 571438 301306 571674
rect 301542 571438 301574 571674
rect 84954 571354 301574 571438
rect 84954 571118 84986 571354
rect 85222 571118 85306 571354
rect 85542 571118 120986 571354
rect 121222 571118 121306 571354
rect 121542 571118 156986 571354
rect 157222 571118 157306 571354
rect 157542 571118 192986 571354
rect 193222 571118 193306 571354
rect 193542 571118 228986 571354
rect 229222 571118 229306 571354
rect 229542 571118 264986 571354
rect 265222 571118 265306 571354
rect 265542 571118 300986 571354
rect 301222 571118 301306 571354
rect 301542 571118 301574 571354
rect 84954 571086 301574 571118
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect 81234 567954 297854 567986
rect 81234 567718 81266 567954
rect 81502 567718 81586 567954
rect 81822 567718 117266 567954
rect 117502 567718 117586 567954
rect 117822 567718 153266 567954
rect 153502 567718 153586 567954
rect 153822 567718 189266 567954
rect 189502 567718 189586 567954
rect 189822 567718 225266 567954
rect 225502 567718 225586 567954
rect 225822 567718 261266 567954
rect 261502 567718 261586 567954
rect 261822 567718 297266 567954
rect 297502 567718 297586 567954
rect 297822 567718 297854 567954
rect 81234 567634 297854 567718
rect 81234 567398 81266 567634
rect 81502 567398 81586 567634
rect 81822 567398 117266 567634
rect 117502 567398 117586 567634
rect 117822 567398 153266 567634
rect 153502 567398 153586 567634
rect 153822 567398 189266 567634
rect 189502 567398 189586 567634
rect 189822 567398 225266 567634
rect 225502 567398 225586 567634
rect 225822 567398 261266 567634
rect 261502 567398 261586 567634
rect 261822 567398 297266 567634
rect 297502 567398 297586 567634
rect 297822 567398 297854 567634
rect 81234 567366 297854 567398
rect 77514 566114 294134 566146
rect 77514 565878 77546 566114
rect 77782 565878 77866 566114
rect 78102 565878 113546 566114
rect 113782 565878 113866 566114
rect 114102 565878 149546 566114
rect 149782 565878 149866 566114
rect 150102 565878 185546 566114
rect 185782 565878 185866 566114
rect 186102 565878 221546 566114
rect 221782 565878 221866 566114
rect 222102 565878 257546 566114
rect 257782 565878 257866 566114
rect 258102 565878 293546 566114
rect 293782 565878 293866 566114
rect 294102 565878 294134 566114
rect 77514 565794 294134 565878
rect 77514 565558 77546 565794
rect 77782 565558 77866 565794
rect 78102 565558 113546 565794
rect 113782 565558 113866 565794
rect 114102 565558 149546 565794
rect 149782 565558 149866 565794
rect 150102 565558 185546 565794
rect 185782 565558 185866 565794
rect 186102 565558 221546 565794
rect 221782 565558 221866 565794
rect 222102 565558 257546 565794
rect 257782 565558 257866 565794
rect 258102 565558 293546 565794
rect 293782 565558 293866 565794
rect 294102 565558 294134 565794
rect 77514 565526 294134 565558
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect 73794 562394 290414 562426
rect 73794 562158 73826 562394
rect 74062 562158 74146 562394
rect 74382 562158 109826 562394
rect 110062 562158 110146 562394
rect 110382 562158 145826 562394
rect 146062 562158 146146 562394
rect 146382 562158 181826 562394
rect 182062 562158 182146 562394
rect 182382 562158 217826 562394
rect 218062 562158 218146 562394
rect 218382 562158 253826 562394
rect 254062 562158 254146 562394
rect 254382 562158 289826 562394
rect 290062 562158 290146 562394
rect 290382 562158 290414 562394
rect 73794 562074 290414 562158
rect 73794 561838 73826 562074
rect 74062 561838 74146 562074
rect 74382 561838 109826 562074
rect 110062 561838 110146 562074
rect 110382 561838 145826 562074
rect 146062 561838 146146 562074
rect 146382 561838 181826 562074
rect 182062 561838 182146 562074
rect 182382 561838 217826 562074
rect 218062 561838 218146 562074
rect 218382 561838 253826 562074
rect 254062 561838 254146 562074
rect 254382 561838 289826 562074
rect 290062 561838 290146 562074
rect 290382 561838 290414 562074
rect 73794 561806 290414 561838
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 344610 561454
rect 344846 561218 375330 561454
rect 375566 561218 406050 561454
rect 406286 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 344610 561134
rect 344846 560898 375330 561134
rect 375566 560898 406050 561134
rect 406286 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 64250 543454
rect 64486 543218 94970 543454
rect 95206 543218 125690 543454
rect 125926 543218 156410 543454
rect 156646 543218 187130 543454
rect 187366 543218 217850 543454
rect 218086 543218 248570 543454
rect 248806 543218 279290 543454
rect 279526 543218 329250 543454
rect 329486 543218 359970 543454
rect 360206 543218 390690 543454
rect 390926 543218 421410 543454
rect 421646 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 64250 543134
rect 64486 542898 94970 543134
rect 95206 542898 125690 543134
rect 125926 542898 156410 543134
rect 156646 542898 187130 543134
rect 187366 542898 217850 543134
rect 218086 542898 248570 543134
rect 248806 542898 279290 543134
rect 279526 542898 329250 543134
rect 329486 542898 359970 543134
rect 360206 542898 390690 543134
rect 390926 542898 421410 543134
rect 421646 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 79610 525454
rect 79846 525218 110330 525454
rect 110566 525218 141050 525454
rect 141286 525218 171770 525454
rect 172006 525218 202490 525454
rect 202726 525218 233210 525454
rect 233446 525218 263930 525454
rect 264166 525218 294650 525454
rect 294886 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 79610 525134
rect 79846 524898 110330 525134
rect 110566 524898 141050 525134
rect 141286 524898 171770 525134
rect 172006 524898 202490 525134
rect 202726 524898 233210 525134
rect 233446 524898 263930 525134
rect 264166 524898 294650 525134
rect 294886 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 64250 507454
rect 64486 507218 94970 507454
rect 95206 507218 125690 507454
rect 125926 507218 156410 507454
rect 156646 507218 187130 507454
rect 187366 507218 217850 507454
rect 218086 507218 248570 507454
rect 248806 507218 279290 507454
rect 279526 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 64250 507134
rect 64486 506898 94970 507134
rect 95206 506898 125690 507134
rect 125926 506898 156410 507134
rect 156646 506898 187130 507134
rect 187366 506898 217850 507134
rect 218086 506898 248570 507134
rect 248806 506898 279290 507134
rect 279526 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect 66954 481674 283574 481706
rect 66954 481438 66986 481674
rect 67222 481438 67306 481674
rect 67542 481438 102986 481674
rect 103222 481438 103306 481674
rect 103542 481438 138986 481674
rect 139222 481438 139306 481674
rect 139542 481438 174986 481674
rect 175222 481438 175306 481674
rect 175542 481438 210986 481674
rect 211222 481438 211306 481674
rect 211542 481438 246986 481674
rect 247222 481438 247306 481674
rect 247542 481438 282986 481674
rect 283222 481438 283306 481674
rect 283542 481438 283574 481674
rect 66954 481354 283574 481438
rect 66954 481118 66986 481354
rect 67222 481118 67306 481354
rect 67542 481118 102986 481354
rect 103222 481118 103306 481354
rect 103542 481118 138986 481354
rect 139222 481118 139306 481354
rect 139542 481118 174986 481354
rect 175222 481118 175306 481354
rect 175542 481118 210986 481354
rect 211222 481118 211306 481354
rect 211542 481118 246986 481354
rect 247222 481118 247306 481354
rect 247542 481118 282986 481354
rect 283222 481118 283306 481354
rect 283542 481118 283574 481354
rect 66954 481086 283574 481118
rect 63234 479834 279854 479866
rect 63234 479598 63266 479834
rect 63502 479598 63586 479834
rect 63822 479598 99266 479834
rect 99502 479598 99586 479834
rect 99822 479598 135266 479834
rect 135502 479598 135586 479834
rect 135822 479598 171266 479834
rect 171502 479598 171586 479834
rect 171822 479598 207266 479834
rect 207502 479598 207586 479834
rect 207822 479598 243266 479834
rect 243502 479598 243586 479834
rect 243822 479598 279266 479834
rect 279502 479598 279586 479834
rect 279822 479598 279854 479834
rect 63234 479514 279854 479598
rect 63234 479278 63266 479514
rect 63502 479278 63586 479514
rect 63822 479278 99266 479514
rect 99502 479278 99586 479514
rect 99822 479278 135266 479514
rect 135502 479278 135586 479514
rect 135822 479278 171266 479514
rect 171502 479278 171586 479514
rect 171822 479278 207266 479514
rect 207502 479278 207586 479514
rect 207822 479278 243266 479514
rect 243502 479278 243586 479514
rect 243822 479278 279266 479514
rect 279502 479278 279586 479514
rect 279822 479278 279854 479514
rect 63234 479246 279854 479278
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect 59514 476114 276134 476146
rect 59514 475878 59546 476114
rect 59782 475878 59866 476114
rect 60102 475878 95546 476114
rect 95782 475878 95866 476114
rect 96102 475878 131546 476114
rect 131782 475878 131866 476114
rect 132102 475878 167546 476114
rect 167782 475878 167866 476114
rect 168102 475878 203546 476114
rect 203782 475878 203866 476114
rect 204102 475878 239546 476114
rect 239782 475878 239866 476114
rect 240102 475878 275546 476114
rect 275782 475878 275866 476114
rect 276102 475878 276134 476114
rect 59514 475794 276134 475878
rect 59514 475558 59546 475794
rect 59782 475558 59866 475794
rect 60102 475558 95546 475794
rect 95782 475558 95866 475794
rect 96102 475558 131546 475794
rect 131782 475558 131866 475794
rect 132102 475558 167546 475794
rect 167782 475558 167866 475794
rect 168102 475558 203546 475794
rect 203782 475558 203866 475794
rect 204102 475558 239546 475794
rect 239782 475558 239866 475794
rect 240102 475558 275546 475794
rect 275782 475558 275866 475794
rect 276102 475558 276134 475794
rect 59514 475526 276134 475558
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 60328 453454
rect 60564 453218 196056 453454
rect 196292 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 220328 453454
rect 220564 453218 356056 453454
rect 356292 453218 380328 453454
rect 380564 453218 516056 453454
rect 516292 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 60328 453134
rect 60564 452898 196056 453134
rect 196292 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 220328 453134
rect 220564 452898 356056 453134
rect 356292 452898 380328 453134
rect 380564 452898 516056 453134
rect 516292 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 61008 435454
rect 61244 435218 195376 435454
rect 195612 435218 221008 435454
rect 221244 435218 355376 435454
rect 355612 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 381008 435454
rect 381244 435218 515376 435454
rect 515612 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 61008 435134
rect 61244 434898 195376 435134
rect 195612 434898 221008 435134
rect 221244 434898 355376 435134
rect 355612 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 381008 435134
rect 381244 434898 515376 435134
rect 515612 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 60328 417454
rect 60564 417218 196056 417454
rect 196292 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 220328 417454
rect 220564 417218 356056 417454
rect 356292 417218 380328 417454
rect 380564 417218 516056 417454
rect 516292 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 60328 417134
rect 60564 416898 196056 417134
rect 196292 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 220328 417134
rect 220564 416898 356056 417134
rect 356292 416898 380328 417134
rect 380564 416898 516056 417134
rect 516292 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 61008 399454
rect 61244 399218 195376 399454
rect 195612 399218 221008 399454
rect 221244 399218 355376 399454
rect 355612 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 381008 399454
rect 381244 399218 515376 399454
rect 515612 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 61008 399134
rect 61244 398898 195376 399134
rect 195612 398898 221008 399134
rect 221244 398898 355376 399134
rect 355612 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 381008 399134
rect 381244 398898 515376 399134
rect 515612 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect 66954 373674 499574 373706
rect 66954 373438 66986 373674
rect 67222 373438 67306 373674
rect 67542 373438 102986 373674
rect 103222 373438 103306 373674
rect 103542 373438 138986 373674
rect 139222 373438 139306 373674
rect 139542 373438 174986 373674
rect 175222 373438 175306 373674
rect 175542 373438 210986 373674
rect 211222 373438 211306 373674
rect 211542 373438 246986 373674
rect 247222 373438 247306 373674
rect 247542 373438 282986 373674
rect 283222 373438 283306 373674
rect 283542 373438 318986 373674
rect 319222 373438 319306 373674
rect 319542 373438 354986 373674
rect 355222 373438 355306 373674
rect 355542 373438 390986 373674
rect 391222 373438 391306 373674
rect 391542 373438 426986 373674
rect 427222 373438 427306 373674
rect 427542 373438 462986 373674
rect 463222 373438 463306 373674
rect 463542 373438 498986 373674
rect 499222 373438 499306 373674
rect 499542 373438 499574 373674
rect 66954 373354 499574 373438
rect 66954 373118 66986 373354
rect 67222 373118 67306 373354
rect 67542 373118 102986 373354
rect 103222 373118 103306 373354
rect 103542 373118 138986 373354
rect 139222 373118 139306 373354
rect 139542 373118 174986 373354
rect 175222 373118 175306 373354
rect 175542 373118 210986 373354
rect 211222 373118 211306 373354
rect 211542 373118 246986 373354
rect 247222 373118 247306 373354
rect 247542 373118 282986 373354
rect 283222 373118 283306 373354
rect 283542 373118 318986 373354
rect 319222 373118 319306 373354
rect 319542 373118 354986 373354
rect 355222 373118 355306 373354
rect 355542 373118 390986 373354
rect 391222 373118 391306 373354
rect 391542 373118 426986 373354
rect 427222 373118 427306 373354
rect 427542 373118 462986 373354
rect 463222 373118 463306 373354
rect 463542 373118 498986 373354
rect 499222 373118 499306 373354
rect 499542 373118 499574 373354
rect 66954 373086 499574 373118
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect 63234 369954 495854 369986
rect 63234 369718 63266 369954
rect 63502 369718 63586 369954
rect 63822 369718 99266 369954
rect 99502 369718 99586 369954
rect 99822 369718 135266 369954
rect 135502 369718 135586 369954
rect 135822 369718 171266 369954
rect 171502 369718 171586 369954
rect 171822 369718 207266 369954
rect 207502 369718 207586 369954
rect 207822 369718 243266 369954
rect 243502 369718 243586 369954
rect 243822 369718 279266 369954
rect 279502 369718 279586 369954
rect 279822 369718 315266 369954
rect 315502 369718 315586 369954
rect 315822 369718 351266 369954
rect 351502 369718 351586 369954
rect 351822 369718 387266 369954
rect 387502 369718 387586 369954
rect 387822 369718 423266 369954
rect 423502 369718 423586 369954
rect 423822 369718 459266 369954
rect 459502 369718 459586 369954
rect 459822 369718 495266 369954
rect 495502 369718 495586 369954
rect 495822 369718 495854 369954
rect 63234 369634 495854 369718
rect 63234 369398 63266 369634
rect 63502 369398 63586 369634
rect 63822 369398 99266 369634
rect 99502 369398 99586 369634
rect 99822 369398 135266 369634
rect 135502 369398 135586 369634
rect 135822 369398 171266 369634
rect 171502 369398 171586 369634
rect 171822 369398 207266 369634
rect 207502 369398 207586 369634
rect 207822 369398 243266 369634
rect 243502 369398 243586 369634
rect 243822 369398 279266 369634
rect 279502 369398 279586 369634
rect 279822 369398 315266 369634
rect 315502 369398 315586 369634
rect 315822 369398 351266 369634
rect 351502 369398 351586 369634
rect 351822 369398 387266 369634
rect 387502 369398 387586 369634
rect 387822 369398 423266 369634
rect 423502 369398 423586 369634
rect 423822 369398 459266 369634
rect 459502 369398 459586 369634
rect 459822 369398 495266 369634
rect 495502 369398 495586 369634
rect 495822 369398 495854 369634
rect 63234 369366 495854 369398
rect 59514 368114 492134 368146
rect 59514 367878 59546 368114
rect 59782 367878 59866 368114
rect 60102 367878 95546 368114
rect 95782 367878 95866 368114
rect 96102 367878 131546 368114
rect 131782 367878 131866 368114
rect 132102 367878 167546 368114
rect 167782 367878 167866 368114
rect 168102 367878 203546 368114
rect 203782 367878 203866 368114
rect 204102 367878 239546 368114
rect 239782 367878 239866 368114
rect 240102 367878 275546 368114
rect 275782 367878 275866 368114
rect 276102 367878 311546 368114
rect 311782 367878 311866 368114
rect 312102 367878 347546 368114
rect 347782 367878 347866 368114
rect 348102 367878 383546 368114
rect 383782 367878 383866 368114
rect 384102 367878 419546 368114
rect 419782 367878 419866 368114
rect 420102 367878 455546 368114
rect 455782 367878 455866 368114
rect 456102 367878 491546 368114
rect 491782 367878 491866 368114
rect 492102 367878 492134 368114
rect 59514 367794 492134 367878
rect 59514 367558 59546 367794
rect 59782 367558 59866 367794
rect 60102 367558 95546 367794
rect 95782 367558 95866 367794
rect 96102 367558 131546 367794
rect 131782 367558 131866 367794
rect 132102 367558 167546 367794
rect 167782 367558 167866 367794
rect 168102 367558 203546 367794
rect 203782 367558 203866 367794
rect 204102 367558 239546 367794
rect 239782 367558 239866 367794
rect 240102 367558 275546 367794
rect 275782 367558 275866 367794
rect 276102 367558 311546 367794
rect 311782 367558 311866 367794
rect 312102 367558 347546 367794
rect 347782 367558 347866 367794
rect 348102 367558 383546 367794
rect 383782 367558 383866 367794
rect 384102 367558 419546 367794
rect 419782 367558 419866 367794
rect 420102 367558 455546 367794
rect 455782 367558 455866 367794
rect 456102 367558 491546 367794
rect 491782 367558 491866 367794
rect 492102 367558 492134 367794
rect 59514 367526 492134 367558
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect 91794 364394 488414 364426
rect 91794 364158 91826 364394
rect 92062 364158 92146 364394
rect 92382 364158 127826 364394
rect 128062 364158 128146 364394
rect 128382 364158 163826 364394
rect 164062 364158 164146 364394
rect 164382 364158 199826 364394
rect 200062 364158 200146 364394
rect 200382 364158 235826 364394
rect 236062 364158 236146 364394
rect 236382 364158 271826 364394
rect 272062 364158 272146 364394
rect 272382 364158 307826 364394
rect 308062 364158 308146 364394
rect 308382 364158 343826 364394
rect 344062 364158 344146 364394
rect 344382 364158 379826 364394
rect 380062 364158 380146 364394
rect 380382 364158 415826 364394
rect 416062 364158 416146 364394
rect 416382 364158 451826 364394
rect 452062 364158 452146 364394
rect 452382 364158 487826 364394
rect 488062 364158 488146 364394
rect 488382 364158 488414 364394
rect 91794 364074 488414 364158
rect 91794 363838 91826 364074
rect 92062 363838 92146 364074
rect 92382 363838 127826 364074
rect 128062 363838 128146 364074
rect 128382 363838 163826 364074
rect 164062 363838 164146 364074
rect 164382 363838 199826 364074
rect 200062 363838 200146 364074
rect 200382 363838 235826 364074
rect 236062 363838 236146 364074
rect 236382 363838 271826 364074
rect 272062 363838 272146 364074
rect 272382 363838 307826 364074
rect 308062 363838 308146 364074
rect 308382 363838 343826 364074
rect 344062 363838 344146 364074
rect 344382 363838 379826 364074
rect 380062 363838 380146 364074
rect 380382 363838 415826 364074
rect 416062 363838 416146 364074
rect 416382 363838 451826 364074
rect 452062 363838 452146 364074
rect 452382 363838 487826 364074
rect 488062 363838 488146 364074
rect 488382 363838 488414 364074
rect 91794 363806 488414 363838
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 60328 345454
rect 60564 345218 196056 345454
rect 196292 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 220328 345454
rect 220564 345218 356056 345454
rect 356292 345218 380328 345454
rect 380564 345218 516056 345454
rect 516292 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 60328 345134
rect 60564 344898 196056 345134
rect 196292 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 220328 345134
rect 220564 344898 356056 345134
rect 356292 344898 380328 345134
rect 380564 344898 516056 345134
rect 516292 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 61008 327454
rect 61244 327218 195376 327454
rect 195612 327218 221008 327454
rect 221244 327218 355376 327454
rect 355612 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 381008 327454
rect 381244 327218 515376 327454
rect 515612 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 61008 327134
rect 61244 326898 195376 327134
rect 195612 326898 221008 327134
rect 221244 326898 355376 327134
rect 355612 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 381008 327134
rect 381244 326898 515376 327134
rect 515612 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 60328 309454
rect 60564 309218 196056 309454
rect 196292 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 220328 309454
rect 220564 309218 356056 309454
rect 356292 309218 380328 309454
rect 380564 309218 516056 309454
rect 516292 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 60328 309134
rect 60564 308898 196056 309134
rect 196292 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 220328 309134
rect 220564 308898 356056 309134
rect 356292 308898 380328 309134
rect 380564 308898 516056 309134
rect 516292 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 61008 291454
rect 61244 291218 195376 291454
rect 195612 291218 221008 291454
rect 221244 291218 355376 291454
rect 355612 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 381008 291454
rect 381244 291218 515376 291454
rect 515612 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 61008 291134
rect 61244 290898 195376 291134
rect 195612 290898 221008 291134
rect 221244 290898 355376 291134
rect 355612 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 381008 291134
rect 381244 290898 515376 291134
rect 515612 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect 66954 265674 499574 265706
rect 66954 265438 66986 265674
rect 67222 265438 67306 265674
rect 67542 265438 102986 265674
rect 103222 265438 103306 265674
rect 103542 265438 138986 265674
rect 139222 265438 139306 265674
rect 139542 265438 174986 265674
rect 175222 265438 175306 265674
rect 175542 265438 210986 265674
rect 211222 265438 211306 265674
rect 211542 265438 246986 265674
rect 247222 265438 247306 265674
rect 247542 265438 282986 265674
rect 283222 265438 283306 265674
rect 283542 265438 318986 265674
rect 319222 265438 319306 265674
rect 319542 265438 354986 265674
rect 355222 265438 355306 265674
rect 355542 265438 390986 265674
rect 391222 265438 391306 265674
rect 391542 265438 426986 265674
rect 427222 265438 427306 265674
rect 427542 265438 462986 265674
rect 463222 265438 463306 265674
rect 463542 265438 498986 265674
rect 499222 265438 499306 265674
rect 499542 265438 499574 265674
rect 66954 265354 499574 265438
rect 66954 265118 66986 265354
rect 67222 265118 67306 265354
rect 67542 265118 102986 265354
rect 103222 265118 103306 265354
rect 103542 265118 138986 265354
rect 139222 265118 139306 265354
rect 139542 265118 174986 265354
rect 175222 265118 175306 265354
rect 175542 265118 210986 265354
rect 211222 265118 211306 265354
rect 211542 265118 246986 265354
rect 247222 265118 247306 265354
rect 247542 265118 282986 265354
rect 283222 265118 283306 265354
rect 283542 265118 318986 265354
rect 319222 265118 319306 265354
rect 319542 265118 354986 265354
rect 355222 265118 355306 265354
rect 355542 265118 390986 265354
rect 391222 265118 391306 265354
rect 391542 265118 426986 265354
rect 427222 265118 427306 265354
rect 427542 265118 462986 265354
rect 463222 265118 463306 265354
rect 463542 265118 498986 265354
rect 499222 265118 499306 265354
rect 499542 265118 499574 265354
rect 66954 265086 499574 265118
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect 63234 261954 495854 261986
rect 63234 261718 63266 261954
rect 63502 261718 63586 261954
rect 63822 261718 99266 261954
rect 99502 261718 99586 261954
rect 99822 261718 135266 261954
rect 135502 261718 135586 261954
rect 135822 261718 171266 261954
rect 171502 261718 171586 261954
rect 171822 261718 207266 261954
rect 207502 261718 207586 261954
rect 207822 261718 243266 261954
rect 243502 261718 243586 261954
rect 243822 261718 279266 261954
rect 279502 261718 279586 261954
rect 279822 261718 315266 261954
rect 315502 261718 315586 261954
rect 315822 261718 351266 261954
rect 351502 261718 351586 261954
rect 351822 261718 387266 261954
rect 387502 261718 387586 261954
rect 387822 261718 423266 261954
rect 423502 261718 423586 261954
rect 423822 261718 459266 261954
rect 459502 261718 459586 261954
rect 459822 261718 495266 261954
rect 495502 261718 495586 261954
rect 495822 261718 495854 261954
rect 63234 261634 495854 261718
rect 63234 261398 63266 261634
rect 63502 261398 63586 261634
rect 63822 261398 99266 261634
rect 99502 261398 99586 261634
rect 99822 261398 135266 261634
rect 135502 261398 135586 261634
rect 135822 261398 171266 261634
rect 171502 261398 171586 261634
rect 171822 261398 207266 261634
rect 207502 261398 207586 261634
rect 207822 261398 243266 261634
rect 243502 261398 243586 261634
rect 243822 261398 279266 261634
rect 279502 261398 279586 261634
rect 279822 261398 315266 261634
rect 315502 261398 315586 261634
rect 315822 261398 351266 261634
rect 351502 261398 351586 261634
rect 351822 261398 387266 261634
rect 387502 261398 387586 261634
rect 387822 261398 423266 261634
rect 423502 261398 423586 261634
rect 423822 261398 459266 261634
rect 459502 261398 459586 261634
rect 459822 261398 495266 261634
rect 495502 261398 495586 261634
rect 495822 261398 495854 261634
rect 63234 261366 495854 261398
rect 59514 260114 492134 260146
rect 59514 259878 59546 260114
rect 59782 259878 59866 260114
rect 60102 259878 95546 260114
rect 95782 259878 95866 260114
rect 96102 259878 131546 260114
rect 131782 259878 131866 260114
rect 132102 259878 167546 260114
rect 167782 259878 167866 260114
rect 168102 259878 203546 260114
rect 203782 259878 203866 260114
rect 204102 259878 239546 260114
rect 239782 259878 239866 260114
rect 240102 259878 275546 260114
rect 275782 259878 275866 260114
rect 276102 259878 311546 260114
rect 311782 259878 311866 260114
rect 312102 259878 347546 260114
rect 347782 259878 347866 260114
rect 348102 259878 383546 260114
rect 383782 259878 383866 260114
rect 384102 259878 419546 260114
rect 419782 259878 419866 260114
rect 420102 259878 455546 260114
rect 455782 259878 455866 260114
rect 456102 259878 491546 260114
rect 491782 259878 491866 260114
rect 492102 259878 492134 260114
rect 59514 259794 492134 259878
rect 59514 259558 59546 259794
rect 59782 259558 59866 259794
rect 60102 259558 95546 259794
rect 95782 259558 95866 259794
rect 96102 259558 131546 259794
rect 131782 259558 131866 259794
rect 132102 259558 167546 259794
rect 167782 259558 167866 259794
rect 168102 259558 203546 259794
rect 203782 259558 203866 259794
rect 204102 259558 239546 259794
rect 239782 259558 239866 259794
rect 240102 259558 275546 259794
rect 275782 259558 275866 259794
rect 276102 259558 311546 259794
rect 311782 259558 311866 259794
rect 312102 259558 347546 259794
rect 347782 259558 347866 259794
rect 348102 259558 383546 259794
rect 383782 259558 383866 259794
rect 384102 259558 419546 259794
rect 419782 259558 419866 259794
rect 420102 259558 455546 259794
rect 455782 259558 455866 259794
rect 456102 259558 491546 259794
rect 491782 259558 491866 259794
rect 492102 259558 492134 259794
rect 59514 259526 492134 259558
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect 91794 256394 488414 256426
rect 91794 256158 91826 256394
rect 92062 256158 92146 256394
rect 92382 256158 127826 256394
rect 128062 256158 128146 256394
rect 128382 256158 163826 256394
rect 164062 256158 164146 256394
rect 164382 256158 199826 256394
rect 200062 256158 200146 256394
rect 200382 256158 235826 256394
rect 236062 256158 236146 256394
rect 236382 256158 271826 256394
rect 272062 256158 272146 256394
rect 272382 256158 307826 256394
rect 308062 256158 308146 256394
rect 308382 256158 343826 256394
rect 344062 256158 344146 256394
rect 344382 256158 379826 256394
rect 380062 256158 380146 256394
rect 380382 256158 415826 256394
rect 416062 256158 416146 256394
rect 416382 256158 451826 256394
rect 452062 256158 452146 256394
rect 452382 256158 487826 256394
rect 488062 256158 488146 256394
rect 488382 256158 488414 256394
rect 91794 256074 488414 256158
rect 91794 255838 91826 256074
rect 92062 255838 92146 256074
rect 92382 255838 127826 256074
rect 128062 255838 128146 256074
rect 128382 255838 163826 256074
rect 164062 255838 164146 256074
rect 164382 255838 199826 256074
rect 200062 255838 200146 256074
rect 200382 255838 235826 256074
rect 236062 255838 236146 256074
rect 236382 255838 271826 256074
rect 272062 255838 272146 256074
rect 272382 255838 307826 256074
rect 308062 255838 308146 256074
rect 308382 255838 343826 256074
rect 344062 255838 344146 256074
rect 344382 255838 379826 256074
rect 380062 255838 380146 256074
rect 380382 255838 415826 256074
rect 416062 255838 416146 256074
rect 416382 255838 451826 256074
rect 452062 255838 452146 256074
rect 452382 255838 487826 256074
rect 488062 255838 488146 256074
rect 488382 255838 488414 256074
rect 91794 255806 488414 255838
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 60328 237454
rect 60564 237218 196056 237454
rect 196292 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 220328 237454
rect 220564 237218 356056 237454
rect 356292 237218 380328 237454
rect 380564 237218 516056 237454
rect 516292 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 60328 237134
rect 60564 236898 196056 237134
rect 196292 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 220328 237134
rect 220564 236898 356056 237134
rect 356292 236898 380328 237134
rect 380564 236898 516056 237134
rect 516292 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 61008 219454
rect 61244 219218 195376 219454
rect 195612 219218 221008 219454
rect 221244 219218 355376 219454
rect 355612 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 381008 219454
rect 381244 219218 515376 219454
rect 515612 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 61008 219134
rect 61244 218898 195376 219134
rect 195612 218898 221008 219134
rect 221244 218898 355376 219134
rect 355612 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 381008 219134
rect 381244 218898 515376 219134
rect 515612 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 60328 201454
rect 60564 201218 196056 201454
rect 196292 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 220328 201454
rect 220564 201218 356056 201454
rect 356292 201218 380328 201454
rect 380564 201218 516056 201454
rect 516292 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 60328 201134
rect 60564 200898 196056 201134
rect 196292 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 220328 201134
rect 220564 200898 356056 201134
rect 356292 200898 380328 201134
rect 380564 200898 516056 201134
rect 516292 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 61008 183454
rect 61244 183218 195376 183454
rect 195612 183218 221008 183454
rect 221244 183218 355376 183454
rect 355612 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 381008 183454
rect 381244 183218 515376 183454
rect 515612 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 61008 183134
rect 61244 182898 195376 183134
rect 195612 182898 221008 183134
rect 221244 182898 355376 183134
rect 355612 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 381008 183134
rect 381244 182898 515376 183134
rect 515612 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 84986 158614
rect 85222 158378 85306 158614
rect 85542 158378 120986 158614
rect 121222 158378 121306 158614
rect 121542 158378 156986 158614
rect 157222 158378 157306 158614
rect 157542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 84986 158294
rect 85222 158058 85306 158294
rect 85542 158058 120986 158294
rect 121222 158058 121306 158294
rect 121542 158058 156986 158294
rect 157222 158058 157306 158294
rect 157542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect 66954 157674 499574 157706
rect 66954 157438 66986 157674
rect 67222 157438 67306 157674
rect 67542 157438 102986 157674
rect 103222 157438 103306 157674
rect 103542 157438 138986 157674
rect 139222 157438 139306 157674
rect 139542 157438 174986 157674
rect 175222 157438 175306 157674
rect 175542 157438 210986 157674
rect 211222 157438 211306 157674
rect 211542 157438 246986 157674
rect 247222 157438 247306 157674
rect 247542 157438 282986 157674
rect 283222 157438 283306 157674
rect 283542 157438 318986 157674
rect 319222 157438 319306 157674
rect 319542 157438 354986 157674
rect 355222 157438 355306 157674
rect 355542 157438 390986 157674
rect 391222 157438 391306 157674
rect 391542 157438 426986 157674
rect 427222 157438 427306 157674
rect 427542 157438 462986 157674
rect 463222 157438 463306 157674
rect 463542 157438 498986 157674
rect 499222 157438 499306 157674
rect 499542 157438 499574 157674
rect 66954 157354 499574 157438
rect 66954 157118 66986 157354
rect 67222 157118 67306 157354
rect 67542 157118 102986 157354
rect 103222 157118 103306 157354
rect 103542 157118 138986 157354
rect 139222 157118 139306 157354
rect 139542 157118 174986 157354
rect 175222 157118 175306 157354
rect 175542 157118 210986 157354
rect 211222 157118 211306 157354
rect 211542 157118 246986 157354
rect 247222 157118 247306 157354
rect 247542 157118 282986 157354
rect 283222 157118 283306 157354
rect 283542 157118 318986 157354
rect 319222 157118 319306 157354
rect 319542 157118 354986 157354
rect 355222 157118 355306 157354
rect 355542 157118 390986 157354
rect 391222 157118 391306 157354
rect 391542 157118 426986 157354
rect 427222 157118 427306 157354
rect 427542 157118 462986 157354
rect 463222 157118 463306 157354
rect 463542 157118 498986 157354
rect 499222 157118 499306 157354
rect 499542 157118 499574 157354
rect 66954 157086 499574 157118
rect 63234 155834 495854 155866
rect 63234 155598 63266 155834
rect 63502 155598 63586 155834
rect 63822 155598 99266 155834
rect 99502 155598 99586 155834
rect 99822 155598 135266 155834
rect 135502 155598 135586 155834
rect 135822 155598 171266 155834
rect 171502 155598 171586 155834
rect 171822 155598 207266 155834
rect 207502 155598 207586 155834
rect 207822 155598 243266 155834
rect 243502 155598 243586 155834
rect 243822 155598 279266 155834
rect 279502 155598 279586 155834
rect 279822 155598 315266 155834
rect 315502 155598 315586 155834
rect 315822 155598 351266 155834
rect 351502 155598 351586 155834
rect 351822 155598 387266 155834
rect 387502 155598 387586 155834
rect 387822 155598 423266 155834
rect 423502 155598 423586 155834
rect 423822 155598 459266 155834
rect 459502 155598 459586 155834
rect 459822 155598 495266 155834
rect 495502 155598 495586 155834
rect 495822 155598 495854 155834
rect 63234 155514 495854 155598
rect 63234 155278 63266 155514
rect 63502 155278 63586 155514
rect 63822 155278 99266 155514
rect 99502 155278 99586 155514
rect 99822 155278 135266 155514
rect 135502 155278 135586 155514
rect 135822 155278 171266 155514
rect 171502 155278 171586 155514
rect 171822 155278 207266 155514
rect 207502 155278 207586 155514
rect 207822 155278 243266 155514
rect 243502 155278 243586 155514
rect 243822 155278 279266 155514
rect 279502 155278 279586 155514
rect 279822 155278 315266 155514
rect 315502 155278 315586 155514
rect 315822 155278 351266 155514
rect 351502 155278 351586 155514
rect 351822 155278 387266 155514
rect 387502 155278 387586 155514
rect 387822 155278 423266 155514
rect 423502 155278 423586 155514
rect 423822 155278 459266 155514
rect 459502 155278 459586 155514
rect 459822 155278 495266 155514
rect 495502 155278 495586 155514
rect 495822 155278 495854 155514
rect 63234 155246 495854 155278
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 81266 154894
rect 81502 154658 81586 154894
rect 81822 154658 117266 154894
rect 117502 154658 117586 154894
rect 117822 154658 153266 154894
rect 153502 154658 153586 154894
rect 153822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 225266 154894
rect 225502 154658 225586 154894
rect 225822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 81266 154574
rect 81502 154338 81586 154574
rect 81822 154338 117266 154574
rect 117502 154338 117586 154574
rect 117822 154338 153266 154574
rect 153502 154338 153586 154574
rect 153822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 225266 154574
rect 225502 154338 225586 154574
rect 225822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect 59514 152114 492134 152146
rect 59514 151878 59546 152114
rect 59782 151878 59866 152114
rect 60102 151878 95546 152114
rect 95782 151878 95866 152114
rect 96102 151878 131546 152114
rect 131782 151878 131866 152114
rect 132102 151878 167546 152114
rect 167782 151878 167866 152114
rect 168102 151878 203546 152114
rect 203782 151878 203866 152114
rect 204102 151878 239546 152114
rect 239782 151878 239866 152114
rect 240102 151878 275546 152114
rect 275782 151878 275866 152114
rect 276102 151878 311546 152114
rect 311782 151878 311866 152114
rect 312102 151878 347546 152114
rect 347782 151878 347866 152114
rect 348102 151878 383546 152114
rect 383782 151878 383866 152114
rect 384102 151878 419546 152114
rect 419782 151878 419866 152114
rect 420102 151878 455546 152114
rect 455782 151878 455866 152114
rect 456102 151878 491546 152114
rect 491782 151878 491866 152114
rect 492102 151878 492134 152114
rect 59514 151794 492134 151878
rect 59514 151558 59546 151794
rect 59782 151558 59866 151794
rect 60102 151558 95546 151794
rect 95782 151558 95866 151794
rect 96102 151558 131546 151794
rect 131782 151558 131866 151794
rect 132102 151558 167546 151794
rect 167782 151558 167866 151794
rect 168102 151558 203546 151794
rect 203782 151558 203866 151794
rect 204102 151558 239546 151794
rect 239782 151558 239866 151794
rect 240102 151558 275546 151794
rect 275782 151558 275866 151794
rect 276102 151558 311546 151794
rect 311782 151558 311866 151794
rect 312102 151558 347546 151794
rect 347782 151558 347866 151794
rect 348102 151558 383546 151794
rect 383782 151558 383866 151794
rect 384102 151558 419546 151794
rect 419782 151558 419866 151794
rect 420102 151558 455546 151794
rect 455782 151558 455866 151794
rect 456102 151558 491546 151794
rect 491782 151558 491866 151794
rect 492102 151558 492134 151794
rect 59514 151526 492134 151558
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 77546 151174
rect 77782 150938 77866 151174
rect 78102 150938 113546 151174
rect 113782 150938 113866 151174
rect 114102 150938 149546 151174
rect 149782 150938 149866 151174
rect 150102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 221546 151174
rect 221782 150938 221866 151174
rect 222102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 77546 150854
rect 77782 150618 77866 150854
rect 78102 150618 113546 150854
rect 113782 150618 113866 150854
rect 114102 150618 149546 150854
rect 149782 150618 149866 150854
rect 150102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 221546 150854
rect 221782 150618 221866 150854
rect 222102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect 91794 148394 488414 148426
rect 91794 148158 91826 148394
rect 92062 148158 92146 148394
rect 92382 148158 127826 148394
rect 128062 148158 128146 148394
rect 128382 148158 163826 148394
rect 164062 148158 164146 148394
rect 164382 148158 199826 148394
rect 200062 148158 200146 148394
rect 200382 148158 235826 148394
rect 236062 148158 236146 148394
rect 236382 148158 271826 148394
rect 272062 148158 272146 148394
rect 272382 148158 307826 148394
rect 308062 148158 308146 148394
rect 308382 148158 343826 148394
rect 344062 148158 344146 148394
rect 344382 148158 379826 148394
rect 380062 148158 380146 148394
rect 380382 148158 415826 148394
rect 416062 148158 416146 148394
rect 416382 148158 451826 148394
rect 452062 148158 452146 148394
rect 452382 148158 487826 148394
rect 488062 148158 488146 148394
rect 488382 148158 488414 148394
rect 91794 148074 488414 148158
rect 91794 147838 91826 148074
rect 92062 147838 92146 148074
rect 92382 147838 127826 148074
rect 128062 147838 128146 148074
rect 128382 147838 163826 148074
rect 164062 147838 164146 148074
rect 164382 147838 199826 148074
rect 200062 147838 200146 148074
rect 200382 147838 235826 148074
rect 236062 147838 236146 148074
rect 236382 147838 271826 148074
rect 272062 147838 272146 148074
rect 272382 147838 307826 148074
rect 308062 147838 308146 148074
rect 308382 147838 343826 148074
rect 344062 147838 344146 148074
rect 344382 147838 379826 148074
rect 380062 147838 380146 148074
rect 380382 147838 415826 148074
rect 416062 147838 416146 148074
rect 416382 147838 451826 148074
rect 452062 147838 452146 148074
rect 452382 147838 487826 148074
rect 488062 147838 488146 148074
rect 488382 147838 488414 148074
rect 91794 147806 488414 147838
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 73826 147454
rect 74062 147218 74146 147454
rect 74382 147218 109826 147454
rect 110062 147218 110146 147454
rect 110382 147218 145826 147454
rect 146062 147218 146146 147454
rect 146382 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 217826 147454
rect 218062 147218 218146 147454
rect 218382 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 73826 147134
rect 74062 146898 74146 147134
rect 74382 146898 109826 147134
rect 110062 146898 110146 147134
rect 110382 146898 145826 147134
rect 146062 146898 146146 147134
rect 146382 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 217826 147134
rect 218062 146898 218146 147134
rect 218382 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 60328 129454
rect 60564 129218 196056 129454
rect 196292 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 220328 129454
rect 220564 129218 356056 129454
rect 356292 129218 380328 129454
rect 380564 129218 516056 129454
rect 516292 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 60328 129134
rect 60564 128898 196056 129134
rect 196292 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 220328 129134
rect 220564 128898 356056 129134
rect 356292 128898 380328 129134
rect 380564 128898 516056 129134
rect 516292 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 61008 111454
rect 61244 111218 195376 111454
rect 195612 111218 221008 111454
rect 221244 111218 355376 111454
rect 355612 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 381008 111454
rect 381244 111218 515376 111454
rect 515612 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 61008 111134
rect 61244 110898 195376 111134
rect 195612 110898 221008 111134
rect 221244 110898 355376 111134
rect 355612 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 381008 111134
rect 381244 110898 515376 111134
rect 515612 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 60328 93454
rect 60564 93218 196056 93454
rect 196292 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 220328 93454
rect 220564 93218 356056 93454
rect 356292 93218 380328 93454
rect 380564 93218 516056 93454
rect 516292 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 60328 93134
rect 60564 92898 196056 93134
rect 196292 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 220328 93134
rect 220564 92898 356056 93134
rect 356292 92898 380328 93134
rect 380564 92898 516056 93134
rect 516292 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 61008 75454
rect 61244 75218 195376 75454
rect 195612 75218 221008 75454
rect 221244 75218 355376 75454
rect 355612 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 381008 75454
rect 381244 75218 515376 75454
rect 515612 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 61008 75134
rect 61244 74898 195376 75134
rect 195612 74898 221008 75134
rect 221244 74898 355376 75134
rect 355612 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 381008 75134
rect 381244 74898 515376 75134
rect 515612 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_2kbyte_1rw1r_32x512_8  agent_1_sram2k_inst0
timestamp 0
transform 1 0 60000 0 1 60000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  agent_1_sram2k_inst1
timestamp 0
transform 1 0 60000 0 1 167000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  agent_1_sram2k_inst2
timestamp 0
transform 1 0 60000 0 1 274000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  codemaker_sram2k_inst0
timestamp 0
transform 1 0 380000 0 1 60000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  codemaker_sram2k_inst1
timestamp 0
transform 1 0 380000 0 1 167000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  codemaker_sram2k_inst2
timestamp 0
transform 1 0 380000 0 1 274000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  codemaker_sram2k_inst3
timestamp 0
transform 1 0 380000 0 1 381000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst0
timestamp 0
transform 1 0 60000 0 1 381000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst1
timestamp 0
transform 1 0 220000 0 1 60000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst2
timestamp 0
transform 1 0 220000 0 1 167000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst3
timestamp 0
transform 1 0 220000 0 1 274000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  control_tower_sram2k_inst4
timestamp 0
transform 1 0 220000 0 1 381000
box 0 0 136620 83308
use VerySimpleCPU_core  inst_agent_1
timestamp 0
transform 1 0 60000 0 1 580000
box 0 0 60955 63099
use VerySimpleCPU_core  inst_codemaker
timestamp 0
transform 1 0 240000 0 1 580000
box 0 0 60955 63099
use VerySimpleCPU_core  inst_control_tower
timestamp 0
transform 1 0 150000 0 1 580000
box 0 0 60955 63099
use main_controller  inst_main_controller
timestamp 0
transform 1 0 60000 0 1 493000
box 0 0 240000 60000
use main_memory  inst_main_memory
timestamp 0
transform 1 0 325000 0 1 534000
box 0 0 108889 111033
use uart  inst_uart
timestamp 0
transform 1 0 460000 0 1 590000
box 0 0 50000 50000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s 73794 561806 290414 562426 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 145308 74414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 145308 110414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 145308 146414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 145308 182414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 145308 218414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 145308 254414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 145308 290414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 145308 326414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 145308 398414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 145308 434414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 145308 470414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 145308 506414 165000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 252308 74414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 252308 110414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 252308 146414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 252308 182414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 252308 218414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 252308 254414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 252308 290414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 252308 326414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 252308 398414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 252308 434414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 252308 470414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 252308 506414 272000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 359308 74414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 359308 110414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 359308 146414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 359308 182414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 359308 218414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 359308 254414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 359308 290414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 359308 326414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 359308 398414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 359308 434414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 359308 470414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 359308 506414 379000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 466308 74414 491000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 466308 110414 491000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 466308 146414 491000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 466308 182414 491000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 466308 218414 491000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 466308 254414 491000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 466308 290414 491000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 466308 326414 532000 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 532000 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 466308 398414 532000 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 466308 434414 532000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 555000 74414 578000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 555000 110414 578000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 555000 182414 578000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 555000 254414 578000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 555000 290414 578000 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 466308 470414 588000 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 466308 506414 588000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 645099 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 645099 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 555000 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 645099 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 555000 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 645099 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 645099 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 647033 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 647033 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 647033 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 647033 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 642000 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 642000 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s 77514 565526 294134 566146 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 145308 78134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 145308 114134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 145308 150134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 145308 186134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 145308 222134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 145308 258134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 145308 294134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 145308 330134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 145308 402134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 145308 438134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 145308 474134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 145308 510134 165000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 252308 78134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 252308 114134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 252308 150134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 252308 186134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 252308 222134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 252308 258134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 252308 294134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 252308 330134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 252308 402134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 252308 438134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 252308 474134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 252308 510134 272000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 359308 78134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 359308 114134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 359308 150134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 359308 186134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 359308 222134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 359308 258134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 359308 294134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 359308 330134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 359308 402134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 359308 438134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 359308 474134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 359308 510134 379000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 466308 78134 491000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 466308 114134 491000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 466308 150134 491000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 466308 186134 491000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 466308 222134 491000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 466308 258134 491000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 466308 294134 491000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 466308 330134 532000 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 532000 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 466308 402134 532000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 555000 78134 578000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 555000 114134 578000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 555000 150134 578000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 555000 186134 578000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 555000 258134 578000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 555000 294134 578000 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 466308 474134 588000 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 466308 510134 588000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 645099 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 645099 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 645099 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 645099 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 555000 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 645099 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 645099 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 647033 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 647033 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 647033 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 466308 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 642000 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 642000 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s 81234 567366 297854 567986 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 145308 81854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 145308 117854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 145308 153854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 145308 189854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 145308 225854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 145308 261854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 145308 297854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 145308 333854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 145308 405854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 145308 441854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 145308 477854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 145308 513854 165000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 252308 81854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 252308 117854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 252308 153854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 252308 189854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 252308 225854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 252308 261854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 252308 297854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 252308 333854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 252308 405854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 252308 441854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 252308 477854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 252308 513854 272000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 359308 81854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 359308 117854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 359308 153854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 359308 189854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 359308 225854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 359308 261854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 359308 297854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 359308 333854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 359308 405854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 359308 441854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 359308 477854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 359308 513854 379000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 466308 81854 491000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 466308 117854 491000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 466308 153854 491000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 466308 189854 491000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 466308 225854 491000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 466308 261854 491000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 466308 297854 491000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 466308 333854 532000 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 532000 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 466308 405854 532000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 555000 81854 578000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 555000 117854 578000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 555000 153854 578000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 555000 189854 578000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 555000 261854 578000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 555000 297854 578000 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 466308 477854 588000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 645099 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 645099 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 645099 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 645099 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 555000 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 645099 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 645099 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 647033 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 647033 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 647033 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 466308 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 642000 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 466308 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s 84954 571086 301574 571706 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 145308 85574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 145308 121574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 145308 157574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 145308 193574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 145308 229574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 145308 265574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 145308 301574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 145308 337574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 145308 409574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 145308 445574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 145308 481574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 145308 517574 165000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 252308 85574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 252308 121574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 252308 157574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 252308 193574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 252308 229574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 252308 265574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 252308 301574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 252308 337574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 252308 409574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 252308 445574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 252308 481574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 252308 517574 272000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 359308 85574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 359308 121574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 359308 157574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 359308 193574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 359308 229574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 359308 265574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 359308 301574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 359308 337574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 359308 409574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 359308 445574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 359308 481574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 359308 517574 379000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 466308 85574 491000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 466308 121574 491000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 466308 157574 491000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 466308 193574 491000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 466308 229574 491000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 466308 265574 491000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 466308 301574 491000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 466308 337574 532000 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 532000 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 466308 409574 532000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 555000 85574 578000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 555000 121574 578000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 555000 157574 578000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 555000 193574 578000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 555000 265574 578000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 555000 301574 578000 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 466308 481574 588000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 645099 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 645099 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 645099 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 645099 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 555000 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 645099 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 645099 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 647033 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 647033 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 647033 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 466308 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 642000 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 466308 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 63234 155246 495854 155866 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 63234 261366 495854 261986 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 63234 369366 495854 369986 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s 63234 479246 279854 479866 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 145308 63854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 145308 99854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 145308 135854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 145308 171854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 145308 243854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 145308 279854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 145308 315854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 145308 351854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 145308 387854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 145308 423854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 145308 459854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 145308 495854 165000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 252308 63854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 252308 99854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 252308 135854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 252308 171854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 252308 243854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 252308 279854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 252308 315854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 252308 351854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 252308 387854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 252308 423854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 252308 459854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 252308 495854 272000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 359308 63854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 359308 99854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 359308 135854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 359308 171854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 359308 243854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 359308 279854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 359308 315854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 359308 351854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 359308 387854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 359308 423854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 359308 459854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 359308 495854 379000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 466308 63854 491000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 466308 99854 491000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 466308 135854 491000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 466308 171854 491000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 491000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 466308 243854 491000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 466308 279854 491000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 466308 351854 532000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 466308 387854 532000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 466308 423854 532000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 555000 63854 578000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 555000 99854 578000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 555000 171854 578000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 555000 207854 578000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 555000 243854 578000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 555000 279854 578000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 466308 459854 588000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 466308 495854 588000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 645099 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 645099 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 555000 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 645099 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 645099 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 645099 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 645099 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 466308 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 647033 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 647033 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 647033 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 642000 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 642000 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 66954 157086 499574 157706 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 66954 265086 499574 265706 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 66954 373086 499574 373706 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s 66954 481086 283574 481706 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 145308 67574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 145308 103574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 145308 139574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 145308 175574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 145308 247574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 145308 283574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 145308 319574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 145308 355574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 145308 391574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 145308 427574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 145308 463574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 145308 499574 165000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 252308 67574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 252308 103574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 252308 139574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 252308 175574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 252308 247574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 252308 283574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 252308 319574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 252308 355574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 252308 391574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 252308 427574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 252308 463574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 252308 499574 272000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 359308 67574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 359308 103574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 359308 139574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 359308 175574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 359308 247574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 359308 283574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 359308 319574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 359308 355574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 359308 391574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 359308 427574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 359308 463574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 359308 499574 379000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 466308 67574 491000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 466308 103574 491000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 466308 139574 491000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 466308 175574 491000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 491000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 466308 247574 491000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 466308 283574 491000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 466308 355574 532000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 466308 391574 532000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 466308 427574 532000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 555000 67574 578000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 555000 103574 578000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 555000 175574 578000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 555000 211574 578000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 555000 247574 578000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 555000 283574 578000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 466308 463574 588000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 466308 499574 588000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 645099 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 645099 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 555000 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 645099 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 645099 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 645099 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 645099 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 466308 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 647033 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 647033 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 647033 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 642000 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 642000 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 91794 147806 488414 148426 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 91794 255806 488414 256426 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s 91794 363806 488414 364426 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 145308 92414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 145308 128414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 145308 164414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 145308 236414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 145308 272414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 145308 308414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 145308 344414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 145308 380414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 145308 416414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 145308 452414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 145308 488414 165000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 252308 92414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 252308 128414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 252308 164414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 252308 236414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 252308 272414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 252308 308414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 252308 344414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 252308 380414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 252308 416414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 252308 452414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 252308 488414 272000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 359308 92414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 359308 128414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 359308 164414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 359308 236414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 359308 272414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 359308 308414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 359308 344414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 359308 380414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 359308 416414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 359308 452414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 359308 488414 379000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 466308 92414 491000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 466308 128414 491000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 466308 164414 491000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 491000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 466308 236414 491000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 466308 272414 491000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 466308 344414 532000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 466308 380414 532000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 466308 416414 532000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 555000 92414 578000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 555000 164414 578000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 555000 200414 578000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 555000 272414 578000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 466308 488414 588000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 645099 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 555000 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 645099 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 645099 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 555000 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 645099 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 466308 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 647033 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 647033 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 647033 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 466308 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 642000 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 59514 151526 492134 152146 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 59514 259526 492134 260146 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 59514 367526 492134 368146 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s 59514 475526 276134 476146 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 145308 60134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 145308 96134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 145308 132134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 145308 168134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 145308 240134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 145308 276134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 145308 312134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 145308 348134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 145308 384134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 145308 420134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 145308 456134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 145308 492134 165000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 252308 60134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 252308 96134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 252308 132134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 252308 168134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 252308 240134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 252308 276134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 252308 312134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 252308 348134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 252308 384134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 252308 420134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 252308 456134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 252308 492134 272000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 359308 60134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 359308 96134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 359308 132134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 359308 168134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 359308 240134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 359308 276134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 359308 312134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 359308 348134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 359308 384134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 359308 420134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 359308 456134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 359308 492134 379000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 466308 60134 491000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 466308 96134 491000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 466308 132134 491000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 466308 168134 491000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 491000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 466308 240134 491000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 466308 276134 491000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 466308 348134 532000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 466308 384134 532000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 466308 420134 532000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 555000 60134 578000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 555000 96134 578000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 555000 168134 578000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 555000 204134 578000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 555000 240134 578000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 555000 276134 578000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 466308 492134 588000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 645099 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 645099 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 555000 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 645099 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 645099 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 645099 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 645099 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 466308 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 647033 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 647033 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 647033 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 466308 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 642000 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
