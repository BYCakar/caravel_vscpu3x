VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO VerySimpleCPU_core
  CLASS BLOCK ;
  FOREIGN VerySimpleCPU_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 304.775 BY 315.495 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END clk
  PIN done
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END done
  PIN mem_ctrl_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 311.495 190.350 315.495 ;
    END
  END mem_ctrl_addr[0]
  PIN mem_ctrl_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 311.495 161.370 315.495 ;
    END
  END mem_ctrl_addr[10]
  PIN mem_ctrl_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 300.775 255.040 304.775 255.640 ;
    END
  END mem_ctrl_addr[11]
  PIN mem_ctrl_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END mem_ctrl_addr[12]
  PIN mem_ctrl_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END mem_ctrl_addr[13]
  PIN mem_ctrl_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END mem_ctrl_addr[1]
  PIN mem_ctrl_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END mem_ctrl_addr[2]
  PIN mem_ctrl_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END mem_ctrl_addr[3]
  PIN mem_ctrl_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END mem_ctrl_addr[4]
  PIN mem_ctrl_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 300.775 40.840 304.775 41.440 ;
    END
  END mem_ctrl_addr[5]
  PIN mem_ctrl_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 300.775 299.240 304.775 299.840 ;
    END
  END mem_ctrl_addr[6]
  PIN mem_ctrl_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 300.775 132.640 304.775 133.240 ;
    END
  END mem_ctrl_addr[7]
  PIN mem_ctrl_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 300.775 224.440 304.775 225.040 ;
    END
  END mem_ctrl_addr[8]
  PIN mem_ctrl_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 300.775 10.240 304.775 10.840 ;
    END
  END mem_ctrl_addr[9]
  PIN mem_ctrl_in[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 300.775 85.040 304.775 85.640 ;
    END
  END mem_ctrl_in[0]
  PIN mem_ctrl_in[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END mem_ctrl_in[10]
  PIN mem_ctrl_in[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 311.495 219.330 315.495 ;
    END
  END mem_ctrl_in[11]
  PIN mem_ctrl_in[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 300.775 54.440 304.775 55.040 ;
    END
  END mem_ctrl_in[12]
  PIN mem_ctrl_in[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 311.495 145.270 315.495 ;
    END
  END mem_ctrl_in[13]
  PIN mem_ctrl_in[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 300.775 193.840 304.775 194.440 ;
    END
  END mem_ctrl_in[14]
  PIN mem_ctrl_in[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 300.775 115.640 304.775 116.240 ;
    END
  END mem_ctrl_in[15]
  PIN mem_ctrl_in[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END mem_ctrl_in[16]
  PIN mem_ctrl_in[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END mem_ctrl_in[17]
  PIN mem_ctrl_in[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END mem_ctrl_in[18]
  PIN mem_ctrl_in[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 311.495 87.310 315.495 ;
    END
  END mem_ctrl_in[19]
  PIN mem_ctrl_in[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 300.775 207.440 304.775 208.040 ;
    END
  END mem_ctrl_in[1]
  PIN mem_ctrl_in[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 300.775 102.040 304.775 102.640 ;
    END
  END mem_ctrl_in[20]
  PIN mem_ctrl_in[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 311.495 174.250 315.495 ;
    END
  END mem_ctrl_in[21]
  PIN mem_ctrl_in[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 300.775 268.640 304.775 269.240 ;
    END
  END mem_ctrl_in[22]
  PIN mem_ctrl_in[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END mem_ctrl_in[23]
  PIN mem_ctrl_in[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 311.495 232.210 315.495 ;
    END
  END mem_ctrl_in[24]
  PIN mem_ctrl_in[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 311.495 290.170 315.495 ;
    END
  END mem_ctrl_in[25]
  PIN mem_ctrl_in[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 311.495 16.470 315.495 ;
    END
  END mem_ctrl_in[26]
  PIN mem_ctrl_in[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END mem_ctrl_in[27]
  PIN mem_ctrl_in[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END mem_ctrl_in[28]
  PIN mem_ctrl_in[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END mem_ctrl_in[29]
  PIN mem_ctrl_in[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 300.775 238.040 304.775 238.640 ;
    END
  END mem_ctrl_in[2]
  PIN mem_ctrl_in[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END mem_ctrl_in[30]
  PIN mem_ctrl_in[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END mem_ctrl_in[31]
  PIN mem_ctrl_in[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END mem_ctrl_in[3]
  PIN mem_ctrl_in[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END mem_ctrl_in[4]
  PIN mem_ctrl_in[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 311.495 58.330 315.495 ;
    END
  END mem_ctrl_in[5]
  PIN mem_ctrl_in[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END mem_ctrl_in[6]
  PIN mem_ctrl_in[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END mem_ctrl_in[7]
  PIN mem_ctrl_in[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 311.495 0.370 315.495 ;
    END
  END mem_ctrl_in[8]
  PIN mem_ctrl_in[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END mem_ctrl_in[9]
  PIN mem_ctrl_out[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 311.495 103.410 315.495 ;
    END
  END mem_ctrl_out[0]
  PIN mem_ctrl_out[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 300.775 71.440 304.775 72.040 ;
    END
  END mem_ctrl_out[10]
  PIN mem_ctrl_out[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END mem_ctrl_out[11]
  PIN mem_ctrl_out[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END mem_ctrl_out[12]
  PIN mem_ctrl_out[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END mem_ctrl_out[13]
  PIN mem_ctrl_out[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END mem_ctrl_out[14]
  PIN mem_ctrl_out[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 311.495 132.390 315.495 ;
    END
  END mem_ctrl_out[15]
  PIN mem_ctrl_out[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END mem_ctrl_out[16]
  PIN mem_ctrl_out[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END mem_ctrl_out[17]
  PIN mem_ctrl_out[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END mem_ctrl_out[18]
  PIN mem_ctrl_out[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 311.495 116.290 315.495 ;
    END
  END mem_ctrl_out[19]
  PIN mem_ctrl_out[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 311.495 203.230 315.495 ;
    END
  END mem_ctrl_out[1]
  PIN mem_ctrl_out[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 311.495 277.290 315.495 ;
    END
  END mem_ctrl_out[20]
  PIN mem_ctrl_out[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END mem_ctrl_out[21]
  PIN mem_ctrl_out[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END mem_ctrl_out[22]
  PIN mem_ctrl_out[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END mem_ctrl_out[23]
  PIN mem_ctrl_out[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 311.495 303.050 315.495 ;
    END
  END mem_ctrl_out[24]
  PIN mem_ctrl_out[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END mem_ctrl_out[25]
  PIN mem_ctrl_out[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END mem_ctrl_out[26]
  PIN mem_ctrl_out[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 300.775 285.640 304.775 286.240 ;
    END
  END mem_ctrl_out[27]
  PIN mem_ctrl_out[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 300.775 23.840 304.775 24.440 ;
    END
  END mem_ctrl_out[28]
  PIN mem_ctrl_out[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 311.495 45.450 315.495 ;
    END
  END mem_ctrl_out[29]
  PIN mem_ctrl_out[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 300.775 163.240 304.775 163.840 ;
    END
  END mem_ctrl_out[2]
  PIN mem_ctrl_out[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END mem_ctrl_out[30]
  PIN mem_ctrl_out[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END mem_ctrl_out[31]
  PIN mem_ctrl_out[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END mem_ctrl_out[3]
  PIN mem_ctrl_out[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 300.775 176.840 304.775 177.440 ;
    END
  END mem_ctrl_out[4]
  PIN mem_ctrl_out[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END mem_ctrl_out[5]
  PIN mem_ctrl_out[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 311.495 261.190 315.495 ;
    END
  END mem_ctrl_out[6]
  PIN mem_ctrl_out[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 311.495 248.310 315.495 ;
    END
  END mem_ctrl_out[7]
  PIN mem_ctrl_out[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 311.495 29.350 315.495 ;
    END
  END mem_ctrl_out[8]
  PIN mem_ctrl_out[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 311.495 74.430 315.495 ;
    END
  END mem_ctrl_out[9]
  PIN mem_ctrl_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END mem_ctrl_req
  PIN mem_ctrl_vld
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END mem_ctrl_vld
  PIN mem_ctrl_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END mem_ctrl_we
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 300.775 146.240 304.775 146.840 ;
    END
  END rst
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 302.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 302.160 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 302.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 302.160 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 299.000 302.005 ;
      LAYER met1 ;
        RECT 0.070 6.500 303.070 303.920 ;
      LAYER met2 ;
        RECT 0.650 311.215 15.910 311.495 ;
        RECT 16.750 311.215 28.790 311.495 ;
        RECT 29.630 311.215 44.890 311.495 ;
        RECT 45.730 311.215 57.770 311.495 ;
        RECT 58.610 311.215 73.870 311.495 ;
        RECT 74.710 311.215 86.750 311.495 ;
        RECT 87.590 311.215 102.850 311.495 ;
        RECT 103.690 311.215 115.730 311.495 ;
        RECT 116.570 311.215 131.830 311.495 ;
        RECT 132.670 311.215 144.710 311.495 ;
        RECT 145.550 311.215 160.810 311.495 ;
        RECT 161.650 311.215 173.690 311.495 ;
        RECT 174.530 311.215 189.790 311.495 ;
        RECT 190.630 311.215 202.670 311.495 ;
        RECT 203.510 311.215 218.770 311.495 ;
        RECT 219.610 311.215 231.650 311.495 ;
        RECT 232.490 311.215 247.750 311.495 ;
        RECT 248.590 311.215 260.630 311.495 ;
        RECT 261.470 311.215 276.730 311.495 ;
        RECT 277.570 311.215 289.610 311.495 ;
        RECT 290.450 311.215 302.490 311.495 ;
        RECT 0.100 4.280 303.040 311.215 ;
        RECT 0.650 4.000 12.690 4.280 ;
        RECT 13.530 4.000 25.570 4.280 ;
        RECT 26.410 4.000 41.670 4.280 ;
        RECT 42.510 4.000 54.550 4.280 ;
        RECT 55.390 4.000 70.650 4.280 ;
        RECT 71.490 4.000 83.530 4.280 ;
        RECT 84.370 4.000 99.630 4.280 ;
        RECT 100.470 4.000 112.510 4.280 ;
        RECT 113.350 4.000 128.610 4.280 ;
        RECT 129.450 4.000 141.490 4.280 ;
        RECT 142.330 4.000 157.590 4.280 ;
        RECT 158.430 4.000 170.470 4.280 ;
        RECT 171.310 4.000 186.570 4.280 ;
        RECT 187.410 4.000 199.450 4.280 ;
        RECT 200.290 4.000 215.550 4.280 ;
        RECT 216.390 4.000 228.430 4.280 ;
        RECT 229.270 4.000 244.530 4.280 ;
        RECT 245.370 4.000 257.410 4.280 ;
        RECT 258.250 4.000 273.510 4.280 ;
        RECT 274.350 4.000 286.390 4.280 ;
        RECT 287.230 4.000 302.490 4.280 ;
      LAYER met3 ;
        RECT 4.400 302.240 300.775 303.105 ;
        RECT 0.270 300.240 300.775 302.240 ;
        RECT 0.270 298.840 300.375 300.240 ;
        RECT 0.270 290.040 300.775 298.840 ;
        RECT 4.400 288.640 300.775 290.040 ;
        RECT 0.270 286.640 300.775 288.640 ;
        RECT 0.270 285.240 300.375 286.640 ;
        RECT 0.270 273.040 300.775 285.240 ;
        RECT 4.400 271.640 300.775 273.040 ;
        RECT 0.270 269.640 300.775 271.640 ;
        RECT 0.270 268.240 300.375 269.640 ;
        RECT 0.270 259.440 300.775 268.240 ;
        RECT 4.400 258.040 300.775 259.440 ;
        RECT 0.270 256.040 300.775 258.040 ;
        RECT 0.270 254.640 300.375 256.040 ;
        RECT 0.270 242.440 300.775 254.640 ;
        RECT 4.400 241.040 300.775 242.440 ;
        RECT 0.270 239.040 300.775 241.040 ;
        RECT 0.270 237.640 300.375 239.040 ;
        RECT 0.270 228.840 300.775 237.640 ;
        RECT 4.400 227.440 300.775 228.840 ;
        RECT 0.270 225.440 300.775 227.440 ;
        RECT 0.270 224.040 300.375 225.440 ;
        RECT 0.270 211.840 300.775 224.040 ;
        RECT 4.400 210.440 300.775 211.840 ;
        RECT 0.270 208.440 300.775 210.440 ;
        RECT 0.270 207.040 300.375 208.440 ;
        RECT 0.270 198.240 300.775 207.040 ;
        RECT 4.400 196.840 300.775 198.240 ;
        RECT 0.270 194.840 300.775 196.840 ;
        RECT 0.270 193.440 300.375 194.840 ;
        RECT 0.270 181.240 300.775 193.440 ;
        RECT 4.400 179.840 300.775 181.240 ;
        RECT 0.270 177.840 300.775 179.840 ;
        RECT 0.270 176.440 300.375 177.840 ;
        RECT 0.270 167.640 300.775 176.440 ;
        RECT 4.400 166.240 300.775 167.640 ;
        RECT 0.270 164.240 300.775 166.240 ;
        RECT 0.270 162.840 300.375 164.240 ;
        RECT 0.270 150.640 300.775 162.840 ;
        RECT 4.400 149.240 300.775 150.640 ;
        RECT 0.270 147.240 300.775 149.240 ;
        RECT 0.270 145.840 300.375 147.240 ;
        RECT 0.270 137.040 300.775 145.840 ;
        RECT 4.400 135.640 300.775 137.040 ;
        RECT 0.270 133.640 300.775 135.640 ;
        RECT 0.270 132.240 300.375 133.640 ;
        RECT 0.270 120.040 300.775 132.240 ;
        RECT 4.400 118.640 300.775 120.040 ;
        RECT 0.270 116.640 300.775 118.640 ;
        RECT 0.270 115.240 300.375 116.640 ;
        RECT 0.270 106.440 300.775 115.240 ;
        RECT 4.400 105.040 300.775 106.440 ;
        RECT 0.270 103.040 300.775 105.040 ;
        RECT 0.270 101.640 300.375 103.040 ;
        RECT 0.270 89.440 300.775 101.640 ;
        RECT 4.400 88.040 300.775 89.440 ;
        RECT 0.270 86.040 300.775 88.040 ;
        RECT 0.270 84.640 300.375 86.040 ;
        RECT 0.270 75.840 300.775 84.640 ;
        RECT 4.400 74.440 300.775 75.840 ;
        RECT 0.270 72.440 300.775 74.440 ;
        RECT 0.270 71.040 300.375 72.440 ;
        RECT 0.270 58.840 300.775 71.040 ;
        RECT 4.400 57.440 300.775 58.840 ;
        RECT 0.270 55.440 300.775 57.440 ;
        RECT 0.270 54.040 300.375 55.440 ;
        RECT 0.270 45.240 300.775 54.040 ;
        RECT 4.400 43.840 300.775 45.240 ;
        RECT 0.270 41.840 300.775 43.840 ;
        RECT 0.270 40.440 300.375 41.840 ;
        RECT 0.270 28.240 300.775 40.440 ;
        RECT 4.400 26.840 300.775 28.240 ;
        RECT 0.270 24.840 300.775 26.840 ;
        RECT 0.270 23.440 300.375 24.840 ;
        RECT 0.270 14.640 300.775 23.440 ;
        RECT 4.400 13.240 300.775 14.640 ;
        RECT 0.270 11.240 300.775 13.240 ;
        RECT 0.270 9.840 300.375 11.240 ;
        RECT 0.270 9.695 300.775 9.840 ;
      LAYER met4 ;
        RECT 0.295 10.240 20.640 298.345 ;
        RECT 23.040 10.240 97.440 298.345 ;
        RECT 99.840 10.240 174.240 298.345 ;
        RECT 176.640 10.240 251.040 298.345 ;
        RECT 253.440 10.240 296.865 298.345 ;
        RECT 0.295 9.695 296.865 10.240 ;
  END
END VerySimpleCPU_core
END LIBRARY

